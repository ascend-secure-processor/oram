

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pnNVPVOI/arOujPkiL97U6I9aCPSoyTEjgpnmJjAwJ6N2eO/yUkxjlqHsbaHU5QhevTw8uu2GKJL
Ca6pfQqH1w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jt0os2dk2xqGb6FC939TDuiJ4FNvtbpeWkKIO5PBtHKZzyGSceAZoiVZjIRafii1e72ZxCM13Y2A
KLJjT91CRz3qfmUriXjni/eFekrD7LvejNqfB3r3KzLV9T0SUzMKo0YFofQcez+BuRcnqbeyV9zp
WFxbUoZFJvcZvNysM2M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T9nw6MsJGqH/ir/VptKsp6uQ/PQx9DuGuUt5euQPRoVpeovqlO1ohmEfwTUM/OWGvLaFsFV1lOlF
l9TgBJW9RbKf2DApED9VdCJ8OD7S6MpupJLWG14bKzGPmYjr1bjCD0OXitax/DGWn+BXD9H2FScU
22RxC8AhhRTOFH/nOP0NjMBWnChE9mJQBeUJ+HHJQwAc6ySDgzn52L9+39mPnnbMe/NhfmdDXwZB
oUR8WcB1VO+wncW/xNSw2qQtbKPt+mypu/AI2R8U3JFuAhokcmehUavAwgNBYJafcw7QLI4Psz+p
5avPLpXr3B9h6NeQ+yYdSg1xeR9xu7icQNmH/Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b452eMsq3LU6MmfLqq9ylli+ZBs3jBd4BzWXyHB89XL/KH+8sbG3ktlTbhX6HEUG3i4R7PFtYe/a
NDcQT9DBH6OpbC+jrj2RxzHef6iQQjMth/bwz2Zvb4bEl0JS0Ofu4MaRX7EBZpu/eF9/DA19QGuQ
fJm6q37USVXXduBos44=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
srzwamru1kuNyQUMjvFQIJwGfQo9kr6wl2O9gBUnLUoMrLYi4YTs62O1Kyw++bTZzvEuiRl/QK2j
1iE0gD7n9cdwsi3ZZhmeHieKRn594lKznJaWEOE8k3cE3mcKzlAOBdoOlRl72M4c6GL0IJq2NgyG
px/x+QfGWQjhp4XZZ4Yx310WI91GQN8+Zy5DZA66Z0uyY7HMAHPJhPWEF1aSWtJvMPUBmooS7Jj1
E/rlsFZWkCu0FIkXPyjc7SV7XsjHTAMPREKAYusMsYCXHOIgw/rtBqiQc8L3nIXRAiPmgHlUT/Cb
GtsXH/CyLhwZrjGiAi72RvbzrERTJD7tHVWPVA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17760)
`protect data_block
Eme0hKynp1zw0MQtsuauBqY6JUvQ3fhT1zXalMJHCPR2a5Yyityw1n2BC3V2Up+npToyQrdXdRKB
o77AxWyKt0ZPeE76o/nREhWKGSEfndul9wjI78HloPxgKqfFFsmfnV3NmKv0cXWI4566p8+lKGyM
MiY8W21RsvfHSCFQIXoDjXPeVPS1eUYkrTrvStnM98ccVGv9focpVM0G3Y/TnaMT2DKQhSpzftl3
Ex59Jg5nlPQ1NB4Dcgm1uM8LY4vMIZ/VMguvnE5lK8ZPK7PYiOFqNOFlctgeMI4l57KYrmFyXSIa
NydmiBJ3VNTVXSaPg77jGaYgu6+dpd49u3TKsDiNBuVp23p/VBT4hvlqa83v/hos/uoLkk5hKm9/
GUwR6BrIzTLdABc77PlLDa1s1L61W59+wzxwG57mVi3zMosnux+NoMz7LLf0FyNYV5VQi06Mz4K3
wUPzF07bgPDYLQzij1p5qhX1lh40TC6K8qHlJEzyDCnx7kWBk7IkbuHonvw9ggjX0zjIsP3XtV1l
qnbHvsiD3uzSr+G4EG94jrnI+SRrk+/oPScSlN0BgxOdGapfDmYl2ldmVnYSpkug733i4JyEmvhl
ABzAVRCUhDX/AEsA9Vz+sSookBaPfILuzOgc4OwMbb5b70YWHWRfdq4gX7+IaCba2r0C0FnrhQ57
WM8yUDJ7p2VtJ9BaHNII0K7xmxd+BF4XlaBmKt4lDn+r83BEbADd0vajFVQ8ov2ho4jxNzg07aBL
ISsmRXswhKMh6cMn1T/nR7yN5fOElSkCTNB43fwdvFAA/+akbatxTddzDRgzgrtSg2kUztlY8xh3
LtJgtnRmcT0CSM22R2YvOdcCtbDGBOdchQrmRA1qVRm87XUzIEO+cLlnUXNvkgKTyY3yfMQy4UPC
+r8ztbqBNhmg/CjdREHbCb3PW4H6vJ1O6bRJFwnQBZQ1/cz/6/jfn0gw3yay8z+jlmXwalzc1pkZ
fpLYpqod/LL1uStRTxcNWFFtbBYbPBPm0ZSVA3Bot+4JbF+81T0nllrgdCLOFWFXRfAwpu0tRDTA
PojSTsxhvdPrYFQtgx6i0nQKsXiRepIt/FEeTHnu6T3w51tRnU0+KUj0jBdYK1/OD4/SKrVoFJDR
EH0QteJlcdCY+wRitl7wyHci3u2vf4OoWuDpeLLMAt+eBdpZCEVYSrrC/3P+fZ9zVAxyAVkEho5z
kxESOtb46/dPpwaz/ASkFx/MqGvG32FKIp6vwVf3+lwQDfznXMNPdpl3fwVq/nBTl6Vb8iwBbsnR
ObLNfQMeh2N9KWGFwgMCM4b4hTUQAXntBuZKS69nK7/CY991/dfTidHhtoGhp+KpzHXvXNmZSTuu
Ye2OyGoXxfg0yXP3vefTsLORvM/HzvbPKP7+TTvhQFlGr1Lq1Ag+1oghdJ4l46qRF2+OlKxZCVP6
sdjoyj/T2UGtta6s+xpQ6epRKle4XZBSxgo8dBAyY83ck1VJOF+Hf+G56EVGGOnjH65wIagPrRxq
2vkt0lCt6lT6rIiKgGfFdiri7pu1GkhLZsLBKiTJazGPrVYg2IuEB+LPDATvwyo7/rtGEWvM3REs
j04EVpwuC7Sb+QJZMDC8bjjY2pNbpDgftyVeVE94lXWsB1UkZlAfgD5e32tiiP9GZNKAejmH6erZ
7PttW7r5JqEfIbT3V8VftsF1lLTFIyIomWTV9k8zjypODm5IpExHQ0YIylaAcqeqyCRLmbkAkIn/
MkenlyIhYFJ3B+z/7K8g2221LkUcdbgmJVGMxi757NRs8oOCBqqPGd1qKh/6AOmOQ1gPqwSSGATo
fgC2Ua1OPM3IxUqWvn2IP2BFMn8Aq+Nejc5O3fESy1+jHpDiu4FbWLXaYoThPWOwaI/hU+nubO1T
yyTpsCjXitDKZfdo+S5ADcnAXwAktBbaQjhwUTfxFUpekXN2p8GUY6nVlZQ6wO/O79jmRNtb1ZZe
J8ZMXooPOIdZlZQNRW/8Gvt2P73lmO0ZLe8wUn6aiEObY3cnDutbDE/a8ixwAZhxLdSnCCYqyjGe
ZGYdI5tKDTnx/fAxN1MVuQADaApcsLbwqEcu9EqenrCJeA10TYhE96s1dj3HSLv45vJoJCQz1A6D
qO6IpLq5oCtZslKaXA7EVmGS9fsCanfund0MCe9pi9a8AKAYp4E6jvYD9qVvZdbgr/lzyPFoj6Ar
KrVhTZFzjRMgp3X+9zcYIfvyzaCJTbUasBdV15EGhf+++arV3IsWGowBXNZ6dyZc8F9ooUthGO4a
JjdMQj1+nSAsoxQPT1QjDMjrpIeTzo0+wRxZOoLeEt045CaQjBTBulJKDvbxtLeZR3P8pdM0kx8z
K0RPILVZEoHQlFHFeJQwApqCuxblCIvBxHuy1KryRXoVRDgjPdjlYNG3sW9j5zxk1vzAFt084N4k
MXoLKwkEIr//ZRcVC7KeB9OVBu70LrEnXARxhg1E4AxRlDukuz8m4G+XWvVhrQ/ZDADFKdtw19Gu
ZpbXcFOW8CkNKN+VJFdciYaqaC8KWdNxKQ6LCR9qyyJxM+LXNC63rqlnTazxgyVkvsDdVpRbm4ja
/JIfamM4HMOsCYm7MezC7lu40P3Tm7d2yOEqvf67nTkZkkUrxu8vWQq6KE9dUYrC+4ba5xDBQmgX
RkZRVgqlsPHfTvXMmB9FdAMsc2uVvSF7Zqji2wIYtADB2GTAdqTZgxx7pXBwp6W3oVm8/CdlWF8g
HWodNFNOvzRWmVon7eGX7tdF/83M3V+jj74J+OMEp9Ky59I9m+grxdiGyhrwuXyVhisLLqovlpKm
F4T5XyJxNya/9jleth0yaUnG6OIqgxSmrlcr17TnxvDxC4JHQ/0HqcTARH6mclcRLUmfyc0hAaQz
GFGUmi5LpMcGSXqzcy3gEbk+1LMy5L7NXhFNta6D44QkxqtjSLnu79cP4AHCZ0P4FcryGezaFVG/
daHCrXJ+S73w/fh7y7L9CEX6rKyOgt6dtI7OcT+rl2eL295SkAB/2NF5Ai6FgMnnRbh+jdjAXKn8
MEeQkdq+QEUADimkN9FdyVJZvz4VOjwpO+VL1KhUPwPHhc+eYmUamteRneWUBIFx6bJeFoo679Ex
yOX4imqTIRg4gIRC+CjlZE30k121c4g3lBBW8fK99VFfaPijlG4nk6XrnInmQd8j4UUArUk+rpxW
1Dy/5+g2sl2B/YBPjFy7jxSnUuJGbS2RRpnglDnMKM9kpKGFb5djEcRyDxnMxcEKOgCPHPn9sa7x
4y4dSdljjEsO8AESVN8TqY8tNz5BKkNH7EsZ2ZojMZyKPxJMjYa1tkjcW5gAw6wpeX8+0f0ifyFA
D1tg7x74ZENWVBn/ZfCcZEXNIKHskwBCah039An5WTCtUPqlRs6e1OxyUTc7F322bmRo9FSrUWFn
sLPX/Yy9hVzr+xdm/EnPsiEBZG2fWBeuag5s0Xr3N8tXyLeewoD4jHA0bxpVlYRTi0arvmEbfLFu
alLQOOT5iaXAB5HBd7nfE7UWwdYDTCVrC8twIQ6QFZr+EKUgpKezJGsiR62dRgGHGtjjFDk52zdA
3j+TsLlMC6k2lYFAJdtcKT7H8LRNBkXd194R0yrAGUNd4evAwzbtINxoJrY9wmRNjCfuDbwUTgMR
4cyjfFbUCxZtY+OQK5eqSzhDdevduIPEfTSO/xwJIThRDBitD1Rpl3gHgZU7nItb7vJAYjCUXzDG
i/J1pkzjFSNzJA6ZbCk8qljsRgMVxQBopGFnEtSo4f0HX3D0JwfL6tyxtYqHSvjvqpnrZCPMjJld
m0JSfXODVDnfyxOPK+sVOu+kzLCA5QHxdE+2gk2PAq6FnlBkvUMt9+LmV8QGJDcP4AGxOG6+qWdY
AEwievd3PYozi9BajWCLobXAuhpqDGFSmT0xDySxhESECgi+iVSagg2IQo0bmdtzWge5CC+pVlgG
sZK18lCq+bjDQuTpNqd+J2/2pVwOHdUSCkuT4ycwL+Fbx7aq/GBBF1RHw9gVK0om7V2zaVGC7kVj
ELuePF+rjXzi6Vo9ZjqzdDo/PDoFFMQs1I/dS3GxMi9nysrQEvuZp6IwOznIB6QZyYWkX0O8NMWd
PYytJrqP1uc14BlpWCaL6dqhVFftFxkCgZkJg03llmICPl1gy7SFN8GvrNfnWqA2812/fXBZ/8zU
izep9Zxevk+MwWOa5iDyWMPTjnJyu96OEChDP4vTh+THYpE7NEnCJZzoNujj3Kte+aJaphKYkA36
sAu6pUzvnGBAGiNg9tse5JPcgWL6wZPFDnDbamSX0nAG23XAbXPDFqP1n0u83V82ztLaag3rVC6j
p03movYXTsnKSWYafSAKS/6DEz48PUzBixGZTHhw0h7kAPy6zw65vD5KpPN16fIsroWPrAECNJ3H
jI5TufGz4Ghu2jvdnaCVIA7C+DRMbDqp6ZGHAFYSpPRp5ZyglOkBQZMkblVvJjA30+fOrKK3Jnxj
VDPQ727hkfhM+0AEDFB/iCPtpc703VVVVWW7VndvrvMjG2WZVR8AWvCQxbmbNB9RvEgPGFUrdlmT
Qu2AzLtKB0e8HtNewM9tI1+B1TpRa/3wMnVSe6V7sxZ5IjXzTV9ekn9PjjhyCUhfO608oqLfH0SS
FN3AH68s4pp7RAjpf5dhoaUBM/SiT2F4yWtvMcKUiOhZZzbcsqHax7XHjTxXIxnobDax90gh+z98
8dWRg6U0lUZQBfFXKxtm32HeDN0C2Xr5Cgk3DQla2PGjdwPOGniBkdbCy0XGxZPrqUXhuV0k1QXz
mjsyHLWP7byIoANcC6Iu42fdcuZK701mcaoRfALLbRXsQGmhMvhYamtdLhLUvzmwAmggE+mMzuM2
mbm86JYvJXmzLdhNY26tLhGTn4jV7OJKHsj/lxSh60NphQgITo+ok7H4OGrKrHRRx+PvI7d+eNjN
0XbXs+HRIvLKl2tNTSWHfKKLpf3vrvijQGC8QnQ+bP/Mokx/0uf1UhIrlZJQovBGhp5vyyHfzQeA
RRg7WcjPHEnkY0AW7bikeQurGeqydS4ee64xmqwbFD6c1trF5m7dS57E9ECRUheWOBr+x1/m1N6x
HUT3YP+eejWYEDvUpEclDW4W2lTBbuqBNiOgeJB6y4kP+4RwiEBxPFfYiroLcMvYn7IpnR85y+xV
fJfQ2NGr6dZAKYmL3Rik3r0TLvHVFVu49XhNQBypxGDKx+75IccWZcDYKPpqo4dLBZAGI98jm58m
K3d83r7kGs6JtyH9JAAVAKcoOt5LXMDrZx3Pxhch23pIXVZXQmJI3u2a624r8M+bTOZ82/o8zD5w
TJGRM8GNIkCsuixJm3DrQaCGFvt4V4Ii9YAG+ek62BgVqheYY/2Mpja2K/7a85dMOr3lS71p3l10
gA8juOia38Hvz7KaOHOP2r3hSZesPya1yTxWV3TfwVg0iN+DcLczMBmslb6S0nW0J9+3zWbIRJkS
wUp5p6KF8ItJR9L6Vjp1co1OVoh6Pxun+tjg65YQywBoyTQ7xWQG2FnmROjQtLr6QuZ680fxwpGs
GXOmJi0iAejA18N6Io1/0T2/OrPbT598RpvU+rW8uvAMushrZj/VsZ+sFogM7ROhu8mjdK4CqWrG
DhGcp6kVD/BohcP6JoRY4SCWa4xiCmMwpce1/Z5ckMPy3K5lijUmqjUnm/z4EaIUnJbL94BdNjaS
sEBuLQx5f6v4gdSlDcIn/jBvLwl6zQUZM8g3dRFy8KFGFf4Vh/wi2q3cPh04InzopuMFtE9Zi8R1
T97IyEq3W7tDDEB0552yDPiFHSEXa53YsjI0X7363sxmr5UYXcebilxvUDz7vs9h515QMvf8ATVc
+6+2obJ1+ARJfwO4GPMj421B02GxqHuOmd55gkbPiGJzseWbqxmKjMoCotjKYpo7N4flALYwrbTe
+gTx3/mTbo2UdgRbpzMGVRDLKt29l7vCOb8NhnYREt22j7bSFfnunA0Yue8GVdpNFTKMscKfnw7/
rBefluQIsw+xVq8bB4CR+aN0gNseMoSy1WQymjDmmpZpLYN3EI0vsyExJE5AxqhznuSVfyhDPyYo
YHvcKw1z2uKVjCNBWZhYOiZ0vyZSB2j0DkN8WvC67mpUdVtC/PK06e42Sr+BmqMqw6Meo2GzY/VW
Vmju1HTxuVpb6SclWPn/I0RSrVXcORRFcQkXZk7LHyA0oD1BbbHN2YInuo0dnmBK+kiZrlvM7fHY
n5QHX8WP3lCUTAnJWItFpi8Ub5vvVEf1lrnpzUAMhsLfl+DYvkZ1yu7fJpOM2UCGNzod+35zJgsW
K9K0VLFJ+0hdFOqo5I2T7WzXfQJRz8Q9o1IIfYOD0MAKfYyT4NFkaVZvL/z2oY+/yjgdmEAUHjwT
CQrDQ8n6I5OLTqbDS7d+OKviuiySx3546DDGxaH+iyi5n/pMyiC+hNT1N8qd2Yp5+mT+ABXASQWy
bNbnj8HxE8dEMLFHh9O5K33V4OYq4Fzs0RkI9RR6Z5WcvQfsGR/UgXtcR1iahV9PFx7cPKiLDUqY
Rq6e7O23eqSH+c+cIUPyeekH6eDgRHoDCwUpwtfTrtOY7DK+yhU422T3IborEvyfnxqaT5tr3fjy
vOVHbT30RWnKKb2a0TOORjrlJCFsZgwOctYRxEUHiKAhmhtdaxG0HENJ/cuXvRspun/eCgqSwmuz
QM8J4mWynhKb8LLBkn3oCj2roGoN0QwyJpkwPT1uYDjj/NQybqhbg2/34Sjk375TMu6xZ+U4coPY
vhVZfvpukDFrQ0XlZnHR4zEijhmrOhdU2uGvqd67LUD8XbIMJNnUnSwza5xVYLJ1Lh6xlOexiAVK
ebuD6x2igz8d93ZQPhT+foiDrPBI3BedQJDmBx0hghoKS6b0gHXoyvvvnipJnSzeid797nRvocWi
MxJxJ+SRouHS4PsRzQjHUbroPt9BJmKFE8bnJ8znMRpy5BPszqlbc+uz9Qpfk95CD0BEc8iNGFGG
4UxXhcVoqQxJlfVHl4fwJ75qYrtHiwIE0ekqKq9Vy+3fv7IHkFafC5gs7x7Lx+ynhCp2mtJjG5PX
IGd66brE4wV+lCIweDYaYRFWYM10l2O9ZTBQliDjew8m8Z4qm+f4dTUhzjnODiOqCHKDXmsce1Sd
2sn+H+1Hjv5Q07S3bbmysxExP2W8aLQtRvOdvAfPDOOvfIaFmpOfcj/aiN0potjiJp1o4eSDe9Hn
qx2Mzc6O5t/JWPpToGGYF1QrvHF8lfvbXesNGjmJYljw+wqrYt+Iw03Mp0SAlyFg/MsFdmFoMluI
wtl48r4ccYtKFD7kR0ZV8q683mJbsoAFOJOnNgimZ3WDyl3tG2ZrZDIDGpPxonsvaEzEv7zA0vpa
3twP8m3Txwl2SSPoxdz38dE4ZW0RmwWil2Z/KlFU03M3qKLvMPgM9iF2YexfkxMBl9xjIGvJ6C6q
NGAJAnZskyVzFYeYMmLspKCTndLrdrGThDq+p+WPH295HS26z7XzunvOLhY+QfiYOgbddah5amq5
LSohXKgMHYq2uZH+mL2oA1YEolB1TtKUgIJt9KAVBFFnVkQsyJyCjZPIcRhhktnJVmsCAmwL7tGP
29uHdPyyh2LQjEsVeEyMt1MBO9uQ0zYi8CNd9GC4xx/H5zzP06BTi10cSAXCMcrAayGHvePSmjzM
EQSFYv/IQAYt3Wm6CsKSBZ4qIANtbjOVhwVze4pXu5h+vWI1j7NgANNGnC8YHVeUSS4wHWs7k+LF
/eTQ5SlRtQGQKXT5zm3PcFrc2lbSmob8HB5UOM2eIKnqHnFVGWfl3d2C4HCM3bEcRX+OJH+ZHzyO
RcPnbqq5ROqH4JdweP25yK0e+xCKj4kRoFwOTREUg7rfY4DWK3dpOZ7C8u9ZOixL5C3UctWj2Rlb
RGqWcZHBTvkepFgfd+3Hzdvp/ofX1efLFE9t4slT57yP0/qZ0CSTEwIhm283ZK2LWJwGmXVyd8X9
LrtJD0wK/L2qwx7MeJj7LkZMsxxijFNaznHPEek7vejTdTm71nTmcWhwyaE8wLA4dQoLZlT+N8Lw
cX2RKCfR28WIXz9IP0lnc2yQzcs4Yg/JO3sTf6OcVFv/YVl3tHvXgzRmhsbJZ77sdGkENESGaZ8Q
EcFhsrW4q0v4ifqtubtKgNIXB+NYs0+g4JKe0wbEKqVPjfM4AbUdivA3vBnonYoTMsjk5guJIKyW
uTtVl9uRRE5DCdHNdoZQFbvu7xfiWL8MiJFTfAafRo9tRF2oaglw5gWziCPeaZaLFvxdjzVd1Uu9
Rfx4GLP/ozGDBvx3Rfnn/Yyuhnml6QAln0pIxK0jkoabN/dGXpgZoAemFK9FmaIpTcY4U5Jc51hn
/mFY8li3Vl6/9SwnJpuwvlDSYumt2nl0dPF3CKQKvd0jpPWUfliAGNC9rpPdU75noR5r0pMMOCi+
ewMnIEPrh3i0eJ+o/s+xwtMDSA+uSe0A22Ugon+vMt37paBR13eX3ZBVeTt+y7YPYgElgTlxbGld
9aL3g2p8bn+6fLLh4QS0BYMdk4ajCmpLZMhXv1nP/RxISR5+qsmPpdti5QdnwLiTHA9CpS0un33U
rqWnRS1ulb5etfckgr3ErY1p33Fyl2Qs+C6KmuyTxXYnl2ktvE3L/qozb8zUYIacgResQlXwhE1u
SoNWWqpYY5lTmoadMgdr61ACw98/jJClf0mRhwoGJGhaGmvWSAolOQ706aJmvLxeKfQ5+6B0hOAx
CLZe/D3vCs47LQZAkzH9snJICLIAlL0gd0lzFmdVSjCn+86KR5HoGX13UlgXg8TRNgGS0ghwIMty
1XsGtNk/ZDURiPBnQNzte+08liJ5EhiDGS6uBm0aMYJNBkCRcSFbQjpGSk01hC1KOjKbj4eCI19O
qAJA0q4uBY6W9ArKLDH69t8b/sMLAKtfYD05lQMORcWAtYyu7kFxnrq2u0c44n80ibgRivM7VcCX
JU5E0qGdTSTsRgGUbXX5zA7JH0EpzKzzLxk33qQLUrhR1xEljQoVLRkS42QVBlX8Hwvv6kwkzk+b
BlMWPSsrKt1wevRw8KIRuJr//XPu6KtU2owY3Yo62kwUqjSac2A4VtPO4wDgWQaAdiWtgVEZuf1j
JUWhQjJ8I10qtbTVGbGLc6woPHw84FRJf91opy4w7kc3OdDZ9woH43Jn131AgSetmKk+hahqFp1h
detvU3O5zh9cyAnplutdioZ7U0G3w4cxDcgo4c6Ad/F/S7ElO4jSXvFGQPiXlPuMbRoPuMED2NK/
lvutR2iWov8YxudEyPZjHXks1cFioWpDiv+65Uz+eDBMJNB6Ug6ut1sXWsUg3TR/KQLwfUifj8EL
26c/kGtOLvtliyrOQVnZHPUeCK3tQVCeTYB9u8rgGgs8n49T76AFTgiXExG35SQuNB7MoqaUCzCM
L4Un4CHg6brGP1U1lfteNNAXe6NGw49ZeQoVHd0E6HNB4vxan5KhI7UjxCJ9TNleNSE/WHlMJc8G
9RX+On3fCnt/D4Q2A3Dpx+IVd+ktGB+UELCpKNfBJD3ZVVXXXRFhRD0agEkrW+YzWcdJehFtH1HB
eiBSLq34y1tN9kTW3+D937MbZx2E3yHNukae2O9wGpQK4KE4Ye+XK7IIcHbhTt+NpjGkZvwcuJgg
xk/a5bHomErLcL7NMCmuJZ3iaQfTOesOx5EaTrmUR9lU18DaKRZNhqxYDXmEzMubKcAUn6w4ZvGV
EPrHppsfNsnYDFF+nonaG020ODIJuniH1Eyl5BRZXWF38ZXMuei+iPgpNiFB9SOG+DvUBaUCfdYb
3a7FZi/0Rkm0STLT9hgfRf92QeB9Nf0Ym7YDE7feHjCydJJyHaOArbBiguzAIDBb+8aZyxUyFDmQ
zCu9G3LHRAj5zOGwkxLxYs0C7J8GUd3gubbO1+yVhS+gUr6XB8rgugztUiSv9ULvmYW0YJUvsMpX
/VDB+28cHtEbbIjmdGplF17lOSHYma7uFixN3cg0zFoXka2dFvA24Wx3Fo041DwFwLJ6hVkjdBWA
YUZAUKLGO9QkZN2hIEQJ+Io1c7DJs4LLFE5fcWfxH2VRy3nMYdaGG1InQmSoPtA4Ek/YTbEW/DS+
LVZmpyuu6bkQVSW6D5SrzlyAGndJUXKkIrCskmPF2HRSTMskMivaeVz/XEJutGUnwSNdBJQ06ZiE
G+zrxLzYazqCko1ZiLwVJdSPtwFveGtD+QWGoQlgSY97+I4N4k5p0XblU51EcXIW7dZPoPmFP53E
iuLr+La56Xxhr6xi6jv/7g1IlEE1ghcCriWkVURY9qYI7yb6b5ohbC/rlOD9rXzfKT/jdPjP0XCB
d1GVoS+JgDgVVY4WoelNHLKvOp8lg2ze5mektgglMQ1pjFEUWc/QTUQeW/M5ydinu2kSskrt9o9X
Btj9+aGSCbif1npbtohczOcfsu6KIRi004Gwem5MG07YtNhOFCU5W5QoVmQriZvQluwzt6fUXmHZ
LRVQS4rPVpnsLVi527oFQxJYvaTXSnlOOdlVBa1R//2t60azaDmpUO5rgr3UaQHsfj/d6l/X+LPF
buCUIKowW0v/MfXUIPZGpqMmGH+5TdwFUWg/APxuvzWE1yF1nDr/0vdHz2My/UKK4FYPS/6NLenP
uJ81vBJ/P6PXl4BR7GMISDaO072mlc8m4RfnH1p8FBeKo8PRznYCOksqtbL7Oz9zScVkVNum2qm0
4Pmvf5MTSOX07RPm9hBOkcYvsE0oXEMZuvjt7xN4GSIViMX+kU21wEyZZEcRQLU6jjp77MGbxxWb
dqPiWfz/1ysha05aRs5p7U21ofmxnkUIqVTMA4grOiz7Kpug+geK1txD8woXR6NbCGddghvMpL9F
ZjrSJ4AuzP2mXL3cbjLxZvrVBUB4viWjc296OAAkNNR86Ha39utDW499VXtDU+VxaK+v+dss2JCY
UcQnb2Y0jwAltIAsc562UHNRZLYdyPHXQz+isnDRsfhOeXiCWgpyS0cT4DUzppV7Vqqz2fXzhjwD
vpySkML9EOAhfePQFyWaV76j0XY8Lo6SX4ZVrY3DBP59x7cnnjj/FfC13aBbAtvyWvNJGifltICV
WzbKEyzNCMUb4MS61b9wnI524owk7TU+W5eENmR2NCdxaM9rqixEeIyogzGW8SBBYQ4h/VNxAdil
uKm5JV33PMRiQR2MJbu5pCGEhnZ6ZQbGBloCDQ9WRq1riBFvjV5t08qeRl4dUIl9XNGEbgu0Rurx
INpryGTLfCfasxI94THUL3bxaa37Jo+N1OPjoX2ABScnq7rO95j28e4uzZScl4msOQjU5f+gBL7t
VtAcixBaR5d5iyz+zhm0rb45cdadq4CtIeFYvx881gMZNI2xYjGwsT94Vm9sWV7vuJBNs3v6Ssm3
7oBL4ZEjZ2Kbqiq+huyKvf89Dm0IXXJqLpazsnJ22pdt5OxeDuzc9vBRtD4BNUZYAi0wjEwrgpER
AY5+QRp4H+N35L4x/gV/NKBQx40Il0QvIbJq8qhNlCNWv+EPb1MVlHjmCEexF/ufP3stFwjs5Yuw
mk+M4pWaTAkZ1SdTq/rQ2sVzOIn6D0XokfHNunPzQQf1RmS4vfbgi3dktR/wG7TUwQv7liUFf8Hu
l5PyJOydEwRgiPRnoIuu2N8MahVbNmVc/G4xhZlej35TBi+sJgnGES8SUZ0uw50Zxt6faGzs2GzD
2A9ML2afaG9Hsp8A204h+FVD4OMShrovJSZv8ABWPAJrNZVdtQTsydfogSzFixs2G/dgHJiIudbE
zUvLw9bSygy83SpQQ/H1OoouhY/9ljiI05iuqXZD2fW/s3MEMoz04WG1IJrAMTL00AqjstE9owjK
sazccL7bks5oxLExPC+dZh/xTZKJG0WwFwiyyDYfPWRR4ihr1nx6TgqWUcxAUIsLAs/lvPKLKyi5
NV/iBTGc5/x5zoGsuwJnwFOI3+luPsav0IcZVHceZq2M1UCJTD1iVERCD6aDSqNoKRGOI9ZGiYjS
BcAyiITvd3P/+dhnMFOQrMoynMyiPIWRVWG6Y71ZuZERJx9dUJNYEjD/0GK2aP53s+1tYvjDOdH7
RUcqFRmMyy1/GYWy6ClMk6qIHr8Ly4SJTTn7lPbFHMPVtV21jothTfR+GNMAq6ZFzoWgX4tkwzvX
esatVG9lnXu/Zb13T9zFzxxBUVDvcRE93vig7pdzxyFGzC30vqoegqLLWAwHiFLR5RTBKfPhwHi5
3mLMZkzkY0Xt8jT+CO/TKNO0BgWvPvcwa/FzzR6y2sA/6Ac5jfcAerJvVvDR8McJ9b2uXa688LHy
nb58MeqJXcIi1mUVlDEB6L/uF45Kd7Dvq9L/jgewHuNu06z7OIcRxkPvfehG9KUT0wlMV/pvBhZe
6u+sd6AlRLrjfqCkwISLVQgHU7V4R2FtanaTlKUeylJ2tMT0tpPWFKchxWhiuPd/t85/VOZxfYzs
biUSgysDjHsnSLY8aYqR7NdY6D608ekheCLkoBPdHp32NQ+lprg6ebwjzb6jsSIJxsAWu36tYEgc
oWcx4TpdhZizevWL5Tc8fa+fhTo3Uyn+tidS9/HueK+xFGbab2Z8fcms82VTpgaUX0fKGAHQv02M
ylCbDPti4yb6RfaFJf5uKuVQzWNTKE13SOErPu0lxlx79gknwHhUB3Q2yux6k/PazRjVNH9i1mWn
zwrXtyYoCqi58nWRLfwQXpHEC/ClVVw0+2N/Hn0IgEl0dbHaNnQ71L1WWcSLByHKBpwPcEv4ZVlA
S0fC6Z2RaQCrOgvPhg5NiW+4NNs1E4r0ZyY34BEVr6UrUfYk3z6m0ViDcvEqb76kdH8+fShH7K+J
Z4S1jklXMzCJGoVbgBo8Ih3w/HH2LP+jrJawcRBWemJURpzWGpBiwLmVqSSZ+MZKz+KmWbB6ig8w
mxJiQdlCmxRtgePNIbNjz4Huch5xlygo/uMLOgB+GRe7Em5p1HrPggL+vJDgPkqLZkICQvBOOvUe
Z1NNOq1d2Jb20/Hs3sQ9eHz8xsDrwJEUW1wP0ymFsz2mHiZy750EVIixXDryYte+6bW3DHFkquLx
XgDM2opROkauLAxWtuYiZtmhO8rHvm8NWc6S88t+NcQrRIWsxrDYENyooSobnnIkZ8tPT0gzw9lL
srossMD6zYi0Qc3pOyt6TkSIAdr+YeTnEzZAz2O41noFfI+ljewXIQPajteODXhK9oTzXhGT02hP
JxZMja5VZHjmy/sdPQxZPGzh+gMmOtgsj+taCeKLvesNC/KpzogjyMGmjg4e6QuwyBiVFv8WujX2
FmScOqN1X+3zcriRJk9xFAC9ku54IMavczzFYVcgVvLDlWt60Pt6+lAyaK+41PMVOGkOrhhHwpJr
d6LH1rybGgK1yWvRu2tBlfFp0a4wA5t8VTNGlMztv6iL6oZIu4qBPLSzFFfXQ+Cq3m2aj4H2MPCe
q8VVO8g+/Hxo1/Vi5B85KBHlVtpsPuVnabdfjkrqhstF2F3fPJ0E1QPQmx3aoOBLOCWOSIoebmML
KfiimKF7+fyWyMkoS4IE9ZVH0NR5SaLBWizQSeB0q89973m5w2kCQYSg2sjmPFm70NSc0y52U3Et
XowwNxIKtyycj4Jq5jWanuJdYKWGragd0z1n2dakRtL8I6ndImfybBNw96PAMjzVBs5ju1+NHyuD
rQ06NTHe11C3UlxI5Dreyx8hLGEKHDcgZBD/xd0gFhTp7h5xj6kK+on8nZ1waB++XKsdHJnOXdzO
zRlSbZ1TcfUMrT+b0y2xfHA0dvX730WlYpHvWSGpgjkvfLZmlLX/jXDXulgJnUk/8sSkKtp18l2L
8kuDdGyrHRqFHOU0gftV7J/ETxDNzovNFoaHH8HAu830+Rk/jQG9Iqi7KO/FHfdcgydkPXjn8W65
qP3SSRkfxx3x/800NELs2/DnqiW1JEZTFSThEon2JzTE5ctNawKg17bP3nUBAMyDlt6QHQbIGpom
vmk0Eu09IsclUvdm7XFk5Q5Va8TyF8yMTqL0nNAEA91LiJJOdsyB5blQIziYGFTeeyVtC+l1szY3
QoRt32gwtZ0lPJrRkbsFR3nhnBbijE9hHYt9z3z3aLw0eO1RQfCQ9W7pIgGyogNF3qt5Ubd0iU9g
0Clnw9Kadi5YQ8cYFQ+0NpQDP7sQgJcjCjlDGhrAoiPL5i6ClgPIwqfF4SJ4Ac912hrvOHS7d1pm
f1piL9yuqbOmYRtIL79kfDds7RaBflRF0zwMRISEK9lfzwm2123UNzTfl8mUEVKED5rCcQaNkjyc
JYLEBCaL8gBID+d3vS8XR0ieEyph9DuItwCc/3gFG7PFKF2xy8PafrU80JaXr3eDFi5ADOFtRpkf
/E9kxSmnGTg4a6n0PaVmJSp9s5kayEgIqehj2JD//JfHjlNzyoh+uQ9NDhfYyUHdzr7lRGRlFBgn
PE/aUxCDRH4qHqAgIM3ORgXzDWcqnrXLKpzLmZRVFkj+FR0X8z24T5s4Xnzqxa2s70gXXtgLEP0u
vApUrPbI+sU9ZXAYtE2DDgsjxEiyZ447hOxWg8q0G8e3Leo4LCROAeMF0tx81bgrxS6Ooq1VSPjL
1+XEaivzXwg9eCKpDGpD66N3xpS41nHP605GftyH3IFXU4YQeUi1DltU6sTK5G3d+LexKqynDRC/
P30Y/GaEfCPOJAjaWUJaEi6Z/ZLxgF4OKdsZePGVkMNqWtkNvArQ9qa7iKXlyrXvUswmIDWe9F4P
wEbcm+b5lATxz8iqpFYfyksDcyloL0NQHRekiNoqNzy0nYhZtmhTkGg0EcrDkh1Fcbv01oFFtaca
vlXzNQlaUsIYPOK8jtaQQjGGG7mOgYYMcSRqiI5Rv1MHz8b47tZjdUHrKUMXJPklpg9ptn82695O
94/W69Dlnfgj8PAItrzS1/zB9POcjpp7AHRVsVIdh2pYknTE0gh1ROTlTwiUuspzQCqPzDfrnqmQ
Ow9D5MG6ZBIqiDELkBs06EqCY3ciJNkPTjGIi5WThQLHR002nBiwlgBmfmEiIeKRK8YT0VbuDGvE
ef4evz8youH69r30gdVcZmNeTHbY89vJNoPfDAWQM8VZOwMQQpuTJwrRFWlRQuhlqkkmwNleGGKX
XuWyFa5e9d3A6akYR9/TaG/W5xmVRQR5FnGtmkG/MThMAxpTccpyTuOs1jdqqbDJJSZ9dpZgyGw/
Py3fIgQYpongZnEPGZ6pWJkydR+jI0BVfw7yTLn00P+O0cZc0PlM88PfO8SGrSh4c8hHbYvW02WP
MRdiXlKcT2DZGWS7RA4pIf5P0NXVXK6OAqMJzm8WNCyP+7Cv5noA3ACjROkOxPImR49sgTtCCbZX
LXK7Dt9HRLHeNu5gqzOicBnuy5GNYtyqtLt/74j/TIFcY68JsNSVvFcoYUG2qhY+jkj6NY0IkHVt
axJjmeH4bDikqLnmtQ+ZIjSlcCxTLt+2D+1cMp3D9BN4IL07HCbN//TxywEjuuP0o/USH1H34fFC
ZBawPjM459wQ7K583Zw7GNArp0GGBGTuQBC1mhkuw8/OvdY7uhU+cvdgrRYvmV1mWiFqPKo3HQ1V
9EhmeQvV6KizaPbjctQ8/kmBGH3LYFdSAzBAfPyQqUPZmA7nQCdzLwJkJEwI3ad2Z0GEywVdwRwM
rWejOfk7Y7PtQogC0m0JlM6siRyU3pP/8zO0FaiDMCjkVqP92d5P9Vzatar6XjCAZngd8emHjIYt
Eky8fjzkOy/wtRUnU+SS4GD3ljiowTWcUCZSaw792K+TMGYVLI0N6fea5N0sS75J6svoTyA/BWfF
BfSuqQcEJh3Q4QgXiH9tiVnCoV88APV9FhWsqIAKM9xQ+oltZoqLLmy7iK80uq3rh1KPYcKjPXZj
yEaYxjfL8QNGJuy4WWQJHNjuDhJ0wc1glLzuSwLu2dWHu4y4un6kd/S48yf9f1y1rzzYPrN6XrDh
9uErQDuvOe5O9PrdV1J7xkOgKFYUz7AUlzeUb5IQN1RlRSfNfcKU+cOAYAQ36WvRFsl9TIkxDlt8
AT7A2aNtfZwaixe1zdwG5EFl4RrJNPoQUXmjSDCgpmpCAQt4RhP9DUgwgO2BfhEo9/WQfRBPfcsp
DKIeIY4oeDoNpZ5O3qDC58LZ6V2rh39hcMHjZw2/mJpq6FeDjVY65jGGTGF/nfr9fbPkn9T0aNKw
NcpzMYmYo16KJkGrhHEeGDWWJiY1JGdHtsVmrfhpdWPztsTIt0ifvAbEoSwoPSdTvd6IgnGJJ2xm
IZ+WAm9ehN/JsADR/nzQ2S7BMFbJ03CXOW2FrW83xrP4pYmqvWJB+9NRj2fm8aashx/uUPsA45Wy
tsvK/IeXx+JynhI3aqSUaxztjDmwUeLJ/XG3CBjT4cpVHqBx4VsYeYiUMKKvFA0IOtVL8bo4ATD4
LqayjUCEZ+hr0/dTCZr70pjbv4dakCgxsnrM6gmOCItN1gETuduKdNdM1/liKDqAE3z/zGt6SX/0
Lw0ZYOB00693pZetJ+Y3avKt7RLWE6EbJA2UVPAL6fUJYP5vogLdpx3AhQZIZZcDB+MUVaWnKcRa
namtMkiM0Nnc41YXRdKz5CyRWVZDEIZFrhkvqCwHvi5OSgbkfm8uqoVDt4JijdOzJju4A1ZXJh0D
m2bwsMXkCjOf61Z4EmVxfXRbAdrRW8gtl1Yv9yFXsQtBFAA5kYn1yKWJZx6X37qhtvxRaRO5F92T
IiVukie8wmGjoo0yO6AeLcVe+9KM2wt8r4Pa5riqdYJkn+vB0oHxnuIx/5wt6MG+JEMACAqj7Y3g
qYbRM68YAdsIYZTnTR54yodXlcfSTWs9HGwxyEpx5zKkkH0OOMOiW99kRDd6GP1sMNiwjFLc015d
9aTkj1bFiHXJO+G0WPulXh0R9Ac6SZdGA64wTvOQxqYmmH9Tlx3tuaxS+rYyKwLEfGfgdS03dPKo
tSZ0rlFG7fJlDhVy/mLXCQEHMM/gyaVpR9J9F1CMP04g0lslwU/90z0bU0ERbDx9iA/btFPkiQh+
eIXY0RJyOSPILGqbWeK7TgDFj/VnUdPa/RNGFBlXi5tTVC4HPvhwGj2/N1tVQXFbTPebsB7ZAvj8
zZ/hZs3GvJaWe8tgHBNZDetFMTIakgUlsZY2YhO8bRpfF5NxUE2IVGFr8V/3JRh2WTV8okhgpdMx
a3WFwvMw11DSwI/2W3Q9kl9R73RpoXXunhzfTufkyNJSqGglMigge99a+F+ykETjoru3S9ID//ml
6lpsjUg1zoGwakrnF5FOetg5uKvMiGNN7XLEqVHLzKuYMdIZ+fNZnWZAnwQFGTRE+T50hRccj7ki
6jvByapX/EEW9jGarYrZrpRSrDnd6EXygMwb53SX95lrqKtZPQFongL3FCs2LrW6Ml6kHxpx93fc
JHkOzPFZ381ny3yAcauxm6Oenc+U/IdzWPa2BhHz/qpNjpqsq1sY610bdtCop5WcH/UyR5bIvgXi
6YexDdJdSewWUBXsjZurqy7/ev2PWJ8FFhjvE11elhk3R4lL8ePcnX/Oxg5IY7sbZJBhBBJqZbka
2fqW+MWUvv2X1mCYaKa5yaJdW+YtS3e2UZojlqzoi09va1Et0BIlrJBiY2MOHnClMrge9VwrUj55
c0iY8GCRa4BpRX9wCepX1wK84nnvYWI+Pze8m4qiDxLcDMmFi1Q2Vacp5CiC/sonbr5A9EzcfAJi
/FS/nSBZ0UdbAO3Nhi7ZI10k596aYS1UtNVlED1pNnIqGcql+anLU+yojXxImcP7linQhGPeHD1U
RAS1STlBI9pLgyo8phjpwBkaaJhu9njZgXTupdizwPEzN3ED3WcYW5e6w1KAY9HasTE3Fy1XBgTD
n15q8qynDIAGTMPoKQrXUBLV7D1QfOpCvKMSWuUX8xzCir/BvWxKY3fCJ8iwDQUO4qjGLVL6T9yS
FQQLAZ0TMGnxdB34NzYQz4LLLMVYvw5+/g+zK+4WD5faGXZqFZYKLq7GFOgFiMu4DjWLmgh4T/Qk
aArkyyzNxU/avHV6VnXHJbyZlp+kLAWIFfEbbxXMj8Tg3BpVeb6I8qLSkjad9Fy95pD+10aHO6sG
gifuIgacOWsL1b7l3q++6YH3lDTVkPJsWGJEaE8vJOaLti67lxWMJbkUOKExyFb6VYnfBQGgnNuH
xalDwf7lIXbEjZrf55lQC4zH/45CLhcuDYpL25WtSV6DceZAoZLs7ihcuJqqqQubuqQ051rDnL4I
7FJqs4zgGJJa4zNK5W6QDSA749tCIK2Agqh/XUnAFbmiDhswd4698oP0SipRvwWHc5uLY4EOm7nT
jkrUvi8Jos1hvgxcU1faua3XoYTHh3Gyc/MIbEX6X4TYfRl3Odp378hYRebt/qhXJfbl/WFJmokL
iPwuIWvdRzcLEXQxims1zOGpSumVGASaADDEWBB+QCrDgXjKsCEc67wonqXJmrVwR9bMUvcl4iG2
eKr/oIoobNc2swDuaerMh0tL7ekk0pg2/K4KoUdwYJXKw9QSETxXRdpjDO+Q561dZZ5gJznjCyuH
z2LwTp3vZrh2mvFcInNYs6LbtWbOVgj8EPp63n+L6r5ZyxB0RduO6Zx85waunBjC15+v1bfkuQXJ
q1i1rJq4aj5EfRTPtIL46D+CZ6+UPOSA4iPcN4cTVxbJoJLyf5pYoTAQczO10g3+sTvNfwYfXO93
FzCDrKR6xVIkYXBZ5KdRarOYZf2blNS1W36t+/XUaGcNxdx36qt1ZuyljJBh6+cbOZZQ6BAUEsqX
d8l9714wSV9+MwE+xoXrMOHICh1xH7KYDjCUeV7qy3ggs23fBpftqLd217Bu0f5ewmt26Xp/Tuvd
MMyJeozBYuRnoJwsrcRT4PmEK9HNMn4SxblwvLKJtnVQNb+z4YyERuTpOXTR+xGWD4Z27+InUXMr
wUDWsEuyGL1I4k2V1U0rha7pJSDMzRyHwkuLM3VcX1RtmIyUdyUkf26uReMDTxFUdq7yjQk4nRkC
+Iqe6IEZLFU66jmsZnc/OsYHOFJZHuN8X+MWFfIbU8fNbhIntFwQ8KQIYiIpdczT13eLHHbn7LII
BBPKDNpJCnJa4C8N0LYXLKEVwnb88a7iUStyJsRQi7FTd4FH93yHRUqONvLCFnUYnhjczgGhmt1D
yiRomoDq9/dh/mWK7f5V8FabFiwLQuXN19Bd0ZAsOymc+HVHZ2XRLpytPuYwwsaQOU/QAbTMk0uf
UQ+qm3Zq+5HMlGY30ldVXab2DVIePJ7KPdUZ0xcnJH5YcmAgqbBDUOvz7dNvjMBZcJzyrL+AiviO
/LduWPDMI0iWjk0RacrCVHG1nxxpjBVS8cP7zJhagpE1BTMBmJsgLPG7lLrtcC0WMbu6KeKbFNnZ
JsN4x/IZqCcZrMCq/AP1MzohEsx7i/dwoFFmtBNZLT3aQiu6Zgze3Spw0H24LbT1npjo52EFzBfw
gNQwrGLSMBz3+YA9nrX55/meorPgDa3Ey/C+hXyysbEuhDSTwgIwrVX/PtgmLRI0Ii06KMbJrsVP
IhInwznw2HcbjxNk0Y/WAh3WbQgh3gtKYbBM75qXbP3nUeTfCpfF8rxtvAyO4jo421WJMpC1bn7V
fN92Rd0Qa4vN3Ij/Y9UOuNZfN6vRveVkvrAcuZj0flCUQ6+xoxaYX9X10iQOpItA+bMcPboS7hg/
/7JisSSTmmRYsOMDfWjy/NDDo4++SVXX/ymVUoqet9uouWz54EDTvToDi+pmwoTrz0b3aOBX+wLd
pKgk3vk+g5vRi9S3f3N/yb+5p5jhVnOu04KseCHFMF8GgOKlRWQrDK/mmaIiV+gUqrx6ufgPrD1T
N9T1MCOkO410MDrmMAzl793RxyLRE4Pnut1LwM9x0ZLoxUP+OlDro35leWwrm9k3lMpf9MUsH1Gr
jW9HMNX9HSsG0ZGfB9qyMMw15qndhRhmXARgne+AW6HIkN/KT0ilVKAPRjo78SMwK/JT7av40L17
78mEPGSeTL8MSNRd+fISJoEj933m97o444ncvsSgNBI/B1UyrdDPDQpNtNhwoNjeEnO/F/Uprza2
VN72Ebqx3lijrapH5mK68/2uW+Iw9gc+mB8oSTca2GdyaTXYvcE3o0MXuYZalsuFLU5Xwy77NTGg
1GlRTdqoPlSN9zjwddhZHeUYgvwlflgCg+CYN05j1s6SoyDHLw+RBPz6Lowf2Irrd3MYjOKxNIow
Fgk97aUO6Bi5XGoG1Xc76QqbcMALSMRWimOh23lA8/8tu0z6ffaOsf2rqz0tzXdOqYoqDaoMFy1q
1gRyK8IQ2BiWeSpKglVK57/2TEdnShJm7mIqK0B8OazS6Y6SAsUNDu5SFbpkYw4dmDRPPXBYIsxx
PbUyKYSbvldzMmbMStM4tExoMg8QF213Z6vj2ShwQHrNrfhExneNeRdRDCJRK+K52ke4WoL/WWk8
FLVxNaOm0yfMzMOE0ZuMF0cVq4RWA688erODV+tcRya2D+88wcIi9CXoL/bhx1WJ7VF1LW8OA5Jv
vvGXqnFtHYLuVtniW8lgl6dFMzLexIIpaHqcVKRq9M7pr0ADwCLxubHwKlW5EVirNW46cvcSpN9N
8HKFO/9hFwlOidHr3UIlVqZgGcCJb8hLu/exqCFbNLLVZWL7mm9HSR3uNtUBUGNf0CtqBptx3X8f
v7aX6RCTLlPvYAc6uCFRcMOeIDHYW8bXCyx+x96qG29yUpvc7LuzbarUD2Whn0yJxGclEu0CJ1Ni
xWUNpUniiif3uwjvec0tLXHXHxUwTqGB/SmIJBdbUbpXJjhzTFOtppRSiuyXDraACTGZuaBoHKMN
dssynqaYVSyZrSDcWrNNWMOyY26WxzhVR9CJKq9ZPWE4iWxhLbhGaVnmovip5ih8VT1oApmEClPJ
W6VTrc3Opjt78fYAnOwtTWGBeOjvbiXD+ANCxyqRUOxKyzxpsS7n2YbAapUzHQeV7sH3ZqJ33xgS
v1u3oCQ2BrxqiMcYlUmQyTATqPuXV/rzZn3xABfh3kcpZ7LIt8F5seMkYCOYlrBp7LX7+vO6IcP/
Tmm4nTQ/naHiq3X71AeYUI1zfJ5lI/CPbo8Za202f5s3rZxhk+AyjULoVNxanGUC6lFI4kD/qgNs
JhU0vbJWhmM/h2V9vR5UgmeYBtgMHuLvbbwJVfIb7AwW9ppSjwHSNGvd6nS0geF6fD//h9HbDDDm
OcIwVpLwQdEApyz75qZim1KKVva618ajoQzwzQnRBydcEnP1SAa+kXO7byPSS/d9sv4TxeevCS8S
GQu2q1I1HCwOYi0mAkZlI8547pSk8+X8U6RCSJOqMa5TGMhxBVTPWf8bClxYbZ4Ll4VH23n+REWG
bkZE9cmi5DXXtAcsb6Q6Vm0YBkuzumMn8uF7VEW7+qjF4YJzNGPmVCFTKJM8IfJO9Y3QRXTx9YA+
zfjlEWQ6ptBG3z7XsBDQAFTFMLWrkaOZOeHTLE+4ssd37uQAjyuo6mQVxFsBUBCBowrK75JaBGc2
Vv68yTmDYDZHwfU/ov2wvyFJVKCHR/Mxkx2KzFu5UoWjKmFJnQ9uWWd21uaM/OOi7Y+/6MKTG4rh
BU3xq+ASYWHGG9YZBJtQQGpjfRg3o7Bo7ZVK278Qh8z7soPlxCMKeKXvoH1tlF2cgNN0JfW9c3IR
1HznxH8FR27EjVCoFPpWOLLzBofN4bzJE7ZHHZyT0Aeo5EJScjRKm75aTlSjX/Bq9dcqXTv6juWu
TPwuTs4BkaYzJillifhrlTmG4OZgF6LdGIIYmrhs6+iX1UM04FooS4UwFBawxkPKlSVfSeFp5GVP
CDebktmawTMSZUTx6oVVeMNZ7YjXuhIJ3cDDwdBSbvOG7UKplcmZ5214urw+sYaS73Xb0WL2wlYZ
KVtiPkmHK6gBPHzDUuF1vjLMu/EW71XcJdwckx+F6u1/DyLC9AsFltwE6V1e0JyU4NZJaN0b8eOM
NkN2RqCxy0FFJ7CNBlq01PW/LalsuJd+YblsZI7bOf5EMmVgl2CnjPwYj7mtbYrqCAiRPzVIobAi
Rx4G54/R51wD96AJq+lvNuw+ARKIWrow7Ay+PU0IOZwV67i8boKpsz0O+S8ERX0Wp2I59SfUUNv7
rQyaB8uYdDJa9KcrojbtYt6LVX3NIN+bSDnXi6gYNGsG7qTJRdMbEp1Gc3Rd4YAyzJLXWnUPk2uD
3We0I+v+DCpBSwdNRAPwZSyKJYgj2N0eXEmiLiKnzMUTgzI0af0rKWnX6rT0cghU2PR7wuqQNNqJ
zM4vFQLdo+QSJchnSBFPT1q5DGSbDA2jzZsxsDLRO/jmtbQ2V0IB7W7eho0vWrqzq3NnitVAmv86
FLhAzvFxszihxS782YvpsOshLcinxrswhaUh+LF5POt0zBhF3qGI+XVqE+IJ7b12yBy5G7r3eTKn
/7tIufKqSynLh58pOXf5Th3C1U0+QQcWGBh9mrnqFuPOBvsk2PuJqayCWnvqXuvon4U61ibts5gV
R2Nz4m4+5Diz/5Fk/b38jjeWtkHsH1Id+A/omI/aA5ziznYdPdYbNGTC8tNyy8DWRtn0G+5VxC2D
CA0wevzAKa95MfIz6mJ73dW9z1ARXVVyU3BigvQsSuGduL++mKKRIpgtabX1WCdKz3yMIx+P1dOY
4y/Si8vyGowpwxmOd8oNTJaQtlld1hDH6mnSSVLyi6wtMgcNgfOsf/kiozw369iturpv1lgx1uZb
zVW6w//tXyXahOgqH/FbpzvEhc/hj76N61w8ZGC/ho0Shbzu7lniE6wDSeX6oGJWN0vazryNqFU5
SKvzuPufgOm0iSFH55RrimHZ+YAlpbXofo8xmGELq/pf8B1J0SYmwiSjXr+EbexBtJH4eJmrr2Fz
oAfVctETEhf1IB5c7WCX9eoLyVhms/pOLKyGhTqSHeHUFoz/6RlKhBdsxfE1W/R8AoMpr95D2qmJ
ksoTEGwm4p0qzP0S6rFNdgHDom5uBoulrbrv3WzkXM92/OS5Zs5Yj5+g3Ed5UGbZt0hOvGiznZWI
cwWVw7yI9ozyjwiLThG9ZIMq68mIofMTHjPjTC3VkREU0PBtJbXuN0KlpjhA1FHp7AFjLV6/gwpC
0hMIrg5YHR2RNZqZIN/Z2FVeAZfaf4Qo4OjBDRjUhXLqGLXMcgJP6eFjsArrTiYeOlcMAOByTd52
W8tEh98SJJWpjClwXUgMrzl8nGmk1SiBKEZJJvbpfu8k6BjaJB2q7DLfXxMO7NIw0cjN2KtgYRnt
Fl5dBBgaJiYsZvApSB+uILeVbVDjw+Y97mlyMlgdm5I8vqhwthiOnoR+CTBqeC0eXMgGKhlrgmS+
y6Bz4NWYQ4t1NPbbzZnDm7TPa2Fe5Fx1Fh5L3wboTxXxDuh7sr0T8OKP2bACccQYCdfsQ2XjYlL3
IT6ziFrSCzoZLZn7F2UU3rDfnNw6h1EiJ55HnwT0poIaU0+orD+vJ2cH8iHr7iuulds+DM2LB+YI
Rd4YZ0qYkBXzEKIgacudyZqcNgb2/4l2aDFQLbg5LxTNmRaGaHrKy7/Nq0W5JCbLZebOPKJt/ETT
MGN8mxYxkGlTSsxmx59jurD09TQLG4rPIcpUwLVTfc0mXTPmQ3Yzhxuw+CRb1OfafQAEJW46bZLr
YYH32nFGi5x84P0r/IIuFrQ5aLyOkAQJxWfJzOWzO5KV
`protect end_protected

