

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
V1ATaLss3xL+7IB2K7seDA6yi9RitRYz53ag5qdvrQJdCjIFqYUaJId5dVVtHD0DOYcDHABW7hIQ
v8c+Q92fqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JSgxjyegQBWsi5MRQkhMNsKXlZ6aVsW2ub0eFRxWKuDdjpxDskXdFvkkPRW8gfb/7zn3yuR0wSAM
GRXuJE1RwoHwaBtkHWGsaNADdwQwJVtSblDHza1Np/UGohmWNs17KQ0KoaRUseontqKY6qmQdoWc
aBe2jeMSzway6YmBYFE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
okGB6ig6tnImIMifoibsWZF2TZuLPRk5MnlxuXDT8N/UFnb2XGKRllM2NtrttpFYLKaUCZeE/WtN
BCLOFNHvLwo2F0d10U0ixtH3AqSpqBhiwSMn4U9Izi3T4B8Jd+wIosHFUL6by9off8V5fFLlgFM6
cTMYiMb4Pyw22wYEZLLHaJN/PgLb/mvesOoNmqI+uTe6FIw50G/trQFL6HkaeY1UuqiEkC+2rozX
Q1z3Mjr9WnzI+3xk/Ec1BuE8dElSvpwFvJ10vjPO6Vpt5wEywOqf+/vAojVlos5DKq/OWdb71bLO
aZNwi3Dc/tmBefQjd9VY04VZ1rZehiZfi1ZCFQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z80u1aw4Gr6ZmqYa2b/TV0ebH4AlJzaoxz1RaRxAjpASOJ9MQdPchu0mfYKmBjBAeMMa2CK7NyUW
LgNnY+cl7c20qN8VH+9rmIxjwdJbj6dnIZ+IDU985ac7xeV3oikYZQ+KYmIC98Z7QnTnEb4rZZo1
j917qQchgNTxm+HE+5U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a9BikCfoqPGhBJNz1f70Yiyj7X7yquoSa26XNvA4R6IzF2fcnmtk249Dm/vT04PGLbQWDjNHwCq8
AbqMetBSvbFzxnydx0xjkALn8kJMuB/7fwxxdD3xEI7iOv6S/cJ2YQBdEHvChtFHvJLV4WdZXdAX
ycHq7luSjNxqnAdnOwRBLcj9p3YWyTD7Ecu32x9Vr2i4pmCnnm3hhjtBy+vPiMsZRfRF23vDPg1j
71P153vTLFNnf6B+LcEJL/9SuloOpe7tygMRCt7LNn0FvYfaso6IQxcv7ZBFsm38MbuIhfRi5heM
8+dySuuo04y28LTeOegW6ronewu1sDu5rpt85g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
OvTRZs21Ol3k9UnJYKQFXdwIwex4b9bK9U2+fGY2Y+Z5P/btw7RVjoP6h5zKft6QuZWfTSViobYr
LWBIxQ2qAiZcpzbuugX8MNXYZtXbf2HbyNwQ1jm8BScfI+mku62ECsi6DRBpYlAxo0/TYl99lXna
Ukro5tAw2Sa8ZHTlsvOHIMNfl4ejAWh4x7SygoGCkVbEGnwn/mjuZYMtE6JcqinbImvpEm9AX+Or
Y6Yv9aClDtHaIkO8RixH5kjTnGZA9/RvjK22E7ZFH76XnRABOae6qnKR7CNJS6fEw11o9PEE/M+F
y2afpzzpOBeVltV8UmhgAS4dfyUGqKarwrPwqwYNkIbzaCZaRrCxxaua60tKmrtTMHsH7aZIWOu6
aa6YQMdkhudUh1fo2pg7R4f/pSmsAdhKpjBh0ZQ9RhgoCWH7+nSW1xZ7CRJfKbM0DMnSAkALqzJS
aryJXoZO9dVZpK6lnRqNWt1VwB+JuLhqI1E39d44uJIFvSo0M1Y6w3M7BI9+xIdKvVXli/CRETSo
nd0K2zl0C9XEsnos3/17+0wPADvLX94+SJ692DaW2vAJtTsLryJSvuYHI4pGwUb7OPNG2bJI0eW0
HbmA9J9mrRB9CfVuFNVwn2JIqOkDrBsRgiSpc66ZNwNP9OeUaoI97mXkJZE+rMWiy7qrOj5ba/xe
NCzlfj/fvc+I6LdI9ZP/JTexuHso6/AHueQkJowlZOScQql2PYkRSaBAsS8maZGxquCR9LXuLPIQ
rUfKhlaCp4+NRUNveYfJCUqnttng5/LA0E/WnLenCGwb36pMuWjkTvo+ziw9DRTD+PZIaRn4DebC
TFtTVMC0H1pUj5lIwh7/Ao7fsK/jKDsAMBHHrc5hn4e5lmlRd8hyJSCmoQRdE5qENmdb71xrA0ZG
6nIyIyRvqECSEY/8AatkyRBGnBi8mi88QdCbHL9apRq7dPGuqUYYHEVS7sdvgyGSTXHbM+uR3o9U
q9NiuY1qSQ3oy25SaPu6rIASoYOzOIDc+gR+KusSHYGH6q8Eq3ZzLarW9Ycul6lCAyyjCAULyyo8
KKfx2ZIjxguyEDPkTJo2EsLcEVHXO6sbd6MdRTaVa4hsxTkbZDcbZRXmcixUTQHKBHIQOfCwOynN
LUOD6igB9eMb1RGp884I7H/QhZVSNDhS63te+r/m0KRlglW1yHjz8d54Cll9uBpoPKTww/uFk44M
vPWwY/HDzbVMwESwhuQbUlWQpd0fXp6LF84iAqA62qxNqOS1ARBeUhPOYw/0qSllqXXy1W6qmIAR
XoYQdoyRACMMwYcQPFClbYZW0jVtWniJujPmxG+9ldrCFrQ0KvKejdJXQaW12Lp9BnyJxL9nDaTG
uN7nTo6W4ekWBy+ETbq1/BLAaJOiKYgNH+BOecWQ+aE/Tp8PcCPHA54RHiiIqgVQ//hv1y/3OGD5
5Eh2WbDzDf/HM11GrV4spzxZXBoTTj6XPeh011jsDaLRQpWdrdpTT1SbSXvtbqYnC0ZPJ3qVgXqo
WIQRqs7JuEZ9ip8CJZleTUf4Vm6xRus9tglIapllkn3ogsJ/2cffBWFrfIIkIdFCfbZ+acnvLxd1
EdD+LTzCtdbt0pKSfyxd1ueUosYO8Q6po6mIiA7WT9KqKeVBJHJfA47eUF5rxPwbX2bm7drv2J0M
mxOzB3AItxS4QKksCLNGP7RqWABHU9RwtRUIZwyo+MhttpYgewb6iR1S4DXAt/BoFNpwVcqYyB7G
DjqUJMeBsXLXV2dLuoD14VdiArBNvzQiP0kCAAu1c6C9U22QWOnsVtaaF9eKyTi9aK485FV3VAg2
IsHImw27nsrUV3Tb6h4k2KUE41G2KsD8uaKISFDknZpJd+BHFr0E4eQzIg0WAmRY+IV+b6C3phrk
07LEDuT0BrzBnolalENPmqVa350cpsNW7PbKDooPIJrxBY1UM1E+e7cbROihQ6FD7+SkINs2L3Lo
rlDL/MaSdpdKqRCGAS088DhNBbXXOzJpRZjjlhQ3f6+PDqXF8bmjXRvIqYgttbVQrOSD3YXiufMX
yxvoUyQTJgQg70nGOxL3wPGSbPbz4WAwgaCtRvoBf92KiAJhP6HzPXsXZp1csgCxOr/uIxSfah+0
6E1ijRDNYeWnnj+PQjN0pSR5400qzPXSNYCIC01UxJxO0ZNyDhlE7Wg04SRfqsC1Ij3kyLmEmWdb
132H9urrP3aPvkvyKaKkp0C4r93AGBj+CW+Srb6fJx5nTkwQuF+ej8eJlncM3aUbdItK7hpEKl+o
z9c5jofZJI1VQq7V5QvDr8MbP94a7O6b9zs99dT/Xf1cxwCSSqz/OF9MMVcopdX5/hJKIJKa6tpl
LudZJLFXTLw5iYiM1E/BLc3m5dSZZXIeJyqgwIJJNFVi4HcnwXi+6NGja7QVACftxTPObNQGTAYO
MHdaO27QsyQHYvwxOgzjbGY2fxuXhA2F0nv14yml9N+C7frNIek/FsmAf78DtTrAatmRcYarl5l3
cg/V1kpag12uXofgpfsKYsWzAW6/KnAEmidxS4z7SdwWByNW8fRI48EjbndcKjkuRBxGctGFV62N
fvx8nuVxOtLSi29PMEciHK9fRlOKiRezsEa5UD/TRlnIyJ8Ek0UvJwZ3x6giF4xO6KnVkI6DHg3I
ZOwI9N33yMZZfJw90dGig6+TZDFYRtYjAARsZ2baGA7B9wDvUNQr9sm0XxDrssIuPNS3Q30hl3Hx
OL2z4QMIu2467/aoFmlXUncDXHOH1HE1FujlTICZawHBJpizuUNJROBjW4ciYBBPN/9CG4IXTY4Y
gcz5xR3hbeCSwLeW95L/O2NZojBL0wacQZ+YkyNMJciIbtTi7bWKm5gMNom9XbGi9fJAVATRAOxL
sWpKPLXmLI2T+X9ptG4TBoSd8AjmETa4m1ZUuepRikZfln5wrXtEtH23BXPG7mw9TNltd6lUX5vs
By7YKMhgMXiD6z+7G31ieEMoJWeeK0iMSxc8eEn2vSx8Q3Koc2ybAvp+BSoL6su/3ZGSLrotyTWb
ZkoP/0wb3FTHGV6nTK/aRt3nGTnGbb3CmR6oStTm//mewedoUwNbb6ajQ7B/z4VY5GdxI/+bh36e
HPR85P8EkGJR3qr9hRzOcQ6PWOckTZAWSUfy8rE1w0agPJNwA/zu6cVxD9yrBB9kma9Kl9sEQ3X6
WvUIeelgxqvqgPhEqGdCqsxGxxZPK81RlnbWgl8buwEeQOTUogyyj/SKoNg7XYXBFmRFVdsCigvw
qTrbPy14e7BT/m2W3GtkGE4VwcPg4shTLc2Wv74F/6oh4osqAcOSJJWOLE2hfkPHgEcnNbN9iofo
9+Apbp9IAJQq+c0Z5Y8cr4dFQJc+DWKWmBhx/NiH99YEWeV8boxkvP7WKifbNk2OZMu/OkZdrhc0
py+R9kU3hmQsab1870mz0l/QO20HbP9BbP2lA+ngsJkWeIRjhrjbImQPrQ8j9GU3XG8JdFIB4CZg
KD9z4s49eaNY1lEIpibhf6GtVtmE+maZd6hMzkJCsmrOkfUSFPdT0/d5SyAXYCPYU06yCCOWbt3h
x1guQe3xcnirMYoBJdgTaNrxEdeHLg9UGiBnOTjJ+jCWJ+GbsaQ4MXEy8ZOG2ICUnupVgvq9QqP4
MnAL5JcJbPQDEoXrO1a9WJ1s5oZHLOhnMMyzdhSxXoqsyFGQSrOQKaETkynhxBwRjMuxMoNV8KwU
/WqG5q1qVOpvdltxN4LTkNdQs/BSIuytRi/CEm/i9YrAATPSqYOjjDdR+VTtksv2hw1dN6uUcaHm
Wa6zs9aOHrkWGrt8GjnaOT67xkzEE6EZv6GGMUjGI69+Rbnog5IIQWyydVOpOst0WPPa4k3TdRY/
RnKcdANyIRnZD5gwNk0qCa5ceJa4uYafwpbCBPzjqYwnOjQhL2h0Uucu+sdFuHEHKuZIsSEhbpDx
ixrpPO/ZvwRG420HGqLA9FPerpLR5iF9GeWdYsarGHfo1a+WWKk0x/gs7+wME9OhWYgQ76Vbg7cS
BLfpbCWHxeVhjPXu2SjyPL8pk7lL0lgcDNS7LWRQ0uMj3EXqInPiOZG68V5/hP0Vf9pU6Frt/g4l
BnR/qKi/Sn6zMAz4y4FEmE05mC0sttF7SDshnMjEJwBeUltNcTebkk2dqSk4miB0yqIkDnUyts49
f4aK21iJ4olkprqCnj6zzGW8UdrutdsBhBdwAMApX9B2QUflyOrT2n+fDuLIDGgA/PZpb1Ylut+7
RHN51U9aiCoUa3Pbegyvpal3n1/DJbWQrDA6/xPRaaofevihGh5duKpJ4kPAfuYVWB03zwvaEymU
DQFpHf+Xc++SXZ/FVSEHv7uqTNaUreJ5n/ATPu21Rb2eimWbOa1FKGjEMnReUkOi4hx53zurfwmg
f2nxGJy3iN9/+wCZA9HCBR0Xjc8WnYRHnDMA02trLZ+GW1A+8MQGRM+tOC61w38jAePnrOrxEKrq
V15+Fa9oQHhiYD/0+CKWjJ4h6ArvFSRp1yCt6MIsUTitxt7MIS83qDJ6v9zrG1Q3RVD75F/pY9Fi
JjAmcHKyp779z07TgxzjZ3JdrwEJqXpCJqb+aiexd/5Rt2FhUuPo85a2Jj9IWd4IanukzGSVX7so
eYiU+7RXGeTO4AgMTatCzKB6FD8dajL3EgzArqueLxWZ0r1xqu3/EkbHwvG2p42GssW+e9LjbjaU
1/ObC4Cm0ezqf8GDoGUeSnQGEpRNENys1fEywjAcLvUiDsT4EMJ8DTYEajNH4Ot7BrshgMEQVuav
B+p+X1WiiZjT8JFUMxIv35K3SQf8XWW6P0OskAfg314vEzpsnjiDnttS/fjEBeE1fO6Td5NmKGwi
8OQ0UDb4/jgG/MlES8edTF3tBp3FGKRWdvyQ8af9LdYakd2MEOLGQyvM4UJ2x4Q2CmRF4Jiyrukp
O8yUarui+gTILeinaFxIehWI0haCeWLTm2dP4WSdZe1vE0WH5+Bl4K8UogwyYVmszb1EhNlctoAj
enPIESWYcIUQ1Btl0PXgHFo94+CEaorOeRiM1KZm6o0esUoMZXt/988/aTf8TKZHZtPnC2Z6pL1D
L3NfVX+bADTgWz8xdQcjKCqJIxUbf6jBG+hou37joE90zYBRkWJYpLgwoa9S242TXIcriHj+5zoY
SmkLv1HRT9oROjDoBxoVZRzy5U7dvhblqFDEk/VTQ6QgFURxEGZNzShTM9TJrVmp0AtKE9nIgsrP
zCL91aRCOXQm/Ai8xqe3oCNzczqUwwweulfESqz+uEpEStB7zUQji0ZZi03hjgKVZGc0SR6n/GxO
83NfnG7GPTv6VRszPAtZZlngQAf0TKt1R/uMuydR0JDlGFIpK8wrXACZwc8cswfOkqpOVeVgM+kr
KcwbdgRLnjwP9wiWDWErmieINvGIRBYBOob93qhBAjHqzHhUUxrnaHBZUlBvT1wzdqy5ww1bSwb0
IZ+601Dd4mPLG0aGk0IeGwfpdmaLpR7H0OVyqtSh6+IzQRC277zi6Nn9lxWILK7T+3B2afTpFyiE
2K9N17zm3TshK/2JDlDrFifDro7BxIrUTliO2JJny70uxxVHZO9+mcMaBU3xk27BQiujC3xtjAOI
Y1UXkqKf/oUYShCqmH9k5wcVjGzKsewi/jgNf1n3H2TfiM9euvE=
`protect end_protected

