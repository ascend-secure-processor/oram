

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BSkF65GdOG5C/IG7S5h9qJkTpr4S1O9NFBkBoFz9KnPnF5zlLHHvk9+acdCXqn61zdPgtM3neM/R
xlsm56NKmQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W3ub6sXXB/XS64utLFH98I9kt3lhmYvY62d5CWUum5jh5hQ2DvlFJ0a3LzIH6uiX3VU6i38R7EVs
7MvVsf87pegCz7myAW7w2y6GhcPahua+82UHaI9gYrtmp7Yb2zGDPygbZjPlFZ90ut30OELil/zp
iGDt/M0M/m+UnyEiESs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PdT1tmlMmHBd4z0vHntNcDQ9q719Wtgyt3SjYA7yz83OZ9IB99rMcCxtbubgo8uBqfEY/jpZJsqy
vs9fPI8ZaeceRG0mtOVGuBGvkFcj7mfnEBI12CT7NhmTLtW4RicWkMCyC98L/Zy4s6EylAC7AHhi
DrZ7o0XKBUVTCSzpVe1115VQM3P70KE9yg+SkGmu0K/T3IKWbrm1DJLQvUD/XeriGua5nRojPt+k
9qkmXgQlTttV6GoCb3kaIVOwXQdLQ2NAF/lvDmmk1kgtQwtq8PdhU3NNRMjJXBAB7C72AdVG1Ecj
+7NKzxx+Of9qsagPnzJuovU+4yHuuKjlCKbDxw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AGoi11uSamOx2qkJmE0N6cTuBhyRtwX4G0L1NRSHrm4OsktOI9nfLSf2WHzeo2dB/0yrFLOG1AgQ
mxalwTjJ7g57Tqenq116PiZPOoyNDt4W5H6w8CGw1sxgYr+fzJT+LICMaDnw2UhahXFTlP1u6ScF
i1CUQIBBpCLJCMAiO0A=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GmIZnHrvWX/hzz2oOz7TqrOLaznLLvFJRGLtULISlnUrQV9TzDFlLrII78YfDSu6Tr5GEUK2D1UV
wZYxl8826gj0g8Y08SMMEe6Vv64STK9Gn2btv+QOPOibed4PwOczQPcuJMwB8YcWkEwC1RssO8fE
L8nD7Y/Fvyl5r2hx3W1xU3un7z/WINHOQlgpEBI3rKo6Ksylfm4pI/ox3uW/r9f72booec7lgDIP
HqBQjQl8ugVoozpeeiChIjer/ftdWB1IFSVutZ61rEVj24U2kQPLDGG/jPIGBO9ojLAvHC4A6V20
90sk6G6LXnpc8Eic9EyIeRR5rKgo5pEnFLr8xQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6224)
`protect data_block
qDsMofjGxrrLyp6H0kWPky2zCG6MmsrhZov4HUkjOmcNOiSimOD+5DuwmJBZ/isdsipxPfm+KLVQ
eGu2KSIVlLG9u/EBbxEFo2JuwH4B8f8NcCOWeRG7GkPloFSvjvwhzUQxgQubDbwSCIcavONIsYAU
rsvzY7DLAoVs/JL+T5PA3SwaapSDwiT3iNQ6OOSB47DHm8Lzrr3vmUZ+ecn7qILlgzJ4rcegMM+s
t9suw+Yr5nllJhsAUDGlojh1s+R87uhKkJYzWJXvzwt9C6tpj7HXFf0l3R4/m6IhuYBLy78NDBj1
cP8MpNMUOM09yJWuVvMIV5H71IAjATLQPxBTVhE7b7vJ/hipeqZHls57rQdtXGKf3zMWkrC9GDaD
+LAwsq9nCFCeRJ7mfl5eb8oqxVZcQkGCVIiBoqJtrTPRZGGeZbmQNi7gDrtPWKvZbXU9lM+ZCI8b
/bZKPeXi2wjWmPlfTbIuQ6wErfXLR1QnvPZMwScx4fAzTLWwD+IajBdKQqSUOhDNX0qSPpO9Y5HN
JUUfzJg/q0Rr9gPezTmIdH39x7XEh6LoB8hooHcVVFlV4WR0s/4AoFiXySS/n5+5fqPtTQwdVXPg
sThAzy8IpgrgnF6tzDT38xo0FZGGGoC1UKGsDNujcN8pQ7Ph13OXEmV3Pwssq02J2xNkbyfaT4rl
yzgnuwxziqtPsp9OQ5ano4WNNTOt5gTFmCQc9U3qkZLm+VefK4YpHGYKmgravDfpETE9ZJCTmuvk
zjr2Yrq6HRGsoIoFuCat4taW4U/L4kVrSBPKe74iCmgm486Pj6bPBisCYv4C4pAaB4Q5ibkzy/cI
3Hwgqo/VRAHu4j20po9wyWk6OxvZHOVQg2iKAZQXtSk7EfHj17Nx0m0uLGeD0jM3mzToGZ4na+v/
2bVD+YDWiaeq61EDd1/SzPJbFPdyfCFSku1sl7l3s6WncT3mApSUz+xj55WBBldZ8O2Rt40M5lzW
057TQDrLOE4UpFkagqtjBrziWXghlJs3QcGw1eIhCdFE94DhhWFVaUXlIY2MS54mlo74iZtYlgyh
m0TRP9rOBFRccuZssCMzreMExJvYiKmajP5Jrj02UU5TZhxketiY7Pq455Q8S/wQHibjRM2zH/IX
JI3fNDoMFHLBVIyFpr79SPwQ6MmIurIGEpoPhbyyFG1qx1xfZrpRPWEFDMdKRkWjASb6SSpcNKJj
n8+nsVXu9Dci/AlqG5QPe0sYmcgIMYCUjXuUJKLlDB1qk+tPEIr5toMfXNs69stoaMwMMxol92o3
qS/vatI9/LWxCVyexvgsZ4L8Gl34qD7Bc1RY+af0QFG6AUwtlWzHnPM9/oyUqPjksbAF5i/0Nwm2
SZBbmqolib5hoFg/scAVCXggQpG9qde5kGxFm62N1lKRQu2c09+ARvbBqEzUvfPWmsBaRlULnykT
MOiZPMNlDszJ5QPJLdn1B4VR1VmugTpx9sArvY2wq3U9hpbLjfUBoTGeCWeNlA//fa3PI/Kul46t
w6h5r9v7OescB1K54SfoUE28nGN6mCyfEAyLoqokaMc78G/Mjx9V9DZKB+JQgZVzlpAXIsfw94FD
Lxdykq1RwIdQ2HxRS8Rcpsi70IT3tbE1L8cB4RLfqLNQ7kt6C2C45hZtMQbeuynp/BkIW0Y78ekH
ee8r/7yjU2NGOv4VjH8/YcBIAOmU6vcUUVRfwtPI/d6haK+uo28PAhpqc358jx0bPb+oWOnWXua7
UGjiZydZR+iEylrcnVPWTkOxyWZ1ivf3EJpBHU4X2Lm5VtnEK6M65LcFCm2+DLGDbpatbLAk+LIw
2kE01w6H2v2NKCMRi4SmsD6MZ/G1XYXF17zOWId4me+sfxngddQ007NiRsVsEL1nMNy8TnRTPuCm
KMk+jwalLTrwIas8zxzmCYmcGcEYYZrW00ssbyt31NTP8vK8mPP+Qpc0xNL4WIfSSuFlmCX89uYw
Ni5/k4qXZyAyu8n7VTVfjg3DR4X7yvBPx91PYm09s25ord/HGXHGwZRveTl0OXNwZ4Oy0NNn1OUS
wDpr4F9/yFm6sIYID8lF1hlxtM8i62tUTIAa7CkShx5EwLgM76qHiILR38s+4cqkMMVmlF/2mDHu
sE+Fk1bl8irv8M72gGQxGe7tXr3MW15QA+s4VtBcJbEBA2LNOwEQdlstRKguZ2CTipBklCD1TW8u
szfvjy6s9aT3Cjsa5Zix5eT5MoqSSjQQlNAeqBzawWtFw5K/gZbYN3eMJxswlA9nVgfp9iBfVtl7
Z0nAmMHocakuaUm1aMJE0+k0sJjSndtz3fuHDt4sQPz/UtNnEHzn/4fOu6y6V6RumEUbVHauu1W8
f7m3xFusdvrtcI7bioMcQWs9l1ddG7+8hGoY6oKYO94iP1pfO4johR2ohen6DNugx1na/0mF6EHq
kNxBLxuJf8ag4ZpJbrebWGAhS0CvSlCKauau2i3YPsij+WTPU0HuZyFLWhdhPw+ln3TbfnNREiCQ
jKou4MwB6zkEvDeAZy+0tm2j1XyR62aY/rfLXDRXVty07TJiNpU0Zr7FEGdMC+qWlGIHQwNyXuLn
4AHrxiPvsgzeEUtFT9nteC6ivMGWDrpXtrFjxORxZP9dTGsWfJ+NrPZIFgB78PVXIxQYCiRX4KSB
Nv9qwLjfOjKV55mhWcB4v21DUFqk6I43V17BDbcbtg28j1rbaUWB8SXmYttu8B2N5GHvEc9cRHBw
5feh6T46pS9lIMcC1/6LvelQXYsprizxGqKDM0njE9BLqsg5ZmqjpzBp0E2SZKXW1e3+c5dSvM6O
jDABh1/fFE4AtVOm9FH/hqjDA95R32VKEFaAFaGu43ZyE+iFWMKsDO93L6dBziSx32avjUOSkwl9
AzZwPTGerwfEfCICLO6o32lR7l3Beu7umCOHRNKozJwsVK/Ooz0Iz43ycu7wE+HcvFSiz9A+b3P+
u+zlTVCHNltE8oAcqA+DJbguwLUqvJRKANcuZeYEMWyAq45S49DizVupMz1+0qnjfYVgaNVAnoe4
nfnx2jrmbHBY024q9XCOAHQgmrGTyL0R9o9tzYj7azW1Cg1rIOT/vH3oaQZyIOlHyhJL2AF+csxR
CcxaoG4R8Zq9PRVFLRVp8JZ+uvO/MfcjrhI7enR9JALC3B3bBE4aUZ807xPgfCHHcCtuE/kIuDEX
oD1Ucqn9BC18KGydqp64p//H662eYZtcah35J93uB+jqzxYEv+haee9GnKYd/TgNQe5pG6apH+FB
MGRXR33NcHeERNxNc2kD3fFElllLb5c56EeJxvkFcvHg/JcNkPn7pJxUA1a+voVZNj82OM4iJuIc
nnHmBK0P551ebW36tuZ7gyvj1qFkNcMgGE1/tbFHQWRKb/m8AXJedkqqhuBcQINQ84PBnBk3Vtd1
72lWeRYA3RJaKZFU4JHiNeyxs9PK4AVHuxKp3n7FY2LPbQUxJzM1RERkCOctr55lDSL/6XM5VB52
VcgrouxwPpkQZTEhx67i1CISUY2gAH4sGzKtYypQ3NRYKL5Fbz+uKas4BpUL/9e4yNTP8nlzuXiL
dnfQ98PmNkcOfxRkwjQLTiUGAuVMFXR8YDaVOMzbC3OqtE0ncWfxMl2akuMevWxFGjMHlR2NMPpI
Nag/Zu5YURCA4wpuXTz2cRNZVm7+vEJMO+CM4i+p0XGRDtyq81eHKjWfK/m3Ff8FrRwfRZFzeB2a
7cnKJMPKcpix8eZH+KM/BWPQxLVotnAQRN4rL8ub7uaXdElXI+eivD310/QehgzuPgNcWJmn0Rrn
a5khrO9hfC9vONNzQkx0yHHRq3aSS4r/dC00+yp5KIub2drP+orREFF1ExjRWSNVc9Flj2DmFzkg
hI36PMNMhAtMQyVOcr/utSHl1og/WLAlllVsOeFlZy4w+gUzu+CECNIn66wM9quHpRlzCc7TEEDy
YqwPNG1jGVZGTbbc5ZLCAvmjjyTwfWY3nI0AtAzR5oxE/ijfj8qvT7L3NMsQ1wN30WdY01yl4/tO
MYwMuZbu9150/yYtLFAXkDPwfvj81zxe3RPAvTQwrYNUt7auL9g6gYEv8pMDHyKUB9jXjbshH0Z9
zWttfEIjTgFUUaSxqhCVGSAo0JxZxD/0ksLtFrYzbgC/MPckJRFUMeJZNP3enVCmD2pCYSBf97py
9ZaB9se1bMc6hZNAkgFtMKrcoJkihA8pbJZ9VAzWc1BRvQzS0BCl+nP1WY2aHNUJK1+VS5DA/udk
jGSeMhQCYAa2osvNmXaJzm2OjUIFiBzCjFCWTrsdyFSjrnF9T35x8jtR2fMzOCyTDSF1yxBchV/4
8lPMClLgd29SRazZlQ0fVVeJGN4YVVbOGdgv/MohUFpMz3JXy/sPwARVMifAkAIxK7EZq/+ZAP25
rmi4cqsf0OSFMWLjCX7KJRxhEDEU1elUmcI1rreQMNFZwIYjGtjHtGVgaLiCWBdsshoaMKIxymyv
kOKpwyH03O+K96cR1HiRe41VV7XWdat4EFDJHWb3QXoIy8hi6rFaH1/pP7VsSj+GQgR4fBc39uTP
zm3A6uaNjG/MrdPSTqbECPAHLs+MyrmNjR4XvE9/wtT+hSQOTnTJD3ymrD0i3MsiPKCw2NGSzeAA
7hMUV7xsLi5v8vwyFIO4YxFXQHirLwcdP/zGBYt6qXMKwlOCCBFQFatnfDg3RLtG2mR6GusTXJqC
zsCUvo3YCmgaSnvIE2x8/2kfdiMVONLsD0yOqqRiU2+/j5DIC9mndnUrl9u80oUHsAJDe3EMM5El
JoYIo55p7iHGyMhgFUYK+LErn2Z1a9OhqkoAeLiDmEqjseX8Jcn51QLlbDNGa6cleGDrVosi+UWD
8JNeJFoWaiT2lgSy+HZVQ9QUaRSgXXkMZSt73Yrfmimwsmcb+u37KNqr8CiiulKuzmwl4Is3YG72
G8G3bXMR1G+i4UwkiWsd+yDrSiRQd7tnKlSbmXsilCPsFVldJlccxVgUe0KubmrvX2KnLa/vI0X7
1wtuZb3KkSMT3IYxFGhZ4LTLtLNFKOx56YzTBn4LqwXp1MhadPAfcWC9GZxAXvaV3cv/Vfpmsjau
Urf0a5562ICPSSicACfkDbiLAM0xYt9LDZGv+UfIn4ftswKzuQ7ed0kFjU3XvaubO4CpgcRT1Hww
rXmy4dOXCcj+AkkMKVHayoMaFhXUdhBeC4w6mOglbidsu9/vQKeYO0/Yi6XAOmrqkzKyNO4prqIg
M0KBdnxdzN9iQROMoOg5oGQqlkUoBJcXQOSqk0X1VyZEbshC8lHzEjudfOVF3d5gSRFeRqbZryn0
+KW+c8lgqEjSAmIJUm5UNWUUHqshYszHcyQ/2G6l3HrChqa/oFx4yxMoM9PAADUwn9YEGHI92p3j
7bgAnCJ24xe5658mkpbt2A/lvn1Dmq/k9qQJr7kIrINR7VxwFMOOp5B6lVtG+rBEUcpXvH5x0Kw1
C4sb/uUYsGPL/erz+CtZCDb0mvhBAnL3dmDxXCgBoQv4U1V3k5g8w2gluLrQODIY5k/a/zCGWFB9
AjYfSPNNDv88XRf9bvlkqcEPVdm30ccgvPzdL4WTSwcb25g2HbOKbxjVWTVFPcH5RyR6Uk8ZNWXd
Br2VQPZsrob1ImLnlPzHYF+IAcW1K15KiQCe92MFUSHN7IX/Sc8g9LfHUqSkpM0P6DdRqWtd+tKT
xqZDT+0If/01o0Dv3+c1l+DdwW4ixhZnmBUrh1MLeC7a5Yuaoh1b+/RfNfWcIVpIM6iYG9JOnjaW
GWHAUxBdAmmmuLETMZz3flSrDDdFW+hAe3ULrGd5zcMwdhMEIUNRigxU9GMXa6jcMu8KMW92YW+r
LOw2KOveFW0befTKc43ic7fc0iqegaCvNuxqCA6FQIVXk05KWsPAUn4nsdTJeXGS1kOoL2Z6eTNI
9Rq602nKkgE0MzEDQnMggLohY/ES6RknUImGrlSwPiGBmxudX+3pvo/pYH4+YXBACRAqiiayMmkC
Iajz4mQpPB27Pda/+yYEcYodyM7jhUo+GPpuGHj+6vmKBLw3k4jT7Ge2w+c6qSebGckMtibALOrX
+TUjJOzPjcsuMX8i2PQBbv4u9nS8jos5xdYAuLS/7yZ15GlwsTDgLxtfN9RBOWbgchSz4nxPnfWh
7WHIOuukMwfdK5PIPe2nNO7JzVQRt5eE6+dUEptOSqyU9lRcma0a6DQ1VcIsthYdnhqg09itqk3B
vODo8x+6GUKh+mCeHacq4ZVJ1zhktwNshw+EbxTK2mJvgdgaplteSWEPPAZQyHx/vm7VuaYPDVoW
qCJYM3Wby5P8vFsxXp7Vk4SaV+U9FBGOmMVP+wbeKVjSHaQLaX/EVyS08jh/V4a24vT002JO1pKB
sagpMAdq7QR7358HQnM4FX8GnAIyx5XCquoOa9RRM0AR9tSHoNhC8VdWvwcu8rpiTaSSPj65YKJJ
AapXBEqTvjqHAelMQk4+Icpc1PtOOEnxGhpjI9pv7wufQgFpwavVopZaEwKAxP3qSFdzEwvQXl0w
/ypLCVu+vr/eSnfbbgnVDSIB+tgf0/vhtoGyCSjzhRkfOi/bnTFfrN/Wad0zM0xBfyzP5kmMdT02
JAqZc8SUpMFFyUerPGLRbiRfsvqdzEWEGFsdaoxvnJOqkkBAsyZvOIftmnIpF/VX0FQDYQImLZq0
lsup/iaI5pX79nV8MuX4mnjwwhrnl2a3RobDS5AUIQG4BBjMoV1ExYct5K4q4Yy8UOCwHeX3da5Q
mAy8Sokyt+yvBRhwGs1sYiN+UDHXzP6zytMvjzxbEsiBYXt40NMOXzaePH8r6l5WQTmT4maem5TR
BW4jG+lu0pId+jv0bBrovXeUWAsfhJ3Bgc52AMpWfhTvTa6jmOVbK2EJrrfWqDBZDnsC1gq6XmKU
iIpZwM4GQqFeD0ae1MMcglbPYnzgLv7xI1TKoB8wK5o4iNNHB+lhvTnyF3y9yp+Jsf65Yw5AEQIm
8XwJucwHNP4c8qvmzIo3d+grbVU1loE2XtuBNxe0f2IiR4iz+4uPWYxxbByua7Wyg9FznaWitd7Z
a/Xt0LOhbRpDos1gTfCgZ9qx6pd3O/UzapW5QIB/4SHrkhK42OdHer1AHS1yiOJIXff0Dqu7u8+H
VSfLHMyfz7f6P9SxZ2IIGgOKmvtVRRctgZKU4qkT0gdCW2DI4RnyC0pgv0arEyR0RXVC916n1l58
AWa9jdOHY91LKkWT8hQaK548Da1oC8nGU1/II9ZPMQcZwV4KxLLIcBFBn3UM/9ChQbFZccy1dynm
1GsC0CXWbvaGxvSflOOQF+qBmW+8gY5ng/bWUUUP5CMx7gwXXj/SRKDKutjNtVvsDpBkVfMFuTQs
NTspBzJd3BRJcSLnaR4VbZDe5S1vFSEk473+gX6yyTliYrWX34+FnoUIrhfXpc2E/k8AEr2UJWzS
esH56gMvaMbcgo5GHUSvNzxbYYiBr1mc+38bQ9aDdOmdQ0Sp8HxV3XOtt9EsAVRpSJmz1odESa/E
NNmlrowHRQFzy7NJppObtuVdwCpzcmoLCXPKp7VUymvyxcD7wf8JAjRfe8MrxmwTeAGm4EmFrC92
L6cNPsGxl0n1Xn+kXQcqIqC2ni2QyD6SknYJEVUFAU+BlT2wJA4Boj0qnoqZRpCIhIlKSZpMn4NA
wZwV+9Wt8zja0wY3qqdUIMshhm7P+zb+bXFP5Y0GT0LfzmdNSvOM8248hthMVplwz89I4rI4fksR
hQ7mxkbALCaTIiGrhYDKpHBCGHfggrvnAEiQNjA0hMSb+7pu/5iVZAj+u7S8IvAghkkCiyLfj+xQ
ODe0kICTgD8Bb++GP3eJTfRxd5CIbv8LU8NEYp/8hwyJ5X+BAWG0ash1+nxR80CfMEteXvt0kwMX
a4Lc1R5uypBXerng5BPAW9F08NLULxUUXngp1bfYDfjQBNAIFeSOqaE0pJ+iSdImhfTwrgaV5+6v
7c6mOjPYqzRsnSJbfyEjL1pxKMzwszMtE9vl98JeoIlPOAwK/OhpwTvC+vwjzm05048KreyUGMvd
HIhPLrhEOy3EhNxjiegv3dxcNeSucmCayIxZW1/KKrEcxGFvb6pB6XYuexHLCeMDvM2TuxhlHq9q
Qyq4fjUetqI8NR78D29zn20gssX4tAfbJOpJoobHk2pQa4WKHz8LYEuPFAQdY+re1MycVLn4jBxI
RT0kJst84sTFm0ca0E4PlYJXoKgypg/auu+XS1pdjubHBPU9eImc6pZHLB8acYQ3WbT0gEJsw8A6
gauL4uo5kWlSh6g=
`protect end_protected

