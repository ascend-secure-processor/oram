	parameter		NumValidBlock = 	8192,
					Recursion = 		3;
	parameter		EnablePLB = 		1,
					PLBCapacity = 		1024;     // in bits
