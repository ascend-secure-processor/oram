    parameter   LeafWidth = 32,         // in bits       
                PLBCapacity = 2048     // in bits