

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mPawqQN/gOXDU6zsccAj1aq4BYEYxxFhhUjJlaBJdStaOlhyZuVZrjwTcwY9QcaxvA8HcIQXSqkl
FxudgfY5xw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ETO4Bu3DwYASF+yGQINNl1qR7RnR/rkfwvmAKfpwUNFt5HDnBDWM/qbvRHphZJnkBDCyGNPNlq4m
itKKKWIGpFGTPVS/BQX6T/QMxnZ2Up4MlL7B7VbSW0XTCCOKl3JOmnLXGH82Ct5vYp//Fkrrr/qt
AmvtDtBVHJT/x317EJw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UkX2abocOLxRHcp3+Z3snkW1y9wMnFsg+IRzmJ0gnXb33/0CVy9VZ8xERv75IzpYHqsSXfAPmzdB
Z8T/P8VGEk8pp56YZAbkHHYBHFcDDbkxj+T8vz+7w+cn5uLx7mEF6NlAf9AzNbCOpKw3b+5CPP2R
LkGtZqJi+lDUWOMX84t5KH/ciZKZGjrcPkfvwsUt7a9lDM7FlZGRxdWZlZRRCCHpV2kYO7bPmAan
NRyyAjUyt+OC2KUuPUOaog6olO+2+RhFvxATLwSZUDX85KuhZk+0tQU7H5PalsCpA0u0NZhyYie7
CAq7t4EYNztRScDN9hDfskVaFZ/oTe1Vf0jY+w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BRP2eOyzP18kec1HWRKxP+ua/ur33aSCVB4d/3J3rmC1wybbXUr6nO29V920cHKI6pcERdpv//Q7
Obd44HjxdaEelav+xhkEi1Ao6pW/5XifnwHDBUEVhL3+xa6luZSm/glkhwMKboEfvIDKVtWIfrvI
9bo33qN+yGuHmLW/jMc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kuAQo83f1lgB2uaOfyuoMm4YzO2rWag41Xnn/92Zw90SlVirQIlCh29sfdCpiOl9AMo1Vq44oCmo
oJBaUCEMDgivL6SB9QHc1h1pLJ4KpEN9mnU8GMbvb2WjFSxkBuGeoAYT1+RUJegRdjom3P409pq1
6t1Hln41j0ZzFxQFOaQLehk6MP9bxQFJLnLGxsher5tIi1+Oxunti1AU1YAWnGdvGDiw25feCRhH
reN2I+DzHG8pA6xvaLPVCHKmBpRvWOs3xBeN7RMdTeNGSoW3QchRU/wgUR+vNVPu9YFBBKvwd5wL
5Wc0HOaAw4OQMphosl+RcdDWEHDWX896yX+Q5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132448)
`protect data_block
9UXPv8y0uteaI8D47Bub5N4yn8O8tOEwJOCnNfXpRfSvyYir7HO71JaCFGYLSPCu4aNIPXcsxPyM
vNh1B41NA6iIPIQzrz0OUasZo/fAQgrMEqgYqmoaGEiFO7YffxwsEeXk39j9oA4+UX84M030ESXX
2ewEkLFsJsK+4N4HKOm+RZwBOTejZgArLhNhqTft9RRNN04n+zXuG0ovOIFy1ZotUzmzRJgn14Tg
ArLNEPkrjE7yWHzGpDCpVNUoW4YDMfHdAiPA/8K8Cl36TnN5bmdyHo+s8voLPm78YXZnP8M9mxJG
ZcNjQ0tfrgYHB1KM/S6lPlvTNjDYecRMqRUgU1yWdWpq3KIfM4pTW+UuMagWV2+5Nei83nuAIYUp
gpRPjQjNxjqgW1L7idWtwAUUhnhCU9M1ANGPy6rjXd/9JsOkRYdy+Kh9CWfJYgXeA5naLlgAhZjV
mkxkTJZM+iH4DxeJlOYM6PH36YfdpkLE5IjJ8SNb9O1egorx1fCUb5Z3YVNEDXwMquB9R5z6DIIe
9Q3hwCbANpzE/7ZY9lGrSdosE0JadSZa7X5rPB1sxnp0ZQVLVCnFyvTww8pa/b+cHiXlPrlKXj0S
IajPxco7hhXTR/B80hlgArewx7+0+d/G19RZdKDvzSuSkDZuh2XOqXXxwm1sPky3REyjdCz+9dBW
fzbXhnmpVuGZQwaXfCPqabMhfmIzsVOifhYrjoY2SIqQBAyMWHvON6wViKG/OP+08ig+xLRojft7
TC8SGB5XFxGEVKj3AF74vwgyDJpn4Arq0Vwy5uaEXTxB9+HfCckhKSs9QO6/YSFBZfDKETJxGEhZ
aDNKsGJVcqS3WXtkMatNNCbYl7ihgFa4mqaRUMqZbqjx8JHUZs+wHQPY2xRIGe/MEd6HY8Avi9XL
eR9kZxuT/oV0DNqPhnPUMicqeIvFZfffOp8T0vCW4cDZoF3pPgAFfKab4pX24Z9oAawwgiROR5n/
pQOEZLo7ZxBuwzWcxW1figKg/WW/zopZ8YQ0BfB9XYpQFMKeJ6KeynARSdhPGQpvZvqLlvHabmAR
u/FrwESZLXborOzDJCmSw4PRWbU23MF7axxVjyP8PhrTdcBer8uRpz7r1EpaOvG/k0HOEnnLXRoA
G6zuJpDFDoYe0KguqUM+EPVvsXgi/wtEwOiflyQ61dlNPs97MWzwovOndX6kx1sQ8du0o9EzxC7a
7vyGq7LL6nsGY1P0W2Fa86BnKZ6VNahlS6DWKeGloo3mtJ3hVgE8SlDyL4pPSV2PU2zWMKBlcJdu
XSLFxDy586L2zjlVtfOD99RDY9yBznZJGu94jm2p011iNYb2u2ug5ksI+VNmOdvQ0GNOT6YX3V32
UANxUpQaHQDnzCOhQ1le+lclhcquRJPs8oG8J7aVqamO5HYVBLqjS0dRxmYf4DO1+tmgMCweSoL/
0NvYS9luYBgWeaSgumow3AqT8Ijqwf4yh1yoPV1nZ+hrpo56OcuXPWm2f1rPhFq0mDAPNUEZCTtF
7GIS4HVEnJ/qlzoYp9ePBiOlHaolx8JIe+EHNGz7bwoN4MKPUX/AQwYtdhQLrMrofRStAXeyHesm
vCZdlTv0aFWfdg3/vzrAV9uaRJPryIuyD3XlstzwZymuF9xdUmOGPy9qsWAMAhuYt5QRpDXaIJyB
tlMgOQEZPekzF30kDVrYYwbP4DHNTFNvrhwDgrmeBPd0DwQUhzop8Pb7D2uoQt82yypKiusLzP8n
Ogh/vUSFcEk7t26v8nvuF58Dqv9dp0aoEDHW3OnOeGKY/+jHhExf2IIMQEP1DirgnFO3u1Ztdo1H
6HkwK5K48Yx8nAIclAjcSLds+O8gpJsFmDuyiLgTeDZCT/xTXKxI2cGeva8L6d7J6+sCYFUz/mX1
gXZ22xpCZTe9Mf4cIMNjX8ifc6z8dc5dN7BBvt5PSDo8neat+h6/vbsp6q4hfx7QG8X7GpTgCR/0
V0xQn6fbOcRLoKAa1aslcVuAHBAvSvOwnpfK8JAOJI38yOwuV0+hDJhpk4Br3NJWLOT3cwU9yZLd
k5YflnZfm25qROWN0yKkS8babZz1Y2zPCQXL5k0ZyVHCen8meSqeWMqHnLtcHye7VbAmoE+6bGWz
rBBKU40Izm+zLhaqL4JVyMd0YKiyQOAq76kOPN3W66W5J9NnATPGD/1PvJExgAHab4uc0xANIitH
U/oOWONhq7+Yy9vP+kfeF5nr4mQU/zXeBs7E7KSEwXNj1KN0dGOeJZlNmE3Y6F18zbxdLHUKdCpd
E8UJRUmUX2TVwQs5GW5gDGQnnEwKUubLAaGHVBFeQnAENXh3vS4Mc+pDBeuFjlAouaphwCk/RYEl
c0c6Nt6L4D3xuTmJMo+d0WF+Hl213eMOcYFUX99d7WWwLqBqlwYJal+Ywn54NfmZM6nrVLMJbUZD
h9voDaefzGGUpI4DcMT29EKLEg+Tt0rE9Su7K7PqP+tHsZBoveKs3OtyG5gCT1GkXJEDwr9wnVAF
3SFJgFrdTEPDArJ9ofC/gF8GaaLvZlgIC62+Q9xqjqgzulXTLRsOehscpNzSX3JEPgN9yaGIUXj1
VQIi9cquyd31C/mVPLM2Ftp1ec8J11LUbwVxFkzasMUVc2AZ92IkyraC9cNTZUkOKNyrS4GXUswu
tFd45bCyM4jfcQ7deZ6TrsaI9lot1BPgHRTFaE4QwnjLgyIfm2xxinns3YFMFQMJaU1SPhJZuxub
YyidQhf1jD7QCfaL5TW0ou72aREq9FpAUMogQZ/zKJTH711sO5AG6zM0u/AC0nG62XFLSjcUMUIg
ahjZ+jZPCRhdYcOZjwULbCZVOQwLxIzYN/a7duj0b+ixkQ526pvAKkHL/JSHeZrg8yYU9xVxImuz
cGsLdzg4N82fp1/rv+SJAPYSt5BbkcNkb/5pY4RMBDxEy7mZmpmTkSCY725VO2+daxdszQFCjNT5
zcYzswhiB2vthRkBi+dq2CeemoSnaIZ5o1p3bTZlUFfI9GslISl3760OSIVAM8ddmEkDmnpAMD/z
Gp75kyxxAQtxiLMAtAH2HWZE7+R9M2vWT9Me7RlvzxBuXbJDzvZd0dErMGrZd9jjxKbCFUZK2GZY
AElwkRaKaYUmbdLCWA2pcZHFSSpG7qPIBEg4tzMq8ckougO8rHACeWzYv3UPiwWOu0Xsd4M/rf4S
vIYiAC6+fyhe+l8Q72LWOoNuiZ2ClOzoCTxRl/IvIE64LjxmNVyf7HbPNIfn2sfSXh5MpnRWIaWx
lGvBWJOQRY+9AUnEpSJjb86C2+BPHi5pYGH2g4ukTtZWxeTym10hba2rcMWs7Cq4G9nj+V65rvmu
q6X3fN0rB64ZqOaZecbPKiKQcJKMd4AWq+WIuwRJijklr3MRRnPO+iWZrySaYlt58OCWlBOh/C0t
aOuaUGWSHuqDCMCwVtV6t9mmGif9mkiRkfJSthFOrpIsZ4i1mLAqbzDeYPEr7/vKWD5+SqvW61dr
Ki9DYRMR5fXKd4JSY5+c9cHlBHNyFMbDxg1OAkQOCoOSRd//wjA6oeHUlU4bwufUN0wpkjjMCfEZ
Cl+RKkFKehC+6uelirJ2JwZxbHahClrZ+cxkslWzUUvMlorOcVrxN18pWgLnfWXI/owiEZDOPucU
NdZlHuVNQxR6aMP+HFFhDSYNWGtHiZdnfgjAUww6jEeAQrVWRn08CPXPPDZANW5vyl8CM27GYeLN
pNV7nPy4jddZlh66pLF+xnBvYU08WxG5g8IFRKkGW1Xgp3/bNEWK1gZzWy8ODWlNK5SK9ksnBSvb
yiJzr+AH3luXkwNj9+pXlWnONSh5TwKxRmAL9HeakeFDQJ/dwAC/hM5+rcdv4PFUDx2pLgQnc8vm
TRGdQGMci/eQC/xHutOk4s0mK/MM1gX3vYEVyIKuONcttBAsWXmS4bfZCpiAXwO6zlDszOKliGbp
9f8LWaA0MQZwChvCVZbXH5u3at8s7rcFcuI1jnK7gyv4SRQ9dpHu+lZOof1Ha++PsaYtrjBY5k7A
ovAJ5mHLufo3XXXjtpyr53/a6Ha2x02wXw6AzZJXOPkyBjWzmQ3Aeg94SSCw2cB+9bdIrOmT3Nc1
XX+/hfWLm9L9QOMn64TQcUHRtT6KLAfEt0cRV6kxdiN3rKlK+6mMvATSS6/FICXx+L2Yt3UgJs0r
CscZ97Kc4j6zVXZEbf2+W53gcMkRGnPaTYwSaSK8ts4d2RZgbel2zo5AoY5dJbrQc8ASP92UIrrz
DWibjwPvTfIJashEm4TxFL6vyz+STS6LJpX9IhTaEyZXjyYz/rscelxQ5r5jI+RMEfUQQhw+dVxD
1jSg/wRztGG7avC+DUAOiYPBjo/yUbTySZ8pKr/wLfGYpcDKrlI6fp7hl5KdHcuH19hCPrMQD5XE
I2mpOJVQptQKjI0vsw1lzno0eXVrhLZwVpj7vsbqimaXz7/O6kMmrgTBNxK5VUFEbH5OZA6AxISK
E2eUdDm0oFnjkvs9g6nYB6rUiuiyhU0KvGJhUv56oXdOuh2wzX3mAWWenHecC1rc4IvyXekicDqn
OI06WFXc1/i+gmAY1cJg/feZN7P2h0jaiUaEQFSm4VRNBNpfHqkqHtb0GMLOykTsg/uitvXZG3VW
T8N4hL0qhKJ9wKd/aubB3vmMRIHGeEV0H34cfrBDP18D+u/XJMM7diA599yJVs2KBuHfe9SV3zuG
jbD/pP2UWGpBdkWccRi0Ar9ZmasRbmPbdkAQSHreFNvcS4Pyn3pEwA6BpC4L7OIcTUVBZwfKdQ5o
9/50fXEcgJ1mED2iwAIw/XasGlWLaSPR1eLjn8EMxGTcD9guwTx85LKnUHbzt1dUDAOwWg+7OPxA
cJlbcIyceMAZXYyhUcLabtjPIh4HvQynA1j0Fy6obtgn6v7iE7iJJZ6CWL4Uo2C0CTKyyOw56hbO
q+0WKlMCZByGXoQdaykTNFR7OdVelwNxB37LrnnVIDlhLnGpA1XyyEs6TbX+qostyCMPsrgH2X5g
v7ucyiEz0hj+2RvL5A+Q06Eyq1A0efiF1RpZXjUD5ei5H+Tg25j5lmJPxi95zSlpCSVqlGVDhMKQ
ATL/HKoxh/YAqHUmIn3rD19wS3EgZLouv00iTNTbSGhRoSSrIKEI5tOLm0hqZui8RfyWxEsYhood
7k9PZeTdmJKxzTdEOLDsjZEwGm5rboD7cdTs9oW9C09+vRTEo9WX1R9vD5zgoCPHocu+7xxoQT8S
g/er4U4fODTCxvdYU52WA2pJ1hZBRjG28iQjJsG60a+RxajHnz2wrsjgEEWatJ8BO8xc795iA9yH
glz/ba6iCDaBozjjdsGVlnRdLWZ6CY7WHpui7HIbZoicHbFX0rpQGsIZSJzfqm5itlWtLnrBWHxN
jXTm4BXjWDq9YFgCk3MJZpu286IHSsIsSvwoUCpwyu1Y9FhDJgqa6YByui9QoQrzQkHvYSEeme37
7np0SDUR2gxidoy3qj3LtMYXy/AUruL77EPBkuu53eNPGbdVJobAn1lHHJrtQXCRCUxnAgpELPem
VAZYuwAIf4yXUv3SIMhJ2cSfJo25xO1CzoyIS2L9/57Mzm8LGpRWOY81TAIE6kmA7NKiWzBC7wzh
KxzQdCJfYuBg0j3huk0NHM/k8Ncl+FE/jQ4T/sCHBOJlg8ExaTLLObZQTiz+I1IZOqAMHrcpgD6G
2didV9EjpCqttji7xj+I64m71spbGC1CbhJ3eLzzPScCL4bYnrhFMfTYDY08KZph+FyzCB/IkTEW
jTZJVFyBzDtPma7tuLfDKIETe25h4DPJbJihJ5PbOWMQ+msCVhtrofeCm2Y1d9DeyG8M+6dzhnMT
bj/SiPwpZaMO0YP6qA+5mhPtJp/9rmNeURoF74AFs/g+aPhYzhyZzVeHKKbIEB2POCbjJNSCqARk
PKMS+SZISdc0aS0L5XrdpCe6MfXfqPTLwY59v8Iq3BkoTvdnGCabXg+pPYlj5aiHpA9v7/UYBdzu
b/5ZVtT5r7w9mPTEUgBskTFkF3ME8zwyF7ee7hhgHRYm3zFVldov+kCJ//3tZ32+JHqkUr2OOotm
X4qR9PqJQeNuXT+AexcB5YaeSEVLZzicf5c8hGP9fJQ0L3QGypenq3Vo6l8vDLM1KwG5U0zNz1sY
p/WDBfoBzrE+Fql2GHGpNQsuS214QCdfLufLlzS5cp9tV4RpzoVO6zX4TcajiaVOAAl35437FYL0
T01yttMpMIlu0INDZplKpDYKptiJhA24+zs8hPrxd/SXaJjW3ZkSlMMayBWgPAhgZAThLdDq3K3T
GrFIdGpyGNCo6SQTKb4OprZ4OyxuX+pi170DQjDC+JAvUayV0MQnFfWI9kuNSWJsqasLYyXQE9P1
KkzMt9i7s/j9pivgdOzctKFKGnEymwzvetxfO+u3u11ZyZ0/F4SOZuKFOsZBKekWv5LJa29UEe77
jkqb2VCHPHeFGxCv0YYl+3b1WRRQvVf8gMSvtn7SXELwn1uCxChPfzFK/TI00j2kMN7La3mHBDRy
uE33kuZqi/XJxAk33RyGJlOj9nQ9K/UDV58taQKX5Jg33Zq5D+3pz4Attq45vu1AYXyvIC0ugcmz
1zyRYZQOipuWcULEiAXaV5tGTqSUKmWRUJJLCUr1oTnoW2Zn66Yw6uVU7KMqNuvNhNHwHihM4Yix
1LytFllncT335Vz67SIRiekiHQb9wUbMHv5LZm3VOBVP5Ovf7wnJvESENvNyrsTe0cvYpplZRtOD
F6HrtoouRKBra161ZSuQLLO/eUYky1t30JhlVt88dhQree9ypi9E0WhRYKHlbTac8vemVjGst3wk
eBXEXX0kMN4rQx8ThhYqSkluRd6DWqncWhBe6YFvjWnGKOi8C67x8wUQbeU6cleV2u5xtj1iCNV2
OjefavgtXB6W3O8CKSAqGniZxM71LFGEJS75OCSeHl0hHQ3o2/QmbKfY1q1qHXBtPIb6kEOoi9ZJ
QxK+XBkktDk09jjGK5eNYmfDEfR+12ks3xB5SWwyvwAnsUXmMEiM2+icVWR7Hw7fGrRZbF7dOXoX
C/c5NP0gWrZgaHlm6aeMHWka/fTpMD06al/SbqUAP6GENMefO7sNqZVdXLKv88HoVDZVndPsBeOJ
howg5jdHcppJEeAUtwkJC1F4YUOsOjnLEuDgKEGVKbyrdj3Luywh1WC5W4HAt8rscxQixoP1kkS+
mJcS74WSzZYlAzx8I79LYU1c8CekTpMj2t5xHCJU38qdJXACJCO1G67J/iHoMGdkxVQsV4YoM57B
RBxCepLnozWXVgtrf1bPcXuH+Pc2tqW9CKhlnmWL/VeVeoGLScBRb6vRZQjirohN/h60TIwOO75t
S6GjQsiAylV4PTzMWIdZ/TH6n7jykMxUz+RehDLiVE5L/2+9n+SR+ehhNMrV5z2JQvo/rY5W/e9L
UH9a5OZ2NqAUahZt4TTI9bZmG19c6In514Vm6BkyVG1oPrz4KaH1k1/dWjuXU3c7mmr5sXJqoSRa
J/jHiW0j++93Pd8wH9poAi4CYjqswmvIWq+Oqpfuri8ZOdfO8CSNMNicjc9NoVdaUT2C2QyMUojm
nJ6bTVow+kJylk0X1flcrAbzIAybr9kQUywcOODKVDSIX3BtzYcB3X2q1jGutJTrGCBhpmri9TKq
PkwpcHbySNwcbIuJSbggttFJxrvw20na/AE4lshpu83FWcbJo7OuCpdt/QcwGomM3g7rf87lZiSo
j/MQg8MrzVQCDcKoqShOaMivcUa8lpjt8z0iOWH1u/XDIbSxAoYc3xCSjGx6WWET66TuU9D3dmpz
M7I2kaHvCYI8zIQwjerAaaD/MCtIOynWTsMYrqSnm/k621yOgqh9oZt2TLpL7IshH3OxXo+kKGOC
Txg+NXQB2aOYD1nC806Nvx+Qm/vklmOJ5EEgSzGkhrD3XpOaLkndAEukFt6j+BjX60NL4Xb99VOR
RHOK44rIeQfCFE8O7xFOjISlUIDpg7nRGhZDIad9tMSWuTFioc0b6e925qtoBY0dHpdMnITRh7gr
vvrMKFEtqyDh+yWAqqYu87uo4iHpz/Ts8DaMdVNoqdf6/SgN2eNcK3iLrp6zE4hjhEfj5DcmXW8B
qu6B0gdV1mQfEbA9iBIfReExjKnN5Uw3IjL5/GeGyEwrr8RfbAEKzyk7ZzIH8J+2dxb9XPmHFifN
HDN2jhR8ZFFHGBn6mPgORtLzPW2RGjAFNFsXKotwK6+cHYZgaZwsL1fpxsMydBEHOT+JC09GzeBH
mTyAZgp3gb3TfJZZAzAYfuDvEAA5+LSZZD8x2crzevtmNADFeSCjgA2YAA52yV9RlMmKYIgPEP2a
QdxdCJSt7bFafTMcoU10HWs4m6YhuC+4IchS/ATTNji54Sazzi2DU2zMT/JHJR/pcabmN+rrJILu
SZ0REaAZUo2febNh3GYbLJL2J5l3DVSDoHjhusMm0M9lrEfIDgkcBe4UtrWzLmNJpFcDB8AHGmwi
WdkfMr/aopR1RWH0u6BCYXUEzq36duwc7LijDPzHs70o+hXJV1bA/xA0Qw1ZTBxwYU/NlTUjB2hl
IfGKbEzgVnZgrfhWiAYSMlYWAUC1nf/IJeGSVT4wtIsZVtX34ZfY37gsUzDihoPMmh8b9MqmG6OM
EoZbp4vbiXMH8ty8HCgWkwK6AU9UaU7YVr9HTAalPQ5+/zHfzyr/hESG+b0GMhYelPzh3vzmqk4n
9DR6HDPwki0bfDAfDdAVr+SbG55BT16JHwmOiySNzciGNHBedkQmC7rm9ibj/IntTcJ1ITTCwGFV
QXIqHsX6W/gsRKKVLB+DITOgLCKjE9Whp2W8/IVaHyywz2ZjQbJLUQ81XhHabqjVTpe9iOJlMKCJ
8QtynrznsW0KcGrjYPKWljt2mqWHTXTXW5W9f37kH/IqrMQhv/61UKWGaAU7EMLKEPBJAYEsoTcI
c57LVqXaBxCM0Vr+E67Z2mabQ0vpnV/dXHepiFiuALiJpRi5BUU71WSU78OmP5CBISY98rOSHMZP
yW1+HeVegIIrNB1EOe6Ie5qUjVu1Lr/k92u2XNCpEGxECtMEAOIRZ0WbIuUUdMhzWhB6FgLl4kNO
oecItFMPn5jK+bemZvVKpxDIRhMceNvy+g/Bipp9kv8NRXJb297JrILeMJIoeYEWKkmuGyPx0bnC
vb+b8dHaqfa81Ai0dqozy0ZOd6rhQeQ4MAP8tLOoCQYH8LG9JFzY4/ZDSlCfan07ShSgw3b8Ebfk
rLhFs1yVWtSHcPrkDiQxg7zIeiixAcu6Pt9vBawJWiAA9cVNlkTzoe8jdcB519qyDdB0VdMB1KqC
gaiTSkDvb+ucik61ttXIqxqHglYzqaRh8/dZqQ152SeBzUiAa9hhf77NDC5A1CJkHIbSWhJuVg8d
pooZoSCzKiZ4S/zohctijjR69hn/5nJ+PMIzA1DKeYvUjmK/bAQuqsLT4VMQIK9K/PrqZUYromv3
5nEoQHZZmMshZ4wcBTa91dTwcZ/gASC4fB30Pb+DaMP1aXdRH2cfTpwdem83RQ3qc5VVLCD5crGA
Br/lDKNE1aTd1iRHQ/WlGIr5I96jo0s8/u2fp3UNcSPF3vSUBohMQidvKOYYtN7/P8o58ziHzf9a
ae6kJcKWnknrJWWCcrWMRZvd55OSYulC4yIc20ejSSN5JnF4KRJAXSGeG1P+sFProEdvHzqBCGmg
BsiMkwk3hI2LH6X4t8eTrQqsgs3yuYNNPNaDI4xc147VIX31JN+pN0dppCTbax3mdmzSb6Dd4o2p
aUuDPh2SzNwbqvo4UnQkXoSQ1elGCwMXRX5rQCLodd1M4SH3F0CQT5/EvUSK4vM52fJHoqgm6Evf
PWA9l0I10LjcC+jERXPm7pg/enxqM84Lx8M0LKj6t+M2SVFrlHEXqUhDVCJJOFFirkmiBOE8VxTq
IjJn94wezFZWmLt5n7vTJESjVKHiu8fW0ivpClRV8Tr/D9OVcdEB+Fu+M3bf32yPS/WYlrJNDshP
6STFraH7qZPsc+zngeOq7VpSGKzg6lBqVA0yAPUKvSbm5d9PN5IuJn6Syo+nyPDyQKSZzwaGg4TD
iQ9L8LA0oW2CPdnJRegRnN+eHvDRgkqgoKzvbwVJuov1ot2Yx9MtkvAF2OuC3q+iGFStlW44XMNp
fmOloycQCaHlz4G5jv78SrYMWKWgnwosJrv1y8Fp2QWokcit/zeuwfOCd6Wess4/A88HZmV5Eftz
wzHNRG7Uso2/zXRXGhUsP/F1DtBWMq2jV5HQLoKuplNa4aYRXMmw2C6jMu9lojCiTMJUkdskiYlR
cD68Vboah6Kej2BwRKH9KlElocau5OKPWD93bmCeXy0vTNTSyVY9010Pf5dvePE7fxlD4dFHVzQz
rsFmS50LHSjCU5m6kk702/FwWxd88qYQHpcDUlPt8vN44nwE/Z8Gpt2AQHO7RLSBAxsQuwjSzUA7
PyCTD0iwMWUdHGO311XIa0h9aq4l6DK1PVKDoyz2+XzFxoeB1vtp3G6xKwKTsG3lht+I4Gh4PXRT
6siz3HapKgJVQeARG9tCf3gP24FBQ+aYKUyI8LqZFgdSnVd/848ZSIELo0Podyx+ASzJzF43OEES
nofSUjmJsYRudu+tvQ3cAoDh/ONHuxZLZFFxsT408nNvgncPLfJsyu7ndNFu5EWU1XXyKG/8GQuI
M4TFfoWlh0wNNZ3D3qHn2bFWompqW3YTiKe5JjK8Dy+sq5DaPwqUeWBapBqCCnVnF9D5wpu9ZhHJ
62bDGyMNDKyQlFy2ISuCsOLVdz5mlwtJ1UO3Q0h3OizdbbHkOt/40+87uodAj9NAWTTgIYErVotD
FuQ58WFLpHP2EPOxcXQ2CirY+DMdsf/19EHMpcSx9NwR9SbhiKJD+8KRZBJMtYiRTSH7wQvRf9tD
0TJzFtPrpJoY6e8FcX4PP0LQaIvJqp4GtF/1W5PmCc14y0gE8tTu9zWkJ5Mj2+W+q0wWhoFzVK5y
sE3ra+1F3DyHjRVhwRLqPGtr0YjqSkt4ALBjQ8qMI3ChST0Q5ewmJKttWJ0O8/GeOHLxPAqS/2/f
Bvy5I5fphL64eTzcS4nqDFNrXRXK0oF1Cn0zZ2biaGTsxFjx3HBHo5paxlbSkILRqPyBT3FlWxm9
0GNCALxt8Pg6gRqA73z+dedupzKFxl0m7jY0SldXIMuxCxAjZlD6lzM0psnfuTbinkQMipGBYTJk
W/6mgpMUT2xeMhsZBeHVGo/14co0SrijBQ4H61LWwJgiUUocPwHkqfSQMi307d9Ujt1YFUaWjrOn
gnwnSMWaqCtZbyGGRL7wz3suNt3CDJRYwoLR67ZiYdcwKoAMj/Xp3zLyjFH8R6/4IytsyNUDM2Cq
as/fRKoyzlwVgZNSjZuwFn2ZD+0wk15DMFBII5lHCRVNoCJ4+V49HV5FFlwxKx8vS9bMpC9p93dE
1+YC92jrLXsqe1Pg2FDZ1OtSnQrh1hTtTgF7/43+pupfsCoe0RBRxDGqwXPS1pvdIJeshlP7mUuY
uO8M6dmr1swju7KADmOJCRl2JZCkLIWJKKv5r8lxihrlV/TfO058YzncNDJvKvlW6+tEJgq5K/wi
uJQnS/iLGcnhJbpAsZ6UW9P1yUoMSuUMLJDeNgBci4HIiCmLandjr77KOP0Klvaqig2o0coup0YD
uWgJYnINECuanaBJVmKux1QvD8hxJG0ZUxqtph68gA9dV9BAhbi5SLoTwd8vu5SdPF+UaIG6INDA
tImRTJZ0rFaFryfIXes+Akc0gNjQK9W6zFgy5Si2w5T4im9Y24+FZ+eiZQ1Fu2bRU6ZKHCHhoBbv
/dJ9q3xBFQfspv9VIXiF02vkN3r/Smb7SNvpgVDkYAglVe5Kr/7X7fJQhyqxajU6t7ZSrCLeHSn0
YDPANA+Ad2Tz6RsGyXVxbGYMRsSqJwGqR9FlYPJBWCGEEzUpVOXmfaEMFAAxxjnym3Zd2QDevWl1
TX9y+i00fQPJLPXrD1CziH35jYaLYW/3nywGHCI1b4JaE0HwVNKt2worSYoy8EIIvh3B9LMUf/fW
6BraCINLBZGf7SlIdRfrbAOS71glInP0oReKqPs8BsXvGwrQLj7P8/WRScUM9HCRcVjEEaf7bIrZ
YT9sAJ2GLLU1xoqTPMMleJCD2sNVQNAAMGYhZaCFiOjEnDQQ4R9RO16ebhO/70guygmMfBsIrZjk
uspKGqhzs4ie17HMevj+N4Mr+QzlB4+Z66XWiqGk2/nLAiLJsNO6Fk3dqg+YYXtL9/V8SU0BAzoJ
4gBQpIB7qw1MQ2Y1NDE0Gu5UR6JaJGc/xDna8XX6aha26niKdhKPEDgQoS2m6ucMCPuBvbvb9ds5
rEkdpf9hVTXT3aIpXvJ/EjcjpXec8IM0Jx7/cfaQrD3MXvNVXbfyrNQBEaPQPI6bYoYfSznT+Yf9
86WqF8s8m1NZlKzx+Tu785NwATvRvgLcKbyQAwKFwhtRaV5GtcvDb6Vdrg2eEejEpdfbKp1YvvZv
Rw+mrUWbLCfECCYQrblBgprnSEC27JwEtD9iitATWSYIEfaO9RUwWMGFrR0m/yBQTHX/QBw5gLaz
DEJqs+zSd+XiiuV/LVPMUxzxKSKUQq9SCFN54cH+lTGYvAwpVFEhyFbX/3hoR5Jpy2h5UrxpT5Z+
1ek7ry6LE7zFX4+AnTsJ3chmiWxCa38fznz3PoZ3uKnAMxAbmaNZfmDY8pLixhBSh89gP398m02g
ak7INCZuDWztZrHA/zH7YL8Hj4wPhdNfLXQKUtc/eGH4hk3omhN4ULdylF1j4KS/6LSR7Ixur6uQ
Qe2zZSPu/mZhCKlDlhvn2UVgcyE0AdbA/piyZpwmL/je68PS+5IU6Njf/AsTa7AqsLd9Bhd5EFRK
tw1AQtCKEAe5Vjy/BgGzHiRv4k2XKvn11NKbCSkbpHCpqgDZFrH7DCSAN/lUSlbBI7ye+0aE8YQF
nyXBsNYcD9NXTLHQBBsdEf6sikt0vA7HgfEcavOzdsWFMZxxDNJAgAFM66CfXgHMbtNCffDKArdC
H0+YYI44Qjyi1DnLQ0vK6zIbpfdbc9MHSAUPfa8kb9c5777HS4hbPRyiKWS9mAVzVx7UPYbcLLFY
yiJFJ5GhGcUNApzG/fF6NqS6tk6vrsZZPGv3G+h1/wnbgJVH5oB743iudTVil/LqwpgIAT0sLvLJ
ENrcf/VPtHJ8h9Wix2uAl4EpA9ztVLVBytfdHzxvtJk+CH80r5/qrb6rkhp29NSerR1pVK739lMC
cbNt87qftwufScen+DsOyXH7JV3YX0bvtU/iTLxUPIqZ/nCNpAFZOoogToBqQqcIyA7IFxehHN1H
AffMOqziVYVdpBr7OOvqlmJtgzP/21qi2mgc+4ncLMKclcLo2Qlbc138el28IjG1KLEgnTxOOdrU
3Bbs/6l1PpzekRpzfMxn10evDZ4UmRHrc6AaFpnPKST5q3vnTi6imxJo9bQjDeEFV8QJKJKfd80F
xLKqyScPHOuwD//KhfcmcOFNFVb9cdRudEYLeAElKJc90ybvvLSOmV+WMTguh8iH9bfspV5k7/a2
7DX9325xrJsnSVDMxFIh3KST8qPZVBAjoCrgHzCmIRx84gtbWrZQ+E6ZXtd3Dt3i75PgoV7IcHZm
F9UgRXj9Rs1Wd12Txx4mTewe9z/qXXCsoCAOR7NxexMI75/QRxmDQQ/T6aO8Qj4RhL6uGlVIJ/eN
CoVrm7Zm/+lx2nTIHluIbh/c0kaoQM18yzwBvNL7qcK1KAkN8l8WiDU9TnxzusKKGeLtnqoxmtUC
xtIVFXovNMwDlNPkMAWxWYesOpPx6D06LOQVrGRk+MrDk68tE9Q2Ms3qiZgCpKKL8ARPT58ZBRwT
4sFOwaEcebsDtI9ML0yIBPDmzFCOqwSMo25oT2seuBRiD6f5mS91utMgaemuSK44OdopFvjEQYYF
cx1TT/tdjRw4BI8QPOu/kpWDSv/K6imU6KbjbcAm6VG4AH97DMBw6hIYy6FKe6rBNTN0BrWMoMa7
2iwZVqiKn73xGAtcCE3GJ39FPeaHvRRIuWmy8+O62HNF0NywxNnTYJRylltjPFSktvj9vgibO/6Q
OLOHJqbqAnSWbiS2qE3d8Q+kFgA6FB31ZA8eDkjuT8sPckBfnHUY+cdHPrtf0wmwWU0Hi7ob3fgN
hdIEtogtJTPbhmOb4WlB2iK1QtGI3041ds0J/DHBQ7VdLkZB0+xQnj/ujCSGZY3ckWkVpEJJiORt
baFYS54YaOZ2BXzQnbZ7XmU4Pc0lyuZhBRmDjJjGGcp00SJubGUI855uK04v9DTsR40nEfFuWD/j
qdQ/edJFt7aYYARkauBoXX+hYmrUgILdpz1ypWGgjHqOId8He5M4vlOoDBTPQcRNs8Hhm5jAnffE
tpedGvUpUhMACeYEwv9rgkmjy0YTeXO0pi87PvMwNwKJ/jKVZOxsMbwnsuYul/zKASRqElD8bf/y
lHkEIeBAKXnNzO3tnv4fGRCTHoJ97ZhRxWdartFmxPcErOk8e6SHpRnKFkWHZGjiq4k5O6BFQGiE
yOuJmyC12WXFkdFsBmqJzAMLH4WweP/0qw0LutJHZmPSnpjnbSvZUJdNqsIXi2Nj7KHs7VFkY7or
xEndJjmINEx3rkvgRVPmp5rwwwYM5oh+F0HmoCF9Th6jVWqUw8euPiIBNb3XIA2OipPmtWGVIbN/
hYeloHCv9judG59O7GoYsCtsET2ynz84rUPoC+cununUCMkgAbFFn+ClkwwO7shbgML1Iau7KMTY
hY19w5cnkZspPngI6seARmKiYFDOrp0y1zDdPS9wbgBDhdzBT4Af2cymv1mAM1+G1jmBkL71eL6u
OT2FNJZ0TJUwXPYsErsrRHEjXcm2qPJbtSS2KMCLC+Kt6/OSYBZTNvkVDTNt8CO7eZCQeb9q9qQ0
dEjfiTfsYeTXjfVJc4giN7cH4mWEd5z0AS2pOY+tHUFeknSARBGYU4lDWkPdYRO7G8IUo9xl1PgW
0zjBb7WG4rEyw9K9CvHQeo8GWaVZbsF9Q2VmBLAwwm6IJPd2gSkprj1G6jDgEVj8oPIZv5fcASf1
zTEyX3+CXv+FTO6xk7ZQt1/KlPRWdRtLwTCLmNJ8YNbOoeCKuMsAn8y5jaH8blQ93w7l5B7AS9Ay
rigAbxJ2bzM4B3lcZBIuvDL38XgtyqgMFWciuHrVFzhJ+tHM+WCDRqCpxLzG7+YmpvJnf2PT/6eI
7qzX1GxglpqXw0jcfpN+iz9St4jSny3RmECa3C/3iPd1kknmMzncrOnT+6CiTeviaai/9i794ucw
ReVd/pd3w/mLPvdTSj6nNVCHuEvFG6ri1jctaZ6p4MVo4/YDE2oApySXp9QfxKrRY8QE7ZeHOqbB
dDLKNuo+ynU37Sxk9vTgR+6Zxq+Wu1b2KWfOfno4gcA5iQq068MciuuaTBlSbKZTTu15EA4BOf8a
YUmEVHZrhOG9smAmjFR2zGlB0jAbf96kJMeXn1cTKadJC3dkuHBifD2pPDSj/FrixheV5cM88nfR
B/2I3dnzwlqkPlMUPSKSzFti0Qw1amfFP9hy5iFtzBUx7Tv0K3KrhsdHZ6U9InAbEVNhK2vZFFqw
yFFm16PlI7QPzkpNU/CGSJ/bTtioh+5c/iIA7WLoENUKzmJZ8ubTCPpYUtFan+AJ1eb0yJPWkBFb
veiJUU3b9YP01LofNA7j66YsbX5ykUeWW3xHU0HTeTnRq44FfmNt8Ecs6V/OX1HwAyqM/l/Asidn
0P7fpqKx+57pz7Qi7TFdBNLqODZ/Az+LbaKjb5blvwmpAaxv3cck0COt3HsWBt4xeuSoA/n3oOoN
hOe6A58YRiW/WfiQtnKWVYdaWdD4gJ4ArITikzu+iCFNAwkgJatr7wS+/kqdYKvuVkt2nru5/HXV
qK+vDh0cnGdFATH2Nb/0CgNcl+U4hVx52AU261XjzWlMOHeTJfMboc2tSxY5BECAUrQ77mwTAmjT
dgQPC0sy3o3ONIjoNh15/o+pEGJuTQJCTKoqaXnq1ClnWc0N2eVrItotRbssEbO58KfLOOyVD9xS
NmSxDRixIqRGu74mR6+t2T8LZ3iOkAMJJ2r440q1BgWpmvZBm9BJapOFbdrQOro/0eWZoPf+tmB7
s+dh0aUTvHlAHanRinYUa1dPxm+xjp96+ao9mZ6YGD8hrILEa4TW7soeZJBdlFO24YXf6CYQP6/m
pb8ekxL5vVoWwolxhirs9sA695zwMgeDEem5CZI0mqbwlJeMKtcPKtEB7mDVKQ9hKaixdoTtl32p
DT2iwi3wB7OhP1AiMgsH6kqZfjoeOHvnDaWVBnqBKyc/ZTI6Bu47L6vfiC4OG5/EtA57m2r5HjyG
fBr6p1B7h8rchYsYgA2m7iJE6ptIysk1i0G+/TW5ocIqkLrIYuXEi6gdkMZY+6YFhfUM1eaWoliq
mbhsqbYgbdJfKZZbvCZ6wu1FsIb0kmmo/mY66nsxfBYtarh7m8k2KMBcLJiftBKIgFxyCUIUq+yZ
Ma2GHfB7bePjTjexk/xpszQAJYOkKZ7LTznh1QE6fsFOXf+TrxBm7uaYzIYoQxg4pp0RQfsUk7ZN
P7/+UJIAJv6GIz/HdBbLJ4d2nADBXrQQl46ac1TSkJkTZOPXfv+ASjEPqg3UVQ5xN77F76Gz4H3L
omcYg9Tu0alCpJyoPWBndcOk0i/ugeCHmRambLZ7Ze328z3KiPj3V91Fiq2pAC+JnBmdiuTUXgId
BqkmeoVIfXKR4ywhvr50J1aHMdBJmvdVhvhyy0k844NSdcc0LGhUJveT+jAufnx9tK6hYsmej8Tn
V9KVOzB3K+krURa9jU7a7S0jkyEf57nFeK6d6XPcTkSn0sYaj0hmO/S3G6eG6gss/N4XKHDG2gtv
7cBOC2ck1sILvCw0DRyENg2Mk0pVRixd3MHq+Rk0cgB/XaLJgAEKpQJ8DNmnRnwxIylnfZniJSr/
rF5XZXEa1X/ebwx7BtvT33TIf1HeHTBG4vzNBN/KDdGXGkI8Tf+hWqN1AabfVO5Fite4lmYvJOLA
LyEiE0lh4MWb2T+2lXAjxhAJTVMtoBEDm19mtb8iCjEUAlyOWyr0jFtAkNFy2gIEu3Pee8k5uvj0
TXzRQ9WtdwteTgr1uk/KgdtyDl77F4EiyAx0rK3GUl/tXth/lR5rxWx9W5tN0qGN7bSqRdTaCn0S
GnnRi4hb0XXf1aLqnqru+jCERhc39d/+thXTt9obkiju/sxnrgPR5iycatK3AC71WVNCFgmYPun1
2T9VeEyD66s7watibtkglh5lvjOpRkShCwHMiV7FeK/R2DjUPmPaxhg8cuv7WBrNlXuQu86oAS3c
bgXP5j9gXBnupksZf60x5/8VAvPUQNw90XHr8xFR3louVbW7P6mc2S0YcxaFBA5KZ1Fq3HPVh8wu
ZBJ2c7OtVrJ8/kTlEAD8js+m2NvUiwL/7NB7SR5a/z1wFWGE8c5ILIONOfqA11VK1azO/6KN5cmD
8RumamvwmqQmAZuFA1j1CLzXMks9vBqakVTJ26Do2c7XapcCwFywCBaY0M8acb03Svui0TpJokLe
fClAD/N5Db8aLZfApAtxhzCkm97FkLQLE1LPDOCpJb7Zdy2OwEkGgpBu0Gun/ZzgaFIzDt8oQpuJ
6uBwvCPzMIEW53oNoFZZE3lwVcKxu++JlOzkN9LACC+yIjGeH24EvYP5cfoxhzPPodLsj5SOOwuS
BQdTiibXiivJADC68OUo0i4HnojJkAlUvVC7N4+KsEfqbHKr+hrMjXl3kCmzSgA/BaHo5mfDlTuC
TDS6+Y3mDwf0UCr6xCb7qqyLKusIxyM1rHcLqnXcLQej8JbrxnDPUdUUmEA2Ea/5fMWNYUjVdSTn
lxrvDzIsfv2Os9pVosBYp/pGmhA8UMYkL1YECWX2LePxRMdJiE6TngM4Fmbphvi624zgjxZr9196
lPMeDdjTyTXvtGdTUMWtVPFnKndT9YGwdOEW8PQICsnuf1uk4mJuQOd3oMTeWcNyH/kQOXkz6yVh
2OAUQ9uBx7nfUUWyDPLf5Z9kGbj/6N4fY1F8Z3eR72PqS7Xmhb+1GI/BgfnSsevJlIkV+lNGVfHs
MiiqBb07SSaOBzSp7NU8OPVt7npfR9lf7DTGvfnKbAUkr3cOGYNJ2gLtXIi7t1ZJr1A+KAxJuR9w
tYJckR421i7TDZT8DxBG0i85lJXqMUosoUkM8T3Sf1n692sCkc/O5WgC9Mrtd0xZSJ4R/u6or9Ch
1wqr9IupbtDT9vEVqlr1sdO/viBxzMiGe756xbKmIs5fzZsHM76722hYJUyOJfH084GsSWHicXvQ
aJk99VnCaFtFmpurEkvmCs9vJCofsVjlvZYhhQTRx5juml0gxZgTNSds8yeKemf0K9kEbRMJ0Ex1
NGt6Fyyc0OoZJyoXEweEUB00K9b1hU7qu/pEXFa2aBKKEGQoNkhT9E45r+xWOZxx6LXGstOW5C9q
D14qRGWJ0z9WO2BkQjDpha8z0IVdUGDCVaDpU/qNJHyhacfmwhVoK/n7VWdnUVZIv810G4ZGlL0y
hxg8cIusJdyEdg8Gn6rUf4xLKjmT/aAsZ2FcAKXx0KVLNy4Z5WZt+6FHKr3OCazhv6Xk18nPTX+Y
Q62vobW2/R/wvhtOrncxRtdYMZ+8PTCgwlAGuDBSByhV9SWtRAghvzN4FU9RX8CaFs+0DnXAd3IT
Ge41ZommIZsouEVtOcg2yKczwl/vjysh5LxnEkWRkfrY/nPGt5oFe3MLzSj32/pIHqlqI/Vn32b0
tdrJlD2LOOlu4B3YyCZZ9F+1IA39kGybHzBlZgLmthAPo5aLL6+08XLnNAsmJ0kvv+g5esiIpSQc
zLmEkTgFYpidJzX3Jo8tFj8EWAQBHEOJtlR3ZfEF5B6lKaP+J8UxNKcCvdoRuTvwjXkNQuVjFHYv
2isDzKHRHFWsBF10WhVxqY0eCFza18JjSdn44j2bxj5T3RWQIWA9Yvud9UKIVzZNsSqUbbp8n6aZ
roP/qRRHcbofcItETJT2uAV1PRLSl97gpD/GOPtCn1rLGLe4lfxaQa6nkm2iTfhdSx7oIPEiDMBL
lCTJ+yurx0C6qfn1YzZoEVjmCSjSKo7VHTzGB4NRUmuEZFst0IgeMn/x3QTil/WVg0wawrfbf/Mt
1CPMVeae1a+dZHOS/ikxXfISLaDdgwT1zMqgGgQ7KeG/H6mrubDDDzfue7RMWjvw6jVhxOetUTHn
jcpRsw9FjnTSoTEk3+8blqzf5apECo88JT/vtNkPe9LLLmYxoTJ5pZRP7GsusW/V+84bATdsplDj
OqucvaQNrRZSbnC9np4hRIQTtFi08j0KVod+TXEO98ks4kNO2fSp97NWhmsVd00Gl5zeqeui7UHf
WxqdEj17wA1xwUD/VBUikCzeRwjWnm1+0pMpCzSPh8ePH59KN6GHFgkM0Fl+Xady24jn8AaAwEnp
a3++z80xHaSD20OUAlgOk3nEovzBM/Rs1UKcQnTnyMkuaa6tbpiDKRAyGOWzC9BkDM/cUHAy/FNN
LncLwp4nqi2GYSudIOt/eCGNm9q6OD0f93VJcqDCxF+P7B+gn0dJML3KkFQ82/rdZRwXlIQuYtrY
s7/kREA4qrzQl8+2KwdejAu0A0/wVqFxTzOIpT6jbtBtTweJIc2rhgdjUNNC606YrH3AGCGybR0s
E6/8RSfsLPXjDYm1LRt34bieiEXWxMiKJ3voL9DF6WCOPQpdKJFWVx0wXtyANNOJhS5fpMDBJoUk
PbwVsZsE3krmmq+TTA81xxX/iYOe3EOAo5BIupN5H98pM19voQNn1RMNWNFWzPMFrENwWTdfQ0cy
JDKDH3oBO3a8kRfbdnii+LKUzBp7SmGAHjEu/Uc+oFAFR53ZtgEwsIVPKs4bVwgMqxNXykSConiE
fyrxGuLLaLs0+ZYQa5HhmODO150noQ7kHwoqJXVHBRNFdMXnh2jwGFv2bQo4XEZ80IYD+weXrEBG
2cxX0ld57iBUMGhgChfjf7xDAZ0XJwfFZcQDoVlJdVwXGdk2yOv+Ip4SRuVRTLa8btjypozAlGAJ
rI/0f0ibHeEwlw26cqqAjiIVsS9BvlW9/Qv48rq9Az9xS67j9FJSbgBLe0UxenPama8OfrhG+BCS
bD7NeTyOGbVhTIP83K1/QOY+77i1B7SZDmr48NHRPVdi3H7uAa/nBJPXNcB8FAbXujqjUMQqHRDV
N/0R3tw4b8tz2NlxQW/kzIdcgae76XlGKzdGNmtV1ipLYs7iJLOWcbXtETFxYk5qcrnv7JaIjPJz
e4uhy+SVhOE+aXwaTQJEFaqG66dznIRHuejvhGw2NJ9rzqldaqHKq8XjombJZocdAO5Daxz7CuYN
s2lo0DF0Goqo+9BMnwTc/oql4CHOqYfr2wCSzcuez/PXMtOzDFpH9TnPA8qldpv/aUK8jgTNpWS0
RgU/fGLOQi8c1qXbslrstqsqWLppXx14gfG7SMyNwjdn+zFObgMul0GT50oPSfuJ5JT45R5Og8Uj
IAzYqCtl8ZuI4Er8v4kjNoxMFVr0/61arHR5HAKaZZVAXPD3jFt8BBTIz/Gb3YolVilmIwImXr2W
5qIHqdpOaSSDqKsvOWOlIzis6XYSMmYfsMNvEez2xi+D9wUr22SwmoGwLPswsZ1cempsegAyGLDA
G9F9XDMyrYVMLh8QAafHNTTMAMCxcLO/Vh5ijgrLd6ju6rDqSKOZTnNbF8JDZO+JNuCUw5P5W3Fx
j1b2zj/gS8sIj1xxUI0iXobNcWrKtCfMvrLrH8d1CSpBQc3OsThFDhfW0x8oARKUjBALPpauIaXz
rDEfS3/NzAnE1vtZHxhj5JmBqMi3i7pN3HUfSXj0j2jYmXF6LpVTWPbMZC+iuVY9dmACjs50NbvB
KC+WEqdPmyALx+Eir02MqfyZOHptInNQzhG6Pl/7GBO4pO7BrvmzmCqpomPfF5pez9FKf+Krnl4t
bZTZcvLQl7OkMlopTaHSV0b89ZEVo/DZDQic9CwbyAZ961+tE36P7/nROq1BGldYPaPHrCCkIDwS
D9Rg4QGvGmoOMaK5XsbcUJp5fwnUwgZ8nXT07MzW2bttvEz1vR5/+Oery51qXjODZZvgZJmLAhuu
xGNNGx4NgbPzZpb1tqARx1iUIUIxUa74EQF73VgG9tgGfVaA6fi4mLHzS2BhP3Dn6mAQQ+XH2zzr
5pH2kp33i6anfI3P0Y936PK5PHlWiMH65bntqF6A83skFkFTUNcziV3tSURBjmMKnlZev4/G4bs5
0fHO2Bko4Eq35qdGooUqdTg8AhdoQALpb1bm58+mHMjSgKBB1V/rm6tdvIHLKrxBYctZHzZNwlgy
j22dXGCgzcG0P+KnCfXD/5gk0DxgzMYQ9vpVyQJ4MEORax8kpPwu3hxVqY/9SKE6a/TafO+/q+C7
FJ8sSjvz8FEQ64hD1d3U3kQudMb51Gyy2xO1zNGknTM/FtMrpjAWTQVBITy5fvjPX/qOF7cWxYXi
QwrhoFzSfnPX0ogVz2wgRqtLnwe96M48B7+9rhnJy+rlxpHv73US8pGm570D+rqCxlAAtpQNMLuQ
phDA8N5K3v1dRmbQE14BzdhkFrVqEJmiCXZCGxk/LLSuCBVAqKtDzAtW7O7Rcub9ZG7UBE0q33/Q
OSKvjUZyU9/cUnBqd8OW2BnnZZCFJSpACcliiWxYHu61hcuIXu+0VaDzo/SKuoygSULdnhLS/GAt
WvIz5VBNPk/yi6z4MU+xhlAC4fG6K95wTfJrGEwwrZYyX1r4mlUM181Fgix3YuZkAJcPa6dTIXjm
9HwpChzEmSWGLGNXSyv16N5ToamhTyBUvv8anjDwWzxjHwZ04Ln9XLlDYZzhx00MhBNquddbkrzT
MJDCTecAsaHcbHT06BQj4KM7iCPzNVOH0lRIaKXbMLbD35ehGKfsIoxgz3dSKsQcOUEFBkSoBogY
ak6DMWCdlshDWgeURR8TKlyWzbrgr35vfV5KmG1PhTRJ1ZVMEDiYG+Hva385ZB4d6ExQPp0sGo5D
MIO16IrPmtX2iMxpZF/0sMNmHP0ApphIeTyKX9E0+i2BI8GnsTfLPnMAqwwz6d8cwPQ4GS0u781o
YDMEp75bz037ADl3bDa2StzZlDaWP+aJFyS1dUiehbS9+zxmls/es6iJUGjnxR1P+fA+NEsIJbC3
duZ3ViZJ+xNL2x1edjBVt6RCY+fbW/067Uan6dzvO69ohU/P9kY8pA9j+siAUg4QCSlGF4YKTey0
hFyb9DCqm0QZQv4VzW+qGYPFaJj6NEv4lNQsNyms/6D2gSqEUM6DQiKF/+xKmGekyLzhe/CnD+HC
X72kvf7ScA9ve2TGhZfyXlJ6ropvvaKO3TK5fJ9cR6hLSpb+amhIxVIK7Kdsn39sRJCQmUgfsxeS
76C2wy0hHKSTaT8rpN9HgtE8MDUWHOMId6sDW7hF1erWZt7jRS5BeFExTlt5ZQW3UM52nYxC9NOp
08IUrdATyE/TRRn5Em53M6jadveyw5xOnU76jlqE1tv7qRqzggSwbCMWTFyJYvbtNquoMCmeO8aT
0SBW5FFimp9o/uXsb1DLPqm5RoGFjT4PiowORXus7JfAYgLQgrOW9QoiFaH7teEsJhZYR001kQvV
z8eE83T+TnwgrQXsgA47MQFL2Bb1a5TAtmaE6ERfLlIvPwEjFn2xUaL8RZJMxlK0GbEioTLUKcfE
1Di9/BIt5wt8cEkwef4O/IUlUzckY39qHqyBalL9Nv+H6g/JbHmCXVVePiJFvW+0U1Tqjr9/aWAN
Eg4Q5idFkYnrJkocEAKIWs9zbIJo/AJ+SSURrWXds1AXZuyuDfKj8vTuYwvLj0kupOBM3bP03ELX
8WLuTLKH+rm8r7FU3AxNROeO/diU39Ns4ZDEbYbrzAd33NPwgmJamJAA6kqIBlvb9Mi8mxtLITkn
NfBaa5d3yI6UmcuYbMHjhW3SyNs72LqxYJh6eZRq9RTRcdWTH+0Wtf1vGLjst9JUP42sK2cKm1UQ
D+diLI01BEo8OI0LlczbC7BFuSVF1bcWajCnKxae/hea2OCFyreiVwlxk7pAlsdOa8vONPhLcgR0
2AwU7OtsgoBB3LMG22+qsgcQZ/0Pi+FMCA8zu/m6ZO4Q/g0tBynAyb4rbHNF/trPT3HYny1I0yba
iC7HOmi0UUHbXAKTdkKrDimOwqbR/AB3A6jwjkvwDcEs0ZTjoUzsMJ68i8g0vy+EHZRCPtuxgW9m
W/dbuXPON6GOgmm/NPVTCNoEFhWMZPNbwG4O4zBXGPgBpRiyocwcGs6ISxgLZHdbx5wxqphOIYkS
FJxAhj17/kRgZih5qX0qP6Vy0AVmp+gC5VYeB1XwpDnVKTXkXGU4msI/ftXxGUPGL7DhnjjUeK5e
D5C3hRYBQgSlfbbXFfSTkjyFQxylkqFn+BgAjLr5JGmaC6zQS+e/gNb1DhIwgY2/szfAYZTFs8dP
nPpcUXLis7BRKlWwLp1yUNUrlHmV5ZhoCUxXxPS4r8JlPhs+kQ2ZU8R952mXBxdRhgRBH/9jSoa2
dWxygjrsxd0onK8zzTkAbzivLnmPpGRfqK5Whla8dsPtlVUMG6fwRqm5JSFdBDNbIGSeXSVtd0gj
pt1qUT5vfC5+c+ArcxSSnWPQ2nXgmuA8pOpQlPUJCb1KF+wjiDjDO1pV4kwegomDFfoLUATyoKY7
gP1vE8Kze7MV5yWh+nVuwB+Ftse5iOTfx2XnrMIZFx+OEneeCjXSEH7Hmg326fbzbKYWfM/BeanI
tkAsCRDLRaw32Ib0ov7jQZZq793Xn3gQyys+GVhDRwVX1nVGhc2tMl2i+S2j+o65FkLSn2v1JlAf
JY25qWbGAkpqonxgK2r9eoLlc5lHZtAiEZ5b+UL/15tRH8dLbUT2vbegbs06ZHzEmKTeRzpOmv3s
07tWOXNLOtfoRmjfpG9uLTYs6pyot3gcWL1nVABGTO40yiAZdvQXFHi5uPbJ1NeUXRTnuWI5lMWu
GZnpsCPOKglsa+0acOBlSWzyjt22IbserRZ0Dqgq25UkMrZPJcxIbOkbDFmybEZjd+KGRcVHbSH1
M45s9nISr1OUW3ETIoh263tFIOQk8yOVD4fvw0S7wkrbjdXIcpWOjXSjDiUsfdcwHEoL4ON8qGOU
cVQga0Xkz6bAC1Ve6GK+tp+R1UARjsCUapkSrw8ynTbqTsoJOK9yCR5IltJg4IzH8Wsw9SF+24MI
HysgvJOUeqqsW+tvxni94XndtLOXKipbt+AYL+J5t9HvBH42Ndvv2qIz9KEJGbOrcnTzvPfCAkcy
43q/Cspw7g+yrB+plI65w1H1pRM0iAN5JglScG1NDctW0aFL+d08qMV0USHubpwj/jHGmruBBS3G
cYziN6eIBfHdY2ZGnwJT8d5p8GtLmbT165Z9teRvUaS9nrmWN4bqCU7NEA2W+6PQ59flFOvaXtv0
xaToiPlRxmxn1C1PS3a0+0jmn7glpr2rLwIfv/kL8m0uLaSfOpL8DAYLMBWDwMFep4feH86Yt6wW
PV8eCLjEyrt0gvlMi7+3np9F5UbiOCFsfgiKXDvnaD0Ny+/3tW1XYSlaabKTOXvKxxUEXooNGYTg
6WR9RNSPf/yUv7bB6JKpMpLJFvT1JkclgoLn2nQjdyh7rHLreYjyvqT1ul5rNoTo8V5iHnA6RZKw
TPkWDbtlJc3yIZkM25kG4nnWSvVl5UvS/7yUEXtthohu57gf5V3SXtuziejQTW7z5FbcSXcg89aM
TGLVayOawmJilmGUByH1LojTOsrqcAZY/hSbL+3d0jLm0CHe6AZ30H86yVDZqvrNA0p+AuRtui9C
GIVAJKOoWeZlbxO6qfAwS9hbIHEDkVgT0D6o39hYA9JcI3W2aEZv+aOHbcDcURgCm4YrhT6Pgfuv
PFTGU/jrp755CzJkevdlhgMgeHRqrBfwoRPjXyzGKBpn0TjUAjPIxzqn/UsKOyCk/SQUh/3l50hJ
DZKpcFDp3f+7neaf28hG7AGX2b8uCgc1mqKAS3q/QN7YII6EBGNgFsQ/miGI+C2d13wB6yaE2MQw
a9e4dpHTryglm1V5KZUk4YrtQJA+1FWjshLl3hn4p8q9ewo4PJbHN2nQ7gU+fKet8OcvNwMNrl+k
3eCLJMs/y3BAwl6mRDiWFdnJ/ZxoIY0wyz9xXWDppsuqOfAibvlpRBqGrnGsnM69n7SVFurcOLrf
RkBNbVep7J6FB0MZkzo60xAcAqV0SMFd7921v300f3gHlYLqAxiN0QWmxlk9xLLjfWrYhPid9Bon
nhuZKtRh9Z1+xno+lLppW9VBWWCSijW0I0nGkpQbDOTMPZlYdDx7fH/2gUteejfZF5K4f5bz0l/9
ZaaZ1Wd7wFN2f6ncEKyrkL1hOELNalgRhP+mkMar72XqwGqRuINp7xAdouJERtkpLM24xPzVicsu
DeupT/4jYW5UjtuvTilXTEjm2sMq6pZ4IfsLJFxBi4UR/Ay7zr1vf2BC1rBGc9ysECBgd0/dxxHg
b/iNfyxpa1bA9E35rBIbEk/mBFAx+AlVQFnkUmPdlmkx68O8bpa7iXygOwI222gyhVoTi5l6bpk1
Nnibd0pk6ThOiOD28Xg+Ssgmdk/zBOni24XWxOC0FG7v5Ec2jDCT7PPggWz1O0j1af9dDrWJHQwB
+626cyjY+RN1zEy/AO0GdaZwdm5i1ez5WAunMV1yD7djIGT01LET/y/nTneADEPp95pMoglPeaKI
iGYQXcWoXPkwDehKlMbQt3z22lvq7tXR7WQkSs3PhjWC0hw/fmTrkX/nJ5hrUnna49jqwUO2mHgM
TqE6aAaykL7VK19I4Z+ErL1oTbj/29F7FD9R6LryJqoG8BlVV0VUqfNITxkBpXdqnRafr4W6xkG9
q7NMVddM2aTa/M+R0Rwb9xzMcUcFUpjEP8Dzdy7EVH7+i0rwVrjoIyv2Db/CePi9G2KOPWXF3AK3
8SUTjOnXBT1riRP/dzCUHcXs0bMYkWHRzhPPgLTfmI6qgzIMvNpmsgJknANhDLvCJYfuEnoEJ8cm
US0vJeY0OrRTKwzVDsx+L4La5tfbje5/6PCIRCcQuvZdfZaScXvrAyd9uTHzc0OHYIPpCNL4/BVF
lDCCzfiXFAUCFkO+qiPtExXhDgnV9V4er9DUIURR31lNnRwut/SMQvbo79k8MaiywcU+E0+AH9/z
Q6ryfL8jWze0/BjWkkE98uU1JGYJ5fjRPd8Bu+bpESHRiXwQYZYkLHq3VXNsXEh76ghnH9+5W2sg
FJgU9BY4gjZ8pJk7+N5e4fJ9Thgndf2m3S5b5RmawFnMedQHCIxjnmBKeiG5wUdD01AI1gHYrWqD
KqN/CnvzyIANrqdOF6c7M8Aq3UEBgRyMKBkx/qzG2nsIPARcCXIj222/lG/AeL1ggQ4PmoDga0Ro
tSQK5OZEMy5N3H/vSEw6dR8dgIjKGH7uau+DIohdueAxlwqvEfQWKUTsVms3hwdImbtgaiMz/2qx
uxqC3nRux94kXg8HnGGk6mSpD/qERekT4fV4gLfEFdvG+g4+MnVNNH4+tUHWXbe/MivpZHlXK9TS
D1+x5VoKkUUZqOjHD1mwIZlPfPESM6RuYHIwPopz7smOvGgxUANvznV59hjmbfm3SD2bI4pkfgWN
bPvazVISWJ+oL7N1/BAGvkN/hDSxNGoUMJnX/gZxL9kSgINgawX9wOyRWSxKpA9z6tjY+qZSbtvS
rSBa3KScCtHZmYe+xBVFy8ZNJnVPRpOgJViDT96YG5T3ZIR7VDTHq2Tk4DhS8EoUycJG9ZzRzy+C
y326dTppoMCRus/3rZDI/nNuGBt57jQ+NqElpiHnUHhaCwq2IMAgxMnA53wNmZ+1tfN5psjVrXhX
uVuGYzaSSl9qM4ZsTXjBtucgqwaDG1/6q4wJDijiS2eIdONkD9urO2rnaHCBc38uHRZ04fSQm80+
SEAAEC2BHpEnz8rMj0kiDwH1yODEZl0c3xMOBzxdSuikL+Cf0rM3INrPyYCanpYrFCI8Covwnzyr
igKtBSkSns/9Dlms3HKFSCPp3cOHBKzG/gRfeQK1Cpo8XF+QIQL31RDQvA3APaNCtE/28mp3Zn+e
CZk1OVNWZyejgzcwYSX589qdSSCwufYwwtd8CyJ8qnTNSqcK37gPyexoP8BLx/FDFdf01x+htaXi
chG1EtzjJc+gSYotyk/7sHAqJjku7ozHU/GnMbtptbmu3JYTfAWjqNaqC4QtP2I0ADZWWF7a91vA
UUJhL1JNCrlZrTftWi1Ucn6HuiyY5EdZh+Nt4gG85bFjo8RLeASGbfsRkdvzNNCgU+PWEesfTJFu
W2BCx4DeRIzMjYkyVy8JkYTkeEBwebUiE5oJKMeuhsFkDt4KPYnqTE8sDkIJriauPlVFMbx1mL+A
xtWxWvwNfbDB5pBYsYjjI2qGT4rNxZMp/AkP+uxUxhpmMvpTGiFl9gbFWaBfpX0eDUyBbEzzCIci
waV/4wL9PWh4WhTKhyYnIgtibWExpg0NKLb6d5ac3QN2L/PWBRAaBsc1sJgScfi7yEa0XheSOBfL
WchkNSYf0spE4ap3ZaKzdO0mlwUotF6wz0dJt8QDpfO+U5EHUksYfp2XVJGAIXrrUmdLmQPp6WKw
Rlb5CNJCBSxCL9HHI7+aFakt71wvO6ojC3v3KZy4XDohfV9F2sr8Uum04BaPKTr4XMmRGGDCdU2H
4Y+Ojeg4Lt8GQ5jNrIZHDYnuvroJnHuYuA8duhrv+zqFP11Rn4nNiH1FmyXx8xsHYDdlPFc7gh/8
0w34XaSFF/aWNCeiu+2irDA1x3EMcOg8omrDoWHmTJ4HERvidGlG3s0DQgs3+ahL0o49y9KR+8TJ
2gEqFNwvUK4smhTqg6VzuT1hej+LZ4wrr0iClLOZ1jYVJR42rGtO17SZrvCR7RLbOxpXmJcLUihH
BJBlHrlF3jmwWpxpYQHX3IaruWkLBuyAB0t97snuJLgefbesudmcmm3KosZWfK1OPx2VGghrsI+2
mOpaOQAcoLkYDJ2FOoNpgpZoFLXxrXB7QtMSk/+ZQAzci1BNjddtb0bZKhf/j5YiBF5LzMyk8riU
y2MvggjLN59pFO6QfTKix50Z+Wp5XW9Fh8f0AgRScSXzomaUpzPsxpH+p14MA8u1RjQWuUUzzMmd
IfNkypeleBZCC1exvfthEmohucoZNmATibPTnjKQfX7FawJiSuFANY5sHpaJomuueojqtuLRYz6l
teVJio+mQSf9YW3mkrtMurqZgVR+jDBmgDyu0qXnN9mTshDe6AxGJejK63I0LosprWTDlka0S51x
CcUB7YY5BvDrK5Db5Zj0Mco1e9ii2UWTPxHA35ElnKJZhyyD/1v/XRt3GoRxbG03eY1OJMvIxBI0
gAz675YZby1EZallKI9XB+USzGhjbyE8NQsulkwqzFZ/h/CnSPg3mTeo9aoEdNfuI8mvD0oke0FZ
PXnI7JGeD4iJ5ohHxtB0LUFZ7nKJNf0J6IGgLqbHfykeddFdB3BhULkRIUmWjL+0k456GxBrZDuI
hs1g17Zk9SRU1VjO6gp5wtZRlyNJKl9yRpBXSO2HSn1NmBiQJsTRSRbxA9Q+Tkjbzjj6sJCNYaRU
W1c/5CowUpBKZBI5JoHJA3ZBPgY04Ss41Gtcebv+g6aS7492d7KiE0S6NFE4BAvkdE58dq5l5PiV
gIdGYjrw5+XzwwQ8Mu1F6b6zNRQe/XA/nCBkGQWNeLrtJ3zBkfjBRT1u+tlD2DsMtxAPTWAY+WZK
bNA6ZjNM5Rl4bsHs+harrAzkeP+E0C0+vP83NgwLZYIr1D8UEEwmyQOwkOo1sDsDzpIpJ70aKQA4
5ilvVcNqLuh5/9RT7FphRaMYcSDw+zqqCGhTOW3YzMgc/BjtqZ2yrcDQh3HQQnCqSoYRfMAlr4aI
aa5Pnfdrh/h8eQ3nBoi88MhN7B7pT5zJbIu5Da7OeJ2jxVX/MNQB+0qop8XBt11EKW/3xuOVV56d
D4Gjf+zWE4hEnAe/066QEU2jY51qH9B5W3f6u+aw9L6sNggMMML5TjCiRAJI1XNf/o3upPpkqcmv
56yb52m7oooDOuI9L1XQ2DJ9mvYC23h0cltxGrPNUqi9BQ8ezrWLznl6F/r5nFgRVj70SgcOO+32
kOLyBJXbJncuYSRbD8Ql2IrYXRrAFHopt3u3KXqDs086UO76jsH8mDi/zRueJVE+fiaFreXgjLB9
f4oq9vksVawcQthMwjTdjfI+xUp07u7scT9DyxH3nTbxSgAExd2CUxmBYPC7sOJRD7dLN6wewTbP
XDanndVhu8sBNbdXj+hFAqcWaZgbsaTtHgr4BoI618mzwBrUaOX5aq2V6tGqOOV3S/gakOH8kc68
L1bgxUJmwMFHeiZJW76KmLjJ/cYtjNcRYiNP6+ZncyD851fPf+huwayX6cq8fYEOYFiE/N0jJJtc
wrRKi075sxyCP/FBLaaZ692jlMzoPbBK+NswlB1+izKHOMhpTp+6Vm+ck1tkJcxGOyTBLhCVIJyG
8kcveIc8fWNGnPOKfyIqiplbPC/jjVm4WBOAcclbTmQvdWUps2K+9aShESZ4Ztq4Hi/YC70wWSs4
4C1vy0xLfk6jME/LuL7NEczxKONTVZlukxZTjFYOz63+CkWEX6s/ArHC0/lY6lfS9kXFGWpGcRux
+cnBAQJfTzdeemsfPVDzofheASgCF+MXcjuVITl6oXlVA9VAdIm+2WXGzctVZzMBTno9uQrODBB9
jFLW4XlEj1Yen0bf1UPHXtfHY1hSZu0Mx7/si9kx0EaPkRspctLxKbh2d2KEbobQn+Tulg433cpY
6xWM1AvVNe9nRS02hFNI2QEy9XADrqMXZnhAj1qoMKLX4HZiGlRH5c2J2CpI1FJmH28m3Wnd+PrT
bLPOTH3s6+XhZynK3+aXluuUhKUpjQ3fQcAq4cDLfR4VvlcUcf22pKuZYizd6LjFb43V+upO/TWp
85TfzBQ4UnAjuCch3gvmnALvsSrblp4Vqafrg8ZWar5hGJWTYKTV5ufRXl15W9mEz00111qmfWkl
t+htncWMDLFleuJPaUggd/q8a59+fro8ZKW+vJrrhX362E6uX//RcVbm/GuYPghhQ7UEF3vkyZIH
zXkufB4pkJ0H1i5qSVUfbuIb6Q3aOTI9/yL3t0QHiU6edTF3NW24fFYc2DMuwTfteYHAD1oFm7CB
AttJn3hT/ngWSTsKIQuIByhOQ/8YUgt2blkfbV1CLnwk7mX1fmHyqAJBUmjO4R1GXR0S2hYjN7Mv
xyuNAsB/qn5SNPDVKu9YaYQfaZCm5C7peANO7BQkPe2JXTqz0/GZszYz0/dveDO6wyhz5XNRh35/
ozn3lXKE8y8AZ3zO0xN3HM8QvozUlRwz95PvtijJwjxLUxl1Q7+5xcYHFgNeVI86hHBaxsxurAny
F/+5yT5+9W5nVA8H8Rw5SbVZ4XuL2SKdM17YFREZ6aMR8Ch2KturvNAmQ0jxADUjFzjOv+xOsvUy
gMRlU7C/YbUY+mhfH+LiMswAHw+gYZx4jbOjUH6avd1aezLcGGemOfzoynwX1dsigI0ihbvjaDgk
sXeUOERb7zhZY0PDV7wBk+HPdzpKdzvdpB9b58hXKYzs5pyyEzlU1GHRwExNG1dDvkcpE+hBaiLC
5ZSLdUnAAkWshCE6xhKKI6elDhDcXunKpi5Ai0KfP7lzR3vw1QkAQWFf9OpSZOyYgMfH3OvvZc94
LaOmTzGi/sH39v2+4pRwnW2NAaALG8enfS42YfP2ienEGg1aNAAk1b4vWczk4hPRtoaAeN6PpYx+
xvOyzVZioKHl2lF7QOaZiCExQHE3B7eRJkK2k7bmwpSrjZ15FuVdPClWyAnZGdOc7rb9e3POT35C
vUIhTIziIGF2rLlia88IE7xjajVGZnHBLO2U1MNr4EZf9/k3sGir7uZFT1CNnYZQw2UGYpCDg/uH
z5OjD6MP+LdLK9KvQODX07B1Otd0boggVY5wYui6qRBHg36XnoqfRrmEy6n5nfvhUzYr5Oi7RYDW
eRxs1ldZWBkSQgvzAMaOREPGH97HtgAAIWYm6w9Hj6PXmX7WIhkTi2jr3C4EhKPwmyuMltav+cqZ
sWc4iQtZPLKqJ6oyI0bUMNFpOG3YDJX4oepjRJMbVSHre0NzKo4dWg4jpqtDk5R5R4iuJ/KOg4Vd
rVP4qiE3UlOkHhKb5pz9OTGMhP4GaWwSHaDczzDkCjbowdgWvCXdidRZbEq6DVzmiOsafHSqPU3r
IN5JTglT+Y7baQohkuZB+PJLhP9GqX5+5VTJ2HFC2fKz/9EHL2J+r0lEbSd9Ezl88G9KUdbkn5d9
07UypYiTVZFstCPnwcCWYqletkg/BpMVh9ijZDzwq3cRUXM855f0VGSrB8YyutaBLVX9x7TG96cU
z4yc8z55qCUHqhfmLK17kE7O+JLenFyDxmMSfZ5LhuLyqr4eSs5ObfKJVfPW6BeufBkbVj+qGXvB
zW3EjaXFL/G8+G8jOzKNZPuCbniipnFSodzCcwbfjQFdZ/wswg7QylAvHMICWu6UMMXKcy6HxvEk
BbhCdFndx0oc4UdY+eboxESJ2kSJO49NWO6jembm6cItKAkrrE8AXC2HyzkvEqugLxiKmShJeTFF
qa0T4psdoG7DgHGqitGIBvlfcXwzkDbrl4SBBmV+1fiBABq773WexGfE8iMUbLCd9lD8MBgUp3dg
zlupHRJV3MwxEGn+YjWIWlj+pBndFXALaYdTtD2iJton0/0VL1/z7IhDT/h23fsjFDG1yukuSfAm
riqVR+yWLmnTkOG8IuvG32CGRa/8/j4iT9o12uSrd7/x1SkaFsZYU9e7tL3n4zOCbWqHgveTvCOn
Z+Gi2Oz5z6t4ybJA2pU4X8lSHMgswtTpjHmAZasukvcSHqSPWck52rqFhO14VuSZEaAf5uhhUKk8
ygC9xqjBXyLa/FWpHlrF/8yWT7mtC0xMhecBFFBU6JJmJVN54MI+7w3nM8tW8F9YwYw8AKcCZEx0
tRstyvwqHnzJJddGWyMxxnbe67s+b7txlDQWV7AstkqAXfFsiENBVDQx6vmjR3otx3MF85qouAlu
Y7x91tZ0KMDECp/V7yMXDPodxejMTFLqMWkpx4Yhnb7/9CABHlLBMgEOdDAinBPuGeXicdC+wEdy
Zlc4jVUYHkTOCESRjK+6s0QdonclF/iIF7WeBcoeXa2+EbEMftBDIeOpne/FmzHFQuGSfc/xt6rZ
G7U55myasYJRqCPJDHcx1mFYUmkiHxy1lupvQM6NEp4e+0OsK2ks3JZ4V66ClvFwW6/pw4fjeEhi
QYRJgLTH1HEbNXcVA70ZT14KKXQR/dllRzjbP6wvOnRTKXddVMRd0uiZqgN74gKIyenn0KRs6RoG
yIJy1qD3xTvanyMFYyWcAluvj5tIWeZpCsKtb5PRKODhK67Jyq4su8hiSRiFF+r015xyH+cTyMtK
vH5C08wukkw9RDLFZa9arMJt7aHZh77puw4VB6kEC1H9mHvkX4UGjT8rDh6fMmRt5i7m3Yn7ihXI
kkUq7SxRcZRpI/5tQgI/K8MymmxmY7uMAzRyom5Mu6yBH7Skix5VGJefaMTpcNOSNxmxUqDkfBnx
QbmeJKq0gQxgxlAYzQ6EUqJRMnixHU3Plsa/R6meF8ftPnyzP+AYedgvk/W3NNFElGIr6idQhkz1
SwcwuKnCk0PutRMUHJ0jGYYJ1yoCTNUjE0oiqS9E3iLJtvZJ3Fz0C0UlTdb0T2TISeRYZcg+fD/H
sKU/2FEFoMYlrDtGTU2S/EXdL4rOsthRjtl4GuaD7voHLXeGPcDFrHXN+k97qnOyFjyNWCnspZbb
VApBJR24R2Y/nd7V2VisochEdVAuavMigIVq7AZBNwPeAAbV6v5XxEJTglI4V2+9qksG3H37NqyT
+WPVR6XL9xsjDVbIA5vWE+bPWLyiv2aXKwf7imq9Fs4CvmTX6GSkeIq1bJ8OlEX6ZvQq2Z7NRyUf
NrM4I9KJL6XamFTJGQeNWorp0Ia88MxOTC7KSGS7amEdDAB/kBOyiRWAZFBKssorjIDaOYuK/MpV
DmlxbFpkDG2PCcf/ovFuql5sBP0x2AulZUtenoWFqw+1RYlfwUnKvuF1OjRmBtrjAZx2LlEyil6J
/6+0BLLuemD69zdULPjMi+a4sCKxtV9eYOjSEBzxY7v4qaysdoC6KW1XwjR6duknn0EW0g/C1jRQ
Ldl7l2/bo6ZEHUyFeFQe2029OOZ+P5uzttNSiMAPq2TEQ1HBt6wMIM3JdUHqNgzwxlzaIKylH7Mm
hnuhJ+0o5rgojfu5bX4h9CSC1wJTpHt/YzxqSFmbGmsYgGpf3c/Wj14topBBa5NX1JBxJ3VoVJXV
NN5/PWFyKCmyRqpqOOJkINj77gA5CkU8g7VVpR1UUVxjkkZA5P8h87+AxERNPjLrq71S1lRRxdEo
KKrQiJptGvxVKeno/rnZoeyYFdD9n3W/eLX0blxiQnYNmjwsG9k/YeYBu7XI28iVP5vO9Ha2l8m9
Yze6VWRJLqt20Dvm5cyBr2El9RnirXrw19c+cvzvDk14AiN0O3cOGIU8FAjpOiHOuOeDAH2E9mID
oVjbWtX26b9BMlW8/9hAcdE38oiYlGLYNUW07nS8FGj5Xxu0/QzRJ9lataEf+pLbFpjaHhpknBIM
tsWbSUQIrxC/Iz20HFYoGP+aSwM2NT3BblW94KJkauNCMu6o8httdMLVyPWVw5vmEoV/WqCnDGzu
pRlRi2aBms1AHSP3YmzhpCuklWdHp+kMNDBFtc4PiXHrGrbdRPQD81/wiuB7ZMcT2FsInFn13HCF
WUh/xZO+NzkLGjY2b1z/0VGuiPjBDBzVlRZgmduMy2puEoONIux8R6200YxW9FoXQX00be/2AKSQ
Irw+djgiy2yOOW7rD/NrXLoeUPoQR7kv+mSVH4dzoF3WuBBcYpyuZdlZEnn0Jeg6jhJoVcOe2jwb
tFVk94nb0fw4jxcFIAsDFdgl44cFtSeNU2RuQrdXZMBKHMqhYqM9NjVK3gd0kNyYkHK28j/qTL5k
sZiORwPJbxIYEduEl1kCoRTILbqkMCYJLEHBGHHf6pF55KJxYiWRpZebz1sBLzUm9InJm6AxWme5
7+g0SxnX53ZJCB/xZ0Q4dxPLRhghKad8czJUnG5DB55w7j5zCzAOtTAq5Lad/eT3qyZFr+5CEaLI
n75bKrWopgBPsQwfGdGvbXUwAL2tkWrluDhyw29n0pOsrkLl6DH0cXebpBJQVId8dMlYJiy6P4uq
O7MKzx0Y/+zu9APyBmSjmEtGHlKvvqjp2fhsvHT8bfqVMxLwWDkBMVGFnmxcalGJwtvg290pfOXN
Hp6/hCUi2lZIxUhs174/kp4tIZDNoXL+iB2DVdeLabmSmdyjdqQhLhg+UzzIlPRl9iTXSI9Q/VVK
WTxpQVMrgWD591dZW7mdMfmdUGkia2iDHvclEmZIQm9EdBTulvTyNyTfFi9s1kdmalzVyByxagew
EmQRAlBZ7KzAnCO3cIfU70OEK/JbthlNe3lZF6KYvP7fNamZ6b6wQfN7UpLj3pPrJspylIEcW+W/
MwlqOxyhReUgJLl6r6on7+mSpyBUDujYr5uml6GCIqKran6giEyAnvv/Nd7ZEKsbNYXnBMTkAF+v
1ty/XIiExh93Mvo7dmYldNV9uqXYn/9tGkzNnnXXUlVjn9v9oS/RHv8RkcWAtMzY1l/u71yffO/7
yjlVcQYuuwPBd3/S3VlgHpELGTU2i5bBYghVIVQ3PxgYQ6pepq9/jL/05NZWCof7Rho6aaxHKgX9
EbYdkrVMK0k3nuOWj8P+BOTetw1XMPxWg7ePNNDKxfflVhdrmvv4JmmGQfWpaM1QyTGaPxg74/j8
bR+z02/spNJgpqaL8D/aN5t4FwPqf1TmcT3/HOr8MgB/UY72hUE2eylecAFFoXn/iGVvJ/4Ae9me
SHLM+MjL57JAQiWhRT5o2x/2Oxq0iiljCjH5x6Jg8jzMWPHQQUjmlYg8pbnwvagDTn6eHhQ+DvAh
dSJxJ+IpjvEdjwZXASl3S3w+g4TJMYo2imfr2iK8LFoP9OJClkyHArB/GrijwzfJ8SpUOLVz8dqX
/mAvMMuXN7Nu8JV5vKlimSO0tADJfIpt0KZzazlGx7CTw64g/kRYRTvU209DZ4NOy/4K6CXrUd/e
GDhJahGkFmtKzo1aAOyqdMZKabhA2mEs19BmrYPtNy3mtUeVkxPeMUBBeAg9utDs+7tJ8ngtGU5U
lT5S571i9OiVaVp7a/e00QFAdEzM+/LMLBPhhlkbJzpr9NerY3GglzXhjn8wTvAJXzo5Ft2ySIBL
lUBfGVEZ12m3xuzt3030iknDyTUzUzKuOoQEglEBInEMcnspVJRmKmmxZ91n0Cl1jq+2nV4W6Qcc
MZP8EMqKMV3KZlww2neJiPftPepvl9iSFts8plw7cvlizMAaZ3fIbAkIsGK6tNlGNqo44DDRMGJ9
WBDxwxEC+DOfhlWvY08pZ018AAo/OVci6evagkH371tLuqOnpLge/xq/8TqRP93Ls/v22ppe/WZ0
9TAnrNEgSCkDMMJ3AA8emjLvTxShK8aeQHIGwf/fEwaKbxEwdG2DwYsuVBAT4wXFHYiaXVi7rVtd
o2lI6HyEMbPvkaFKi7zbzRVcdf2KpMjm0zViOzEg5jrlb77BrDQyH5b2sSd/VW6a7RPs2eY5MlUG
Pt0Olw8e1tCCqQ3TcGzJCqNAwtHxdzm7hg4pKJAZ58HYHp/xA3EV2krFHbhiAMkpoieZ7ksfTmWt
xF5mnyfRk5QRu+lVwq8/FQAi3rRj3VSJqA55os/JDXPkZKwRulUgYy9J2IC31k1b9256E+aCtWXV
ogQ6ZWSMW3tg1gnTtv1G9r9Jjlwpeg2ywgZn1EmtMV8WpJhCEqU+HzKZy6q7ZRY1FLoAkOWQARMc
8PlnYra+iMgw0qUiYMxkN1iRG57y0b5OiAGT+HRHrY4UcW0XtzpB1W2R8lkgUZJwADCEUx1QscsK
bx9X2Zdk/YTTXgz/A12dKInQwMQiStaMj0WtJ+xgWRGh79mDIzxX7LP06rVnBNM7wFm+mL5qBUTh
IqBjZQmI1EpQsQg9Telg6nXK3hf3iKDC50H13eUrSNEm2TkxcLLkyWXblG3FstzB0+o3b1Elew9n
/oWsLjbQHp2oSYwMqF3fXNPtXWh97cHDuUiahoZRg/+J9KjYPHAORSnnhUX1oEBf8TXIr5JW6vHQ
jxXLu1DNbeufI7BC2bhf2H7g+YOJHbqahLfwQzmeReW1uAvacwEIo3Wow0sc7jgCyQX45vA1pIHF
FIsohF/bP4pHWkitw7PzRzhhplzs6IR2s1uXWJIiUcRJY3pclTWQ+Bu3s1k7uKh8a7nJ16kJD7Av
pB9Hz40CanZR3d6XlNfH26BcIf7NJCG2SI+yTNRxyLxV8manv/hz39NY3aYzolQZzKpCr2FbLoEY
yhrWWYvDI5Q10/SEWJNrlLneDM1h3UCwpzi+B/cOGOxM2YfToZ0Hg5LYz0IDBVdnTPFvtD86Nf/l
vpb+GojkenbWykh4fArLTcmFCGfb2ptULtzH+5luNpJgvcqpitcDPHh3KSTt78vqTaVqdRCXNWCc
3Qtm7mZvyowfiymQCVyXVNUc+q5GaKvbxNvAlIy4sGypR+/Xhz2ax03f4zOeUdGl0SSmkq+TCLQa
dm/L4oKEOMg5+xQPxoT1dHmTuNkq3AXHMD92R3A9xb5HFJZ6Y9k+yc2xpxwY1paPPLqEUJ0Ozg+k
kYYMLy0rWAV/e7gij8JNF0XDuagudZoCORcm4t61DJM4zM5+4YzM0CYW5eVOkCn8WY0rz/UUe+AW
ZETPK7U1AHa8/vJObjppeVd8Lyr0xYEB/U/nvRjwvRRsW9tSuheyvpzLxuahSGY2IXuYEe6lnhQX
ZnO2SaLnA/mUT9h5faSh4NOL+K3DLZL18i74ULDgYFwXgV7qdQOlA/Hfg0A69QgXgsWs3uR7uJle
XH0yu5rM5XDYN7sEORjBUzFmuuiPzUOiRYujyxNlTZCeZzjhI8y+OIicVvydQiWY9oOBOZnyHsl/
oc567+Y4DXFUDQ2zcnyfj0l1XUK43d2BLOotui+gWWc7A+Gqv029Ec0CcwtxdYA+lOwEm9nWJU9n
agcC+vTrFT5j/hfOZ/ItFJRAGbI7A/jKhpoFJl8hIpZb1jcLz93FQ97kihKdJQtGKkJZ6Y8e+YSx
zULe2Pdiqs6vJJbJZo/CbwE57+PhX+mS+XI+oQ9U+nz7W+8HUxGGsB1w7PmaR+e5JaOuL4cSsoEb
h4gtzsH+y02a+rCCOkJbWIrYqWANAfdkQAT7y9iBG2Ah8wl2Vynlrj6fPh4fXOz5NdnJVUGNrNPJ
zQv4JSRkNiS/oFLxkZylhm6Fb7yegvXJmKeCWettt88TO+vwfE7TxSsv26ekl83ZtET2EMcPnZp/
SuOV52YXJ73sW8tzLxtmnqXOFU0O5CrK8rLLcWPfLKHQkEusD++P7f4jwfOs4h7Ewxyp18lzjKpw
INyDTOy6TTeXbyou3cHbYSIkS9c2sIwix7j96LnBahu80p7zGupXl4DP4KIzIZBBY6c3IUg3OvRS
c2nagK//Y8Sl1vX4nXRFytpVZtCXEsFajUCQ9yNH5jZ4hwVgDLn13zrFaIMRboaZUoiNWInP1g+w
p4vtxeTJ4/uFtpYruzucnlNjnzr1/unr0kb4YQmRtxvB5qoPk+Bgteqy65UPWAg5OHDPNmaDEIV6
sP0T34EJTXgg4VPF34BNkaR0O/8Tc+dQqMc/P2JRohVSKy4migfGpSLbUK4n8yHPcy2YKRil8fOW
NDgyWVaQ07GiW3CZBBpTGpOkWHJBoVukJXLwBCk3xEZJ+HHzkuyvgU8FDsLt5JQr8Z+mJJddxQ+W
R8GQS57XSNPALKbEH3sC+34AEBtEg2hfOx/tGEzLwylCMQmzHJ3FqUC6xiq0HHqcTQmjeDaj0tEu
wfXRQ7FmfgZQINyMTrE4KNoY2oLbz7XZNr9eehM3rcW9/SPuK+gfnjCWn14s4pELKsETyZurmZWy
HuojgHe3E7yb1rcy+wr4K1HrTCfaUhfNYhvs/MUBs+8bjt21xp8S6F/phVn4fRjt3Nx/nexy++Km
7lkDKpoA9Bv9GWXXwt7/IiE7AzILMZJZYc6UShPMTkywEbdg6QQ7X5YBFOHcNeok8CzzNcIekTNS
7KGVXBosrUhqNJ6uZhudajBg3EEqjrtPuG50gTF6cSjJc5RLVbosxYqKMR72i4+acMSTco8eSzfZ
kkSTfSJTXTVa/ioFhp3cPxvTNauVLOto+/xhEP88H6fXgbeLpu19jB7+QI+KvkMz65B+BzD+IdLr
LgmQ1kDpa6xo3S7q0Y/6Sdxeq6pUcMd2QOO1f3bQmO5bvS5BwRAt4qOF8oE9sOxL9BQKgcsXggO/
WaOLc38G8OFKiyC+6vFYqxl2UFnK6Y8GhBx0pVGToxzwCBq3BixTrQEAcAUI/tSYJJUQm4YmPOXo
pRhiqIqm+MuTDS1mG59JCPhppflHK/UWRAEOtJkgCBWlxyShL01G1URMPS2yc/EiuP31nHDRQoW7
E/LvADMRASfzkcfNhf0oHEt2qaTtOhc63sxetQm9QxkaRGafvXlsMPxUQKt79RCy679PHjxs9hZd
P+a7LtNiypYYragfDt13ztDYOQXVPR3NzhfX7fUXYAZaIX8OC+9nC4e2iO/sCTXzQt9MgAwv+SRt
nKtategHw30fV+sdYXFVRTWQNPALYv2gh5D9eiPSHeuV24g7sun4lVqZbh5YT6wmZ5in6Fzz8N+0
9QAqD6z1g6WEQEtsX2hH/ladnyq/0w7/EV3A+kARD/xpv9oIZAWE7VMltdMAAj8yhPtFZ28HqZPh
g4suUEWkn8vjrA0RBHSpx8YGH52Lx5/VVrUC2JBr+KhvmKwGTogiVl6OQphOpxOXNcFWwrydRTfE
5Kh0wMi4tDAQ1XdXNKq03hY9EI06kRiBvxQrnfObd7skQm0aBDik2cXve7YgFdL+NhOZoxiS5c8a
6TLfzmovpm/pqHRnXaNeFmw4BtYEdNfpgOT8w41cFZtqZuUKpMAa6RBtHWxKfR5gtFcNP4mkjQYE
y9UXS0n4+WyIWBtO5GK2NOl8R8ZfRMjRELYdGKR4UIgQ1e+aMiGcLzRxAt8U47gnHqjAYsVjenn0
DEARukuk3pylt2b6ANB/yrPdrlnGQFB389t4CSWpRhrjiuw/y1vcG7GgU8ON0hfYwDnRDMi7PqbN
zQ0WyIYbes7mp14kHe/UXlNCcQa6D/Xi6gK1dziL6jWQ6+cZB5cpdCpuIymWqcPINDZrtTwqM6w4
MRRKVOIoA63hC7qnVaxnYHU4SeaX5qW2h16uoMaCP9DPihBg1S8vl8BjM5DrDlvmAak2cATX7Se2
B6+wYIsAJGQUH4n79i1O3/ySmH9D9J27GD6t6EBmpajGI6kIBAz/nMIJAx00zmilqTYGhnjYKC1i
dFOPZ2Q+jZ67mcVYHphRB+KqiFYeC20zhBuKd1Y52iDAkT7BbrpzI3XDRoQZeFFEYH8dDerESpK5
xx6gMMxkNQTjVNtUmNx/d1t986BTe9w7FNPlKaUAwt2CRLbor533f0N7vxA+BD9USQFQBoUQbzck
xdp6kLHTI77PbyP6gG1Wzl1MaXoIjL6mwyalg79/PzQ0cC9++rTcVP84lGqZsfl+mr5gf8bkGSrr
A7+uq6B0dp9jPQQJd4edEEloOOPwlUa9XVwsZAEFAwyM81N2sSS5XD9riPKlQL393FcGMMknX1m5
+A5Knpa2DI7qyZQuNUkNGWk4phdIJp5hu5NXJ67RaA6w1IotVM27/VtflN4vjZRX1eYBt+Ufmci4
3a0Gwzhy/kddCsiLvisEry82YdB7LFQ6DpmQjTisPKkdqqjofFGGHTv7pcskvSbnkuawiuZzIGe+
TTeb8zBXjhb0/9RIq1lbSdcxMmNmo57i19uYnzIcsCGiiOnS415H3w7rSIgHAC9dbtQJou4XSevC
Qjqo43+oFmxMN1StTWlrZjZi+Lxn3zstlmVXUe0SB19m8d5W1nwE4/97CvqoeC5Z3+CCWgzlu0EU
temsk2bo6C5mXx1fP+ulGVzLIagGBtnJrUWEIVG2ClFP/UzAgkRBDEOgxbn5ETk33P8pkkoTQfee
Av4i/u4DMM+Ftb0GxcOtifJaxJyRtNDpu1f/NgYwyOWv/VUP0ZK17b817+9hy5uZh8sK5y7nXkYH
Xh/bVDFaMaLog3gsN0FTClZO5y/L9Vz3WLItDJY7lLQAc3kqS9y50bXHpC2pQSJAXdzt5beUPwsC
iBXuaDu0Fy3ynROBZ0jtcXh4uvFy8b9iCQbU/1w58Pn4Z7ojCqr+OTYvdcj/6bjMegdT/Z7ET45S
P8zlHs4tYcM1yhi965GU5VRlTnDGI63NiFQjVjTGzTvwxgBB0C5vLQVYkKmRCHNmfwcuZ1REB1Xm
hp+ZrrrddVy4R9rv5/tLLGDqWhCUxIO30rh1G63JxfB1P4wSjBvKpoXeuc8b92MJCVCU6gjVC/l6
sFLEjigs3qzvJU+EmqE2u0cxN2LaaIspQKpwswReueU0j0FZn2kbVJVS+BGdKdczqmlsSbG52URu
ClDetQSGw2I0GV6hStV6qXh6JKtJCBoJhW/qz2rQDA/HvjT+XKKbJEVjxgt+fQ/a9V9/qasgYAS5
lZExPfZPh1lf9fBEGDAywONK0tzZiQ4+cl0fGc6eR6rW3tsOzn0bEkyQF0Ws5gElEbQG7oM1vNpl
Z5sFN92yk06LhwPCLYT7f8Hz+rhTlPpR8Ah4K4B1mvqjB7CWPX83iRZTU45Q1qqpm9efvuoJH1k2
U1VVRJ+GBbNa393UDHlzkkpcCmQZdqhXigiR9wFxAQDodzUzOkd7UxU8OA+3WYn/TqYzVjs1d0W5
+jJJf8dyG0bIwkkpqdfl3c9+qvBtArPFysD63ghP/GuYK1mfpboazwgFFtclEeom/Ssrd+r5MInz
kyr4ARjrMbIKkQpSikQbC1HFo6o5z8SE65cCoDulq75qeqrTlOmO/CZG9FvDptY+nuS07ODlIQg0
Zjti+V0KBMVHrF5Wc2wj0ptpa+8J/xdkC4rL87/SQZTvX22iAl3C7i6R2RHA4Us2ykCVamVnVY5A
wg/vBXy5X7KrQN3cZmeunAZ+ALSx2G7HGlCTqLWj+JRUL+ODlRWdcRzdS25e/NZ+lyeVN6iXoyo6
37hyUY7bOkwvdnmWRbvTdv6SPs4IRTX3k9qkbYymLpdzPnLIEkIRjUG6eZpjdgO+s0oLTIElq4Jl
iFbl4xn5EJgiz0kMitefyn4sKrxyEgJdw4n159VaxhNnR+uQVyBv6WKt79rro6NI3FYa8ZSqbjAS
2ms+O6NiatH347thXuNeMHU5fVxGvjPanEqrYfFiWieL75C/vupVLs59R6BYo+7V7G93Jtn/1Dg+
t0GjWbdu9S6Q35oB3k9zgE0SUJeP/FSHKZAvgMYgk3oEkdnjQVUnfua8RI23EP4LqYJBM5JH2jv9
hchejWs96KgtX49Pj771Kc75twVU4DrpW3HT6ASwFniNHovn5u6Jolc2I05XIbR+3Vci8txDArxv
X7x4L0zfrO5+GvoXdQmpzzKdYAPpsHyh2XIitiZ3Q0aUPwNUa1ksrz9bePn/1FX/SoJz6w3Hmv6i
hzxYspCOE5H1/+SQfB5nukmsxgp01P7rwY/WWlBYkwYHNW7Ym4fFtVKWXEwEPonQD30oc4Q4aXGO
JjxAGDij8osJK+y8SjlhJs15jD8dwXFBPsBjDrIBYBs7gz8sxduT9SDmXaYiT0mQ3LSaX8X5STVX
y4Ggqno8N5c/K+wort9SN4XfnKJG2cuB4/RL0WqPgicGbiP8SH0Vb1KZ6lk3fiLx1wJ85AzcEU6l
icnljFUvBvkiB5eoTtAKrNtlz4Gy7tQ69efcs7ojkOESyuvgR0n1AXtI6cwkWrACJ+RpvB/4OM9l
2ay/r1QbNKnl39ievp3gFiPhCt54kGHCNw0F51nCmbWACCn4fjauv8zZ81P7V5yXRLe5f1/Pnp/z
73cD9yEjbfaH75jRllz1Hr6vSl3TaxpgEyim55TlkthsdAeEy+4S3hPvPJJEN9IUcSJ5ZIUmqvaW
XkMjqW+BRAf8TeisR3EMJxTWcWBO8U4M/Cj0l6YGMNmOY3veVDMFIDTBjHu4SnrvsSY/89v58s9b
2+jom7pHVYrWwIeQXOloA2vUVUB7giaSj+K6uYsuc8v/k5PNmegHs8oQefh7+YzMFyv36AsxLKmb
4m3lHSxVbJ6OQL41MIWf2Dkv+7QhdNEY+Pb5/2DdLF9oc25bmfIgWCUpynf3urMdNdYSEZ2MOCMT
RZjT+t2nHDz6PrMuH9NJ9gBah84CBWjM1Ho92yHjK5IYt5Xm/1hvNUhku63VjowrlfLk8u1yvUZ3
syYOP2Gf94ggylYj8w2qmtHZQIOEkh1o9+0rNHGXtTN1KBKDxKOce/JEm8MBQfbht6u1BE0MmE4I
bkGmISKuW6YsagM0QuG1PmwIxqcaP24cWRVdGkCmTUEyf/XZtpIxCWH99fOwQ+LThIQXaQNGRzxZ
nvVLwQlJnGAzKYow0GegLCq/ewMGTfE4vdQe34g941LDD1e7aoqtK9/GjbJ43T8m6/86NAlxXSMu
nkAdgN/OqyCLth0Mth9iG0uYV+NPe/f5n6lFtAW/lvRVwgVxkp+gINv5Fdcx91WBjFo7CowyxB87
8U3jI7EglEG/5WWWx9sDtVQrX9OSQIcyVDUYyT28YTJRrQgAw/xguGcAb5lPvfzIDeTRAQqi7u7L
MQSjcEnWoWWQGnwPkQlTvwr+xZKWE+GSM0kMZlBkkA++xc0v6BO2DYvz3VzzfrBm+Sz7LpG4Sjvu
Ewc+uKSlNp7rUFNPkml+se7MOIY9sZ1jNBH986n2KuqSBMESfSh4D7/USGBKGPBaHfF7TnTOL4vQ
J5Fc5lBPWkecbYUaBidd+E4j7OInfUDLYbvQld2Fl+uZGCCZVGpeJo/bce95b8OEHHxkVLExZl4S
YzRIFsFMaX2izWf7+9vlFLEB1MRUdrKIiCNSmPzitdPwo8ft+XcL2NC9EGDp70hix34FA56QKaVj
jaLLXPdds68pURPA5t2wQx3LJUAz65Nxcex10Ef9QpiJl5RBkKQpLFxXqsL9pgvRbAlVJwIK02aq
qWclU2FzxsT4AD+/3cdJYWxItkn6ii+GOMxWHx6jnMWBvbhi7TWAN1H5dqb1Xis2vGjKgLOG+H8t
Wsj4S4+DVj7T/v4RE4iFHOBvGxNk+Y9dvHgtQOsaFAeHN4qnw7AqV7a3+FT6FmCr8/q32YICa5N6
uNYycaP98IeB/qf8gRMVWlzGzXcUyXZqI+Taw9ktPAF40Po+kzdnbiqaIorHmllPp5p/j+Nb7rTa
eOirwAGGm10xBQ8mNmBv0zOY/VK+URwNvn1lA4cmYH/uO6RKItciIDSsLtNUemZs7BSftB4y0YfQ
3dWcjIqJxOUu7GqjwzDv3qDo1d4A8ZZOnMoc3Xv+MLsPOBB/yDf4RS6mb2fHUBlS5g1afW6BEpuM
POkKPBlHMfIjzz0sEgoabygY9tJuQ5gQkMr0zLbIxCrt3igJujYBZMyJd/ujpd3XaHHg39KqsT38
/xXmDGVgERF1Hg892JPGr9P1zaplGSfcijKgOYPWIqOux9UGcMEyOw2vsNQYWiPpKJMz7RJyRcid
DrwKiDewOjndA/WifoKbR7Yk+VB4kwUoY3oGpbG4Drdu0R2jKmSrHTkHXNay3IvkfCvu9A02IZ9l
BEY223ES3qE9JrioGQ5SjwQzAHfHMVJk5Y95MsJTo2edsLbTZofEU6wMZ/qyRyqLj9FzoD/rcjmZ
Pq8ZMC4z5Ylt5nfFZe5GUz/AQfL4PXgQkPsZyvvTN8DqDk5C8kw/9TJC/yme3euv7i6MZ4iCaRLJ
Yvq4Dqp1sdxxDWK80aGEJkzAs0TQD2NjVhwnSHKnClY2oO+UIid5/AfH0oqAb6zLUSl6ilz6L2RQ
8q1G2rb2x96/jMXY0Nz+Ii/ejQW8zCYu/qP3kFLC7vUloAFnTetfbni1daj9OHvBJ1F6tc34GBIj
5qbK1pLJiSh/SHoJfcyfTQYrVrdCjgLVQtVPeCqCGfFYH3E7XxOjx36+oNemXdeC3Hok2MXrtJxS
JekdjQuaddpB3856uRm77IIl79k0rT2hbeQ1G07xWkIlBGE6QqgTPO64oUyjdwN2XDipklozLKHC
9oa1z4ersw0009OtrFOopOwSnFDeGAASKacbEsL8RctcJPDbNqUJEeGKMv02opOX2dbCy+F084b7
h8VElagShVbn0EXZO922QiOEWHxz2F5t+3+Q9YBnQ7mW37fnlvUs2GqhhCnKdWr+ps0YVRGY42Eq
4PxSzuDFFXotCYQOQ+6znMY/o5dpknpz0HemR8ND5i3UmwDmx3CZ+bBY4uBbuFHo19+cp9IVfYAe
rUerU7mW6iCHES8ltu2E1cY7whUGkl5+DWl3RU50E0rGbqutidHU9DR6igXCJqWEhvih2MS53tTy
DgKzGTkeNdKyaWCkvkJp3aqel7M+QgMKxAoIs69zl/m6/FKvLAq8utaWPrbHoYFqIZfAArXVa+mP
LM2N0GVho24Gz7b/T4EwiaoLv/4+rtl4njuypll5qUNDoI8f2pMLOjEnDE2I6hfKJyFIn76aA1JL
iF1dJSTBk/P7LUAbYt8HwrsvMgE3v0gBMxNTu2qRHxO3URi1LaWwQrNXny7kNlhrREkfRc/5Dgdp
JZhGekfAM7lbDSE+J/HjW1AyZ/Db1x5sP34nnU242oba1lXs65MH6k5UtDZprd0p+EO2R0Fr2kyS
uWJXhVklrVsk8g0k/Soh2wD32j/bNyJYI6bv1sLy34gyXUJBuOLEXQj9iYZCOBpmp6hDcBtDAL24
2P9708YDNTuooMH3kDruUWYITWig8bIgR+E8dO2Q/gSwEEAR1KaxONLadpmPpgOsFRIOGFFTrMC6
PHMG+Oqd4NwmjPaXZTQCpQoDIBRuMklWeqtZR2jrvkX3UC4PlLn7BPBDBK1XVtr4DEWXud2ztMWx
4dno85PAci+Jvq1udpb8en+CucRkkIKR4iP3Sp6B4TBTIMnzXLkaVHu69LRjZgn5jWrev/vO6pcg
vuW4rdK/x50cJHmO/65C5g547Py1nfk5Uz1Aqs8lDJ2srTCFWcpnLwvwJlOlmilNNzbPyY1d4UrH
GICHnkswuDouGZammbiogXsXLaMX0uEHS9FkRtamhutpnPZoiQRTyM85Jd0AVp5faKwW2VLpJPgS
b9OfFSqQpvR/lzdwuDmCn7Cah1Yub9k2qUgKmnUm3FaryAAQyvPi7QB3SU3IhM8Z4UHdBLodaUGx
b69Ljv8Q8a9GD+HGQJoodIm+s5iA20qVfaTJav6v+WbALLbjWu7qonNv1DAEpkMXu11zXEaYL3JN
GpgjE90khoxjlGIVJot8uH3mAA2N6OJglxOpA8tpBPQfNT4SE3as4/HTIh2DT/w4JWTYQ949K1nl
6BuN0VBFE851AYLfscB+7qNfRTwuetGRzkHi9O+Oln1h59Um/MBevzvdQ3wWB3aVzW9vR5Y+DwGx
qRlUbvWmHEwGWo1szgIgOFWp7Mm71GQ4OkZpzhcT+/tr5o2f32Vruhc3GkliM4jAKtwoNhUdOatF
8h5ni+lF0oGju80occyWNnwc0ae8ooAUzqJdbjFqGE4Orz6Nga8CHqwRuTj6zvvDQYPJxiov9y7D
YLaYb4MP4tiRbkmhkQ5UV9PMJ2boYkUTpIcLrKVleezTz9g+nq3S1GS2lPaAZi+7IKXJs0Bq+cfU
w2bx6jHPc4K0EIQC4b8MrmQJ2SX0Db2ZcHb5sALkEOaViDkMD1w/tSLxboBvf8tzoUkds2qfPGIy
MhUuHAALWodmXtEljOcwD4/3d0VaIsQ4/cvXUO0Ui3iyEWu4XL9rFZd+iNIw5n7CffIf2tYePfBI
QfGVrVbYNPfwgJQNPOSzshyeymxO0EzgYPXL0FhhEFzaYkyKsZd748Lu5AIEsbhn/6WyKZOTMdBH
ZloeVPPOkf9UjwExHuZU4amGWWuNFBg1Dhj5ZOl+ZjxWP90jPG/9kk7+B4PACRwkfoxH556QNJ9+
7xFtuZg65x0+J8+WBI5RBQMxBgRnYDRvbqjvwdMxKIlWQwjhm61WAsuxhC4bF7ATAEBNijXkJW9P
drf+CtURvLyml5aOvXX0blamhq+0/lET/z+BQgPvdtkjQiEp5yLkBjb5+JcgO0GsrsWAsDlrHcOn
IbY5PD/yRqPqXhdmJEUkgDmeRJmxj4Nmli9ic5y6q7ggH4WNHLN0Ed5qHtCUiXhfIICbZN+azmpj
G9xdP+JdxX1kp9ze0EmsjkwXsD0hITQ0FUxbl1erzNl+IJz19Gb45HYl3cKY59gvWMbyWZe3cXlE
eFrVmN1gva25PYa536Ik4xXNhkwBT83wLZY/UCiaGp9vqOTpewPIOIkdshyy/Eyw8o40RAO+mzXQ
BNF4RnJSIQ2XflETOTSbBANFmV/tjWngVxmUYqHnJE8PCOVbsLgxygyvi+sowtcppIzXWjNS5UdQ
zy1ypuXunwyGjjPRzaxZAB37LKBKRoya95aMHk1kcxKDeoZ9wbsV4crVbp6gstQkgXxKzLZlQLwb
qtj+/baW1nXwnol70kQH4o30DRrXG0rI9xAD6TnNruhdmNDPI9bP+v07sajLabH9nJp3sxLn789v
CYEPqIUctFZoYNvAZqssH4xi3SOEhApuwcI4+C4OZw0PD+EKUaGvBxG4I1C2gg5RCeW6eoq9wmto
zyikTclDH8xVUiPTNg2fsFUi3LMauQ43De9GTxQwuUJSScnrsazBKzjlK0VBuczfabHRVS8oPdtF
awd5pHETx4hWSTP/Kg2gm5XwyLG5r7TdzjqmdJSXGN+emoPTIlBjji7otZW5wsmBDkvZvRyePRnW
8b1ssnxiNArAnDYyigqiBBGWCOxLIGovoKEc8IAmli8u3L1vOaHrkfBjpxMdMt3Wrn22kq6CWNVs
LoER8pA0C6BQG2Mez7XBiLH2jNlAeNmt7dixmxKiw9dHSHZoczTTZJ5leHDAn1N8VInmDffIE7aF
AGe5AV8/2v3sNKLnA46ZRRkU9gIY6QhSpu0LzivL7pppbgRC4MkBU+99602oYeewIWRr5V6y8ri1
fPUSbK8K1a5ZfBh/DXJk/r3MRcuErpoMpOMuR0cz2byQtESh4GKq0OUp8IGRoVrfxQhWW5hrJleX
ehuOq9sKFXlPWZbGe4SSeXetRQ9NVTdPvhue/C4J3WKeok8udKwEySrtP/+bT7zmw1RsXCO+FuA+
WpTP6bbXtjjP7PqBq6FJcPjWkOBWh5v9E4giKE5yovsLVBtCL9gx/qiRWDVkmtaKfLg15fWcU3Mi
BNGv9PqVczuQ9ZOFWDHJiOIoJWBXN653Mz2KozhpFTsRAFOCUp1UnbDbXYcSnJcrxH0kga3NS5OB
9X2AGhnu22GgqVMj56aM0UYQ8sLiSzEfARBsUOCC7P90wqCwcW63xSsuXK3iM47IKWYT/OiUiHIB
kdhlVDlUigK2W5rOc1Y7km/imk4InPQ4IIzotMjwt8L8FnZ1HApAwOMdiQegOpdUc9xZGuNkY8/m
oEDFgqrFQMqX0KdKwpS1qyzlGuq1iKKDNzow38YKwrdaVLQlQ2eZXkVh2/TV3IALnxa+09WWlKG2
p8W4GCJm9LLgMcW/WWgJdx5BYc91whGcBsH9FGZmmeHI+v8VlBpeP2mpcaBnMD09UlItSC+idIup
Y8+drqjkg4mBUEcCB8QfDyaUEh0tgl52k/NCaRxaJ+VwDWdryMuK/gIrWhb1mbp0rJvjqag+BKdy
YN4450x5NqWOBw7EHfYbbWACCTSoiwMRWPS3qTiweasyvitQFTGgJRpdYT5h4dMHCKfp3ubrGQ5g
bN4nU58S3Qga4XI3lbNWxPIYQJRU4RcXP8hhh/LrCpXBiSjGee21jol5S2TD4JNKYr1Ip69ITitb
vyPNDDVLLEsu7DLxZqjZPYZULhAwyuUh2HHxFvVNYFvNhn2ad3rosBWn7W1pnYkScq6SNoPN89vS
ami0fB/QgVJ3c3uUMrmyBS10s73QL/PI26/8u15nglt9+xFOI/+94vboC9dCBR46LpL1vAH0u5ZJ
WxVNeA84DQYP2Pcq9mLqxSsAKHidIqsX9vj1+jVSRoyGTEeh+nYdXz/4BvpdxdMb3nAkxdEVE4gS
YxSmW7jOJAKcrmm4cyVSKbB0vh6CVRMZ4TJCfgo20OGqH0a3mIcaBlYxJxd6AOs7qr3EK6Qpjned
e0Rp7dQz9ZVW8bxVNiqk3fi2g6OBzvOct8MwoNfRl2UdOWry/xSX2a1TNQkPxOg1XhEhhkjDXeod
5YyVdcmmYo1eJcF3YfmLO9/GpgZ2wtO1gVxYUPWEZqmI0YcaElhEk1dHA8A7l158uLEzZoQ+x9nY
C5gmI33gc+NS/dRVePKEj3eURiguFpfOTiNKvaj45w8pyma8bASTA4unME+mY9sipUNN3xjWt+KM
Gd8bSoEMoWm8lbFZ0KJPmL1kNDlHhPeFrcarqV9z0P7nMv7C9t6SBwXdiDYDZc9FRN+LZSJhj83q
IurAqzKvkFJNtswZqRZaWJ6HkxptvBtDtya0/uIUSWJTVYfUNNYVhlZ2TGUsCIArysjUF0fCxLca
XNDII4KNcDelEhVNalhF4o1TqZDkjbfAPsuoOwgRjkkSxFDdW0af6S3vo/6ldMej2OKRk7MlsxZT
gCGuDUpWCrYqpL+If6UW1fTvomuXow7aZDgR5iUnk9YZp8z4UUKnZkruHgDp5ehRdiHGnMVoPE9q
TbxlNn4CbOsdeZ0miG/6LGGbaa/L1EXjowEsTbohiAyd+nnuaI1VwSQsfJ7kKuBkavS8S8OaFhsH
jltiefecSvJUYa6uR201qCEPlmBCWiMc7j2om31yjyeVQ3NcyYGYl3WUQQhwTqixmgoRjHFlgDkT
iE+EGplC8XgB9hU6ytdKUs9T/FWX6HWWIYgvhBSqzUX0q3qH4wrhVqlZlxE5XRSDXh+hopR46oHV
0T5/YEna9fbEOVyDRtdXMkCu2Lp7ZeNGnLF3ogCKEKvWCTo3M1ygqDZm+kBwfKdQwBZ6ewwGaQDO
nzdbMJLZtIi683yRGh54a5b8J7T8BumfutOtDY5xV3hQimV7jhASACudsNYp/UHc87QD93n23yWw
eqCjpJgdxweUUO7uiTytyShAGhfrQsROhJDKQAXAR2LsFxVBjQA505Q/p/x2oQv7T0B+huNeTEek
rNWsK0Goz9deUMA5G+MNgnao3scF723bylV/kHP9Y6uXyaQ8Qr9ETVjXbFjHarA5+2JmKNzA9fQp
+H9Jr4nZ5BM4GzhcQd9nRjcrE6kuB+H4XPnmUD5zoVdoONgI8sn/fpuqOUPq1XW+0CyUvmeIDuAf
Lqp5WYwXvc16zJKTYcsY6rUvDhXeyj4WwIofNnFh3goRkUvQa1xdiRvfUik1MUYg++oE9gQBL/CG
QRu0aX0E2qWeypF9wHUpbYoaonGnf8waDOWgZ5eJoaMbino8uYwO2q8O3pIUwIEFJuzgOv9D17aO
0Wgc37h72aBmDHSmaKyBNbwfJE8xKojEqIUXUDxXutbB5U0mJ0hW/tYqCPm9WEKNdB/PPJe3Y/zN
ZMJ1FuHIMK5+QIxd9RMPyPMmNWQ13HjRERuIrZukIgZBlAn7sT3MT8d8dB8NsLCBemc9vaVeuD1T
1UBolkSiT9WUbwEk7jIV3JIWfv+E/9yekTIaZ8x2KEBXYOdQ1Vx1IkL4bm5Vbjpg+/hV9uaiJdkQ
AnEO2gWjwcpf2Yp7bTHAY38oDnVL5rkQwVxBYR2fP34Rcsp/2YmxmtiC3WI4EzYCgXs/aqSnBwUU
vOLeKe6QIoUzdAMfvE12/bS5uoe8qeeQa02v08Ff5ooMVhImu+TKEfiw0UNYZ8af5B1tQeLW5jO7
rwhnVsKh/LAXOYlUWeZ/nX84q4f+Zf1QO5LN/j8l4p8j8HO5SMNprFIC7QQhaoT8/quUGUGwIJKC
cQxrLO7FSV6KdxPTudHnEzHcvpXKdhP1o0uJnyTLnR6t4qXbxLlFTTs3T2DjqgHv6ZH8QldT1K9D
2S74rD5TurNbsw7VmdKscczoP/ABsuJsY6TTzQpgKtGI4B8QJbqFbiq4xo3dkA0XdQDWFNnQhV4t
Lo4iIw8o7sLD9fqydP1D4PQn8KlyMPNFieljmqeayRLWKs4qsmbCTUuoZDriu4zuegABvxFwocsv
WgFV78Qqbm/XMpj5/Fj7JflicMnwKaYOA7KOiDdzlAYr3QJyWHn6Auu85077sFzGacGFDyQuDahv
x/Sfs3t4WC9DLGMqhJhudlnXswib73Y/BeHFCf1+FbRBlsiqPviuCMCeXr2KluPAHYmGsx7OyzLF
6H7BmZfaWTutOK2M9wrKzf8zOQl1/9Lmg1KcBCYM37MMA6cZln7OogWEbnbDaaXbxWivjYWyK62W
imdYavkUht86pBusa4nokrvdhctHeXLa1IuSGkEKFcU8C9wnSuNPOSQMkcV4PPx3pgcWC/F9Cfpt
Rdoe/uqo3yCwLLmYXYzsu3MJ5S0SM9z40e3jTEqrw8IQM3VbyompRT2Vwu9SFwEJC1nzBY8H5t2g
r+o/0IoKWA07LEuNzOZFR6+zV4m7EUlmE7yuNAWOIj9XY9q24fWQhrBlEKMuw0+Eu1s5c+0UUknH
zhWFHmOnsL2PbBUPXQWweS97qxMhCe33ZaFH9comqiEu1yja7ZWweCfvfyqobMnohxNKzOfUHUtu
F4vsQBOdmdLFrsTybm3c+hSbqmSuSvfqArGZYnN91m4lxrBS+ylj2sK0ph9abdYKgb1zBNPCgHsK
RQ/2ZFXq4ZZ6whs1RxZ5Gv+7dUYPggi7C/K0WY9oTYlcAzkRlaoshEKbIySZczpFiR43VRImuVzg
vIhmAflSa101g+ErQn11T/cSTcgu1RLI5ZrPWvUhA/YJHMB6kl/z+aIRqnWFK9D1cKBXqqEaX6Sf
MGchrXvP2k5n+XXmFEbJotnJyw5ykcggQLzhMCjWUF/xt4drMafBOSeFC7Qy0Zaq7oIFsiTXX7DP
5iKGOjBrJG1293Kk/pwUb6RPHJ3CRclCQYfWeHESOaH5MVo3XAx6+8jRMq8aMDoRovv4ABVS1q6z
wqop2CspM9tbZYpkcoX8qDTjdWcHRXr4aFvv49ydpuj5exK8KZq/qncts0ckkDOZC76I4h0lKHru
U/w/jQEjTgEFQAxfhIbnQR7ATjTetMiEOIKW7ku1Q0Pvm199RzKTXuXQfyN3xoua9zrPcz+Fu2Zd
47tmdDd0+J7ZTUFXGzkVN4DENInFYMRk2LL5lWJuJwZn+32eMoP8b3SIcFDQYIFOalVry2jLTmZl
fq/F9jNxe2e2UGgf8LTpAYQxK/b9TkuZ6f6daPlNc7jVe25jM054/pMbGelgFJPvIL28qGdtPqGT
w+XM/c5BgMznMwl39WO/3xfrycWWtHnN07DBnKYpIXY328FlIqW5dYRHUh4osiy3e/MvuK14kSh7
fME/RRcmOmHYm9qER0nAjRD7jYK2QW+5CUfmjoFJdeW2T2lGGGx7SW4gmty60LGBYrsfsJFQCcfv
7J9isoE9eU1mOzo9rWjMwEdNt+TbcZZFwluPTWVBmS5ZDWL7S2PLkq6Lux5LYIeXvDneCDkUoXvo
5y3pGSVCeJWmUms712h0+9XWnt7XbXzVd5r6DRPlTECyfPt3XlhaHvLiFy5k0WK0e86rxDvkVyUF
Qe3dsQzf+oMP/H968A+xtBCcA8BCGQ2MZEutDvH61uXj4A8xd2QwIBfamrZpaFzjq3kfR84auBQE
AydD75KSXZLjwHBK8c12HqyUiBW1qrE7qfXhkEdmnWiLkwcx9gKi+hqdkVP1vXX5ln3qHvAL0Av5
tIp90SxSpYOO3kq/ZDohTAnhYxTuKHsoV/VfNnPPCmRrtOHB0oAONz8muce11YJhWog4/vGi8gYx
4vZ68oyqvFGpCY89bzv38q9E8h8X8b1efzPkmV8m04sHjQAzZX6tWYxR6vBoj8E7r7i9LpFmgsJY
FAhYCILJP+ITPrpfmqEaKOOOK0yIOEQ2QDF/7LyjJEMZaiVBCedCic6cw43p/GrSIyJam/yVqiQf
NIDUydUa1rX7S7y2NGOWHzqTR1XJBhO5bn9XhW42IkQpjte52yeKk30RRh+7br53zYHhAWcqxyUR
i0npApUuG/RJT6Mf2f8mMMS9VN07yfaUmerSmiBqSN6qfyA1cdgqOUBABMtf1VhGnRI6pFfWan1A
cW2qvrK2CM7IBxNuhrpX1n15/NvENXIjq6FZw8YkcGabFZ7Puf+VjzBNgVPSmWiCp823eDuJbO/l
qKVoQS97kf8I/WbF7tP3LrqmDvsIs7XxItIck4JBmyQkwMxjVVhKMKDuyljVAPrLGm/wzAICAq1K
DuDENh/j11ERw380RTiqzRoA/5IUR1assGUzIpSWOnal0Wq9JKKj7wSK6HGWsfThGCypLhSTKzaP
nx1cvjOYdAXsplVF2ZuEc6aQRiU3cw/PZAbgmo9GIgXbrNKJnhBJarVUXTWt04+FhdMcbTa3hlyU
ZYl1WhP+NGPvtB0cS4QluYxj5G4UuT99mi4+BdG2WfQrhrjZakuWnLPsZhJMuJI+VlksaFBVXWmF
xGU3qeSt5sVryvQDA5fY7KI3RjoTEW33BjAYI9bB1njoH05lzsrEV5V5JsDVXNIXyIFEKsfz29XN
GJHk/catSrxbLpO+czI/qijKwjXbjT6Z+RUr3frkx4K+p8q9MAU9P6ePcoJgB9H8TsMQ9WmKT/xf
jtVI/Zo45m8hp+r6J6HTkQNCJiKabBrVT/duimhYhvdsx7uhkoSKmPhdElzu1JRFFbc6vVgITy6s
ImRKc1cAcn1mt764s77Ras+vtymqxBabipaA9CsWgSM/sEjTICRmS7ZyQUAjPj+UKc0yHN+cJ3Vs
QL7p2PT+Q3BqhS4T1pOCebj2L178IXHTReANy5yVn2glxqrjNph03OQnsfRnZTOW5msuVJfZZqLE
hQJK4cx/eFTGiusv0cfCPVitLMBKX8iGzTyRmkBSLqy3lHD+0eZujkBOwmyQA1rH2LvG680lJX7p
UaQia+OpMv9Uw7Pm7Pw6M/kwBvCF8SX26nhLO2x7JTyzt4FLrZSq5jAISx2UFpwMOSse2cJ+lA5J
XLDX7MpVbTfnwwXB6d+lsDu5Em97NTQxEW9R8aA7SXZWfWIIZ/n3lSzpHcFy8HdCpeN5t/NZJ3XR
HwjdhTkZIRneBSzprpKvCyfONs0wEkKzxdKfdha3+evI2Q5S4kTPvORRO7OidreX9teJ+IuYTms1
fGZNN8Zbr3w/vkiz9SvTHNAMTCNkk3hC6XlVhbwIm7LcnF8Bk3z1R/1NtvYKSFTH3sLZ7PZho7u0
HjZyO6XfBH7oL2kEUkcA2SLHjfq9lxMFia/mWulUB6tZZu6MErCvhMwqBhbzWiEoEUhb6wKgPIwr
D+X4ETKeCmuVR52nu/HCsbcwjXoWeJQw/leqqOeoYx2P7BK4j0fkmsuVzFJs4C0GL9ohv+4UBjse
HRW54a8yjTPx99Kgsx7fQlOm3xjfT+fd52v2e2yg+yyXxOjRFz9x/COSV6gAO9SHRUq9zm7P5ZRB
hnxcxd8pSAkfMbSjivE8BPWw8bttlcFm2n4tENyXy3p13ISBw0lCOg0gi7XTaRoftRJX8vPHfo4I
1dKGxWEe11RnIonC8yxZBKf3TuwXjnnh+I/e92HLvKhtH3uXZd9d0zJ7JlJc4TCSstHTUMI/JuXy
tWwOX1E7LZ47EIQKaQVjr1TNcCyI/PyvhGf0E1hqLHF1+GmVubK1hqTbkdun1G1IjmAiYfX7t24j
CiMsf9ZLBRZLi+DCo4GJFLIgdLx9LCGZMnRwR3wnIOYELpDKvUcS3oyfh1wPMxI2Jo8FRTE3qOeD
YnEBbzHi6tPOyt8SE9J6osiaEvzDlcVdlZGvHmMi4ki51vJrgRsQb41qEgnxSaM1dBnybjbsV/gK
AMnJHyLC20TIH2rUSo21YyVVVIqQqCySMQxv+NB5peytWR5O7cEW4a5IlY6iENIGO8IWAC4BkRuK
hXCRcMADykT6xc2we7Z32ZgZUh74xdcrTGp8gGAKzSsWfvgYxPVi8d5xsmLW2GIuy8Jhnb7MXMX3
JtZs0JpGjEf64XfyCDsx82JIagXPQH7wb8eBRqPVAV6oVgtjckWiVIJvrL6vUTw0r7qcHmLr0zd9
KsxqQus34p58w4GpLebY5GclkyWuVYnRa4thrivedjFalfWu/yJbIVllW7x3LgR7uSYDBwD+hM8y
9Nmu4s/BeQBJn2z3xaB6ZefJTM7/o2kmImCcfSczLDRLmck1K1SB8azUFIrNLSxF9T3ZCcAp++H9
CKz0GBCe1PzS7lKGNSAlE5OPhPl++oR5T8g9m0+GA7WhzNGfhKKP76uZVDTNV5b1a2fQ69e+x+1R
rubX125X/MQu3S1ouRtuSPOhYVb8h0IMCCyoZkgwSgIbFxh81Vd5ZWPtOx7P+Kri/7NRW359nscx
x4ysSp1U04GSuF4tO2EMbwb7oc8FtblD6rcxQBoBaAb0yahaghmy/lhMNA1IZ3c4hxb7M3P3a2oT
E+piyQ2oJ010BXctUVaxJ32gzsLie3xZADGqkG18A62JoFssK1L4wV43HHJ9WeCNquvkCgz18okg
BnSfA41IvVQy5Oq7zsXJRs8OwED90DAHnLDTD5UNTlm1VEGEav3jr1S1mCoKQlJ7Lwvk9NjItYCX
XF30AInZkHut9RGHIgp1PKcQM2zUSnVp1H9EGfdSx434SbCoGBq7ulja0pt7wvlDhm97w3Rowu3O
YKF8PgLMudn6mSLA1pQzL4MKrS+J+JBqEyrXUWTXLXYrxXFIOxr/7qOjzC60oPf/uqSM4E/8eFvQ
DZCU+LjiPL6gxrKa2lyyVdZHDEvpF/66Y8vGDeBZkrFglOOfLsQjf0g1L/Wz5n9h9xxMo887VMyf
X353AepjBSV5vWDWZFojTe7xZZoR4HRhS4reAEVhnZNQpsvRwYw1cJ6BeuDLPBYrqFKMWaG2zXcp
50aFo2TvflO41WzwR4WKzF+ie4ez/yex/HJMgWyd+uh0z/Hi8OzCem2rmtlGJyZOGwJIL5Tbp56i
DA2kZ5IXcSRlsDXm6PJT2FJfcYgLaNjMUmSEYQXwYQqk5MHV0QWKBo0zA6Sqnq95kIVXXehVpxLK
10jZTPQqALLnkr1hpTLDxjdbk5Eh0UGiF/un33FPftUO+c4HQiPM1NAxU4JVf8ecnES9uc686R07
tDFMgZ+52BmTK2ziNza/pAT6W0dZWji4mKobqLSBq6/W6qbUW7LXf97HkczgNkWhRmR75qV30lLN
WUMZFLMdl5BXZOWpKUvBWuLDB7cJXzc1LNaE7Xa+PtCyQo6nKfZegdElagrHzgj7cDXDxZzXAfCG
7wQY61bL0DrYCZSb/aYPwigRquphYe+A+zjhC9SercMeW8ZCJlaVZ949KjIdsEO+pzuMSPiHF95m
KFGLE7bf5hqfYSjJpT4b3rtOSqh1Sz/NDDmm23C5+Ff7nddXVowFS/o0jJ9Q2In7XUiB/Jq6PcYP
T2GRi5EQ8XkSODM1fMQhA9uBE9ZiRCMJUlLH/Nu24DAzAgn3AadiMiOcMhhiYXWgfdxMheQzvecL
b2BfiWDX+yf6DaynmPTpDNrPKyn8JqPL0g7qwgZB9TLyQ781dRZ275NdBonIxcVUOhoYFG3hgzTq
vKYt7qKl4BrqjQ561SmLh5xDKquF5RBzHMO/GUg9RZpf1GT5ZKKNGThViiHxLiSXzCLyrkkPkfMw
n0OwqL/fx4TpeOrxqhSvHw0L6pBgc0kDZ1okiN/BoX9HsStktcDngl6F7o85w/qIeJa34yw6m5oW
dLzYbZtl8s1Q0zjj/dVJm354hgcnLwmYMB3D/sN8UFHlT+S6M3bn0KCP8ycO8aOpq8oOMZQaTdsB
UqcMNMfGUoDhBYzsTnMp2G4Vj3wj60WaO7ruqBc5kqbidx7we6Sda3mZggGH9XW/OYgWAjmDqqiX
emsixySx+y4aqpzThUMp7owZtZrxL9m3PgFmH6gioigi9YFOa7yf/YLkd0YAC8CoSnMTWx7C8BX+
ssGRZHZROPtQ2Gr2ITsehyiuv3mW2VC6TO6yz0c9II1u0ddqiQgIJhlc7QgHYc4HfudVqt+KiQ+E
qCni1rx8ATwsRrc2VA0AiYQYPBmMpYly0Taegf28mOTleLuFkPFVnLkVnzFmstbQt/JKwv1Rt7BG
5fLk0yz3VRa+b0DObdozYYepxhu+Umgs3LWcovS6D4LxorhoyHDOpgJdxA6v1Ldj6nZyahyxvntK
ZNWYwehG1OAOt8U+9x6WBp4tFlWFb9ikd+m4mMB2kutMNh5KktkXC3LJFp5T6YkSQmPPQ0XzWMfz
2lQcpgLv75M1hz/oLM+PJOmgQQoB0ux6AZrL66YC2YQcsD2GOM3GHDtcVLhGJH6ewVyhWYGd6O4I
Aoz2h14lmR6OmESHI4cTXGEQeyEe1zA8H34rhug+xsyGBMPqZp6wGJ0YTl/WulRAB3BltzejK9R4
TI5cJefDbM0n2tkIuakVgYEZj1brmENlKpE6vjrEiV1F/6Ej++N1SPQi1hx/oR7Dow+4wQIDmmus
SUm5UOsVdXraDV8eqV8U8AfeMYsKJqx2cyjS1qQrlx609V9v8p5VqeDLF5TMdm2K5uVUgQBK5lIJ
orFHn83afbsdA4uT1OXvyjH2baOq7LcHKnM5Y5Fp/dSp/SxibBh0Ih8+0Ju5yyLdhvkyruFMDipF
XN4AISNjNthbxBseVP62NtkOmIHHheElH2yCmjb1wO6sIA4lZ0iKtjv1eUOW6INCGJpueNLiOnMw
CX1icQMEpZQp+UJiFlATGbAvOj7O5GCaBM5d3NIZQUL+QCNUtFIhRrzGuoBAPeMUhqFoOkWqa2Q2
qFrL8wb5+D1c8/OiCscjGab9zLINOKdLczjtcAWQKwt/r9ISDqp56pGdWIRIuEZi+2P65m3pQOH9
1zVHTq/lz9HCIh8w2MgOENnOj7E2/SiCtpNwHIE2W/aEqZozmghMzI3SeHVmyq9zVwwVwy/bHPT3
EDmjMfr7a1cb781Sj3DW1qGFgVXs3JdUhWh6oETZ5cyMAyj63k6Kb0hMIPDVnOTYtGdoeoXLmV/H
AgHmZmVvPDo5EkxNpdXSd/g+W6AaWJXma+fzKi5hVAvAzXRFTp2q+xE3jMLbXS39WHuDiYwBjt4r
0ENS10NSuds9wsr4rpseo51/UO+1n7MyAQy/6TiTYUAEBChlnoKU331bX4OCR+DQ8o3ZSVPNSKlR
uVTtgj1ngvHGZad7c1OB63002sh4ops0LCS4IoXzoYu+ENpGso266j/5E+CBhj/DZNugzIHR8IgI
ex4GMSQQtEefLwSKgbqZ1f2Vi9Iso8Kpyl0sev09Ee14pY7vGgw9bQJOp6BRyNxcj8hhjesZmIw6
4NCMBX+42qt/JFA+luLtuYXSM6giTDCBWJh6jnAFFhPMyJ0YbpbXDiXiYDBCcqfxAmcnopahX0Ec
lhAwUOiQADjO+IxUaKoh1UpxawoPQk1Wq6mgtb651gLYNXZaQhxDMT/9Q1e7QDAULUiXaaUefR9I
Vc2ECBuY2+Jvap+bMbdsfde4VKWVW2XF43A4DSQtqMukcVb+tiGeUEgP4Ut6scHP8KSpi/j5VAgA
5qDQnyRPJBCD0AqlRSAslcvxouQxK/h5lP7h6ADEXjz0iDubjqimIXVQMP+kXysWMRQkqk1GG6q0
de9PPSPqywO4D1+0vFPK/oawI+cmK8bcXKN0xxvyfosou1x4XLsHFQaBN7neG9WNAYJBIWE9TAeg
vmvYmtgh0TCMlaZblmzfM+YjLE29O+2BsJqHLgZ7Btqe03PVAAZitB216N4SshxiAJuDt8/KPAf7
2LWNg4oFCQywI28+BUogjXrXh2pmq7LDlZlibkz00LZnLEGSBWUp9kGw5GzqYmJZ7Z/xTYwZqq5w
LgoWc33b5wxIQ56sJ9pGo6SCPEyk3psOytxnlsWDO4EjOGDruumepLwmO9WPJeD/KkTNLinZG5tV
Fa6Dvuq+VtiyUWJ+UQtCJsIjmtAe1so9NIRCikRWuBm3s9SNb0gUVeT82nL2s/Xyc9b4SPjhjnb7
k20VO24Mx4XQYFHDlPfaoOg3rt7jM4DIV2th9cGhpMqh9/W5alpr701YMtopVS/nFCDUFDOYHqki
rWRNkQMGRXcsvQRTp8DWRF6PV9FVgUckIufBhD7HD9jwiYdK1iMaLa7DgnoV6B0vTNrcahVIBUtP
vKblPsuA9H4x7+CuERzdSWkpVcWCTdH99TJMh8a87hX6k6yXsv91KUUmGwaZU2Y1rr9M5U6TyH4J
V0N/rtHBqdWSqcInn5hWM1dASdb2HBdbOqosSTsUp51E9m8Aq9kFkvANq3BpePsvrn1Jem2/OIhF
G1knKoNrbGyrPqaUqHF+9YGSfKrCS0E3lw42lVU+cp04H55NZgXVNff1HkWjHc7q9oZLjIVg8KCx
9ZLI28XaHq0zS2iC/y2NY2GwkoMmz9AZsSHtB4RL3UymV5hGvFOF4bybFpZOZqEHITjqSYi1PcF1
/59dWUyQobJ1Rkyb+CBQprW5j+61ZrU5KfBmllU/a0RFUaPOW2xb79/5iTM8X8oAEzEmgQM5wGYg
mpFiIg69VJjTn1ub+8HpMnui54qwy7TMCe4DlmZW3w8ZYhFtSAcOKO0ZiE+pwuwNZtmDVsAohxDO
3N2OkOKmw8VsfJKAgeZLvplFlRT6Pbri+fyLhNm35BjCw6hMFrCxNYlqLoq8G+ojj7kcX+9YQCy2
FUX8/VRSQaldpi/1aJjM3CEJs9fLCUAd6ZJVwo39A29EnlvyHtpYLbtiqVUqlacpMExKGhy1xDDO
hcVstaN65I1jIgRvgZErTNHfrmJDZLBk0GwReZqzyhWx8zSo5K5yhDktoEZsZ3BWAnBnTvMukj78
n/zmkkKuB4tMq+8V+Mjzt8sThLuU2g/rCm5tOkbuwETi+2f6Gl6lCsKqmiIB6anZjr+6JuIM5HgM
mA8vNVL2bHAu+T8gYI7jjnFh9j1VGFpmgYt2F9MFH5EXi7mrN7R8zBlxRSSVpUdUGP5su5uyCGS7
FGg+ttds8/jAX0TveODJrhiLJtz3poBDFPm10RMWD/lquTiRlx0i9FYtowXToCmeTP4RgxHtJ/wK
XvqSwFcOIEML1R7JC0HJbCDtwg8AwYj2vvsSCEIxEOLNA0etqQoAMYbQ5RZeZXJMEFzi2ussZ0bN
bEecRAI5MrhE9djb+5CQ3H7k4PbIlNxWmMQpRGx31qsOzVF1SeodwIzz3Ibk5rOWivWj6gyguX2b
F1kmszY0a9ATdwCIuADzMz52KN43xVlZVb1azV3coSpyPS8UaIlWOwOd23/ja2pQZcdgI5GlDNqi
6CA96bTh3BaT3DwXFyxa0YtyAHK3oM/zwt120WD7SLeyu4wa7GFk847/vnjnP+UQ9SxFYDNeE4xv
t52ZCup9++6bAHvBs+A1VF9n0eGOA0SSDB40NQ7gWS+jmi12ZELJpkfiRnjTMITDoGcQYHRm7Q5T
TbCyPVMsUBvr9wADrXZQDPFOVwyHc+MkC8sAuprCkx+U99r5delgzSJ0JITO/QtK6L2vJRMlSQCG
SgfcpuEiNKRtLBE/QcNXo/RGcIDfb9X6vEgjAe/xTs0PplI5ZDA9pMr/pgXmFtxByKTZaothSyJu
1jXg3nJY8eSJ+ZRme27x9ymNrclGPUIeNIBu4rCDRPqRt8MRUrGKu+kja2xvcKKU7eyCl2D+sjZz
MGDNN7MC4jVC3gCBaIbPCEVqP+J0tyxP9JENC1+T0Zn7JnIjSrNyxUeW8O2sRzikmm07n5Aa2Bxm
BzrEFSGCCwpcz9teel7zIEbLCHlA0zpUkwHfkn8oYru7mTK7+tLJirAeFL8a+ySa25PNVnE8lHHJ
Gcc3w/w3nI/cd/iml/jU2aIDz2lvjvLtGSt5OHMO9k+dAFERuWcbRAgPJMHB7PN26mVVDqwtCoxl
/IcyTh74oIx64x7SBUAwrbJFUC4ojBwDam8oT4wY7nbhk3oxILUEZs5GeIhxk36KIxZJcva9Pxk/
Mc2w7Y+soUtHQgJAAPV3kjwRke3f7CkajilWTrVj0agjLnx5JLKn9pHvlnw/W+3DvyQQB/tSJvLT
1Nqt3W0Zpf86FNYm9O2nDG5EdZ8hKyrCmsOg1rUz9jZberADhK1Zrbb366MEYhRQhAzdKEKrTEJR
fF8mgKP53QaHt/W+7LqS9DDn+jKXky5A8VDnaRXThiU7D4+oiqp5CccgKf/ywh8fqrORVaO1VEiz
A6mMr1dyyKERLYtFL2WeKsARPrWH/LPRwMJCJa9M7A3IkrPTeDRodTea5A5a1nlbVCCnG3sQTLUI
jp4I9R0+56ylVZ3pbEG92IbsE/PjjgTV4A0U56YltDtU6ehYupelXk89SUkNBhQftdrFs1nd1qa8
XWBuUhEH8rMQh21VWZu0R4YtErQFzpDsBmcZGNakmoecsiSmVhY0r6uX4vOZXQCFa1wwhhUZL7uF
ZY7i4ttfTE2It7X6fFkyaAjameViQAOHL3tsfehnbvN/TUknn9tg/iMdOiS87npurG4jhI64SaCh
U1JS+o7iinpz3XDxRugTQm6/a2puH2KyM1iS5/z7rW1aKNJscL3ioRxaow2gH3RHhh34hF6nW9g3
kZCAQZm5C2Z6gnBPi4HpwL2/9SWHqJdVKLL+5fbIfFRs3eE8Z6WLtwuDzi2C35UKfF/GlmuTFRAu
C+RMJN34ZSx5Wya8ImdUvniHgi66qV8/P6GKmc4sp4R33cpKRGYpdsh7HqxqWpEyr/dsoDvBG6K8
Gd+0esalKegoSqEbRv74CifHLvQLz7Q9UFW/dFqw9mDEtRl+lEKQWwW9aetFqEuMesLaeJUnpya/
nz+aY99PvPIQ3UR3HnGW6DgqDGje5dN6oHXBsDr4NikbE4J7C3qQS6NwVNkGdTOSgEiTosBS1DU5
Mc+4or+6ts7p5DQXkUQNHpZ4q/PYa/gF4Y7cJbuRE5EPH/W/MptSVLqifUpsQktw4FQ0su+9d11K
phoW+UvoE4WCeTrliHCvBNjdj7vR/8c8LrGHo4IJA96YbAV8BhAfC03i14whmgwJsijbaBDUpWT3
Pd3IqUV3F5+zoKyOawLhenLDQF3h6uR8AJ8AcLcBr6YRyzvkQscfjxVVaAeS7G1v7NI25p+a25aq
TbJWSOvErYKsvW9RzRFPeM4M2yutvOc63F1SzYTpxUXzGQis1a8ScaTR6kvtEeusMZntsG4WvVmQ
v6PS1spF6EDaVH5AEAIuoo+J84Qz7qu+m4jLzlvIAMeYuztMICRHuVKekU/LuGr3zaeTDQuv/8or
YzOpc5a3yofZr0+jmg7iaRkXV2vznakfZzkwM1jNqz+cFioAfNvRejxkYKGTZR12ciLcDCC9JPNT
hOxinGwGAVXlGFvbDaZnxTfmq8TpFeirez2j0UnOzPuyg1qNMV8iPW2Rr74B9dyac/NyxkUK1sAs
PliZu4wUfuOn0jIDt+5hvdKG0EsDojncy/VGMAxkx7KaY1o7SkmrDPkx2I4DjErO05UsTh6kG9oi
hTm2v5tos39+BqnVvNwjl90FN65Uo6Pj3LKkjjOzdMHq61ossUDJ2wMQ17K1bWxsVenrgqxzSLmw
ap6ZMEMniHvBqQw5xgK8ooan5jW9Zp78av3XpEwcNg1EAo+UeV09UMYrWN8oEcBIz8dsIsxLeE3+
5dN0JxGMQ45Rago7VGiV5QxGxEoVhxDYXXhuYuFCJl3ouGMq0aJLM+78T37jzg6N0bn4ejq01SlW
J8g4ny5EsP+zk5Uq6rh33BhMknnLVobYyFPlGqceTYR5ySDnWDlo0Uzng6p760EGzfNwK9sIjbJc
/pHHD2p7l1i+8DrOkxroA9pON+uRK4B+LWA7qMVDa+AzngM21HNWtA+85Y8ZkOyQ7VuIoCu4YjZZ
/ZbyXAfBJi/Jsq8DLDWIkej3HEHyYfmM68zIye8mLLN8Ea8SnBtOtszNqdhIqXYPUonPivoszO57
GBW62sAUGUTRXoBthPd5c6/ungtWQURjqg38eaB93FVIIGQ/YRVvbDYtOPc/WcIC/LJEablFHLyX
F6rlpwd+Jv7+ZorxD1ticjFKE3YC9RW+YOWmnjzCm3Z3Rs+RqhG1fzrsYRxTkrWq9QWy6yFyECDk
xtiiu7A3VGtbhN5OQIJOzyXvaX8Dwv6fy60e9CPohc1X8+FVBH0faDG12QN3jz6tjq/xhE1jtZb8
rf+7hT4zCglsHXI5E7CCfEkUP+LOxQZIu4XUMs0jSt6KUkJ0oAWOqx0+nObqeHOuf4IVAj/2IA6c
x+LYtlUvm3KpKR6PYd32iK5BnB6GeJ7THzKURqnMjffDfBUnket6ru8cv6dkReeWOpVQQtHcN+/Q
Z0VMQ7B07zo0x3EASCrA/5SC/pOeKjs1jKKGvtDrM2zTvI0UNGuiZEW9k/yg+foGe3B41AhxpGX/
D0IR9Z7q8yER+DPDMs7nhoDmv7fednfKClvNJ6sLwByROjOnCVlijlTPesvBTqwDh6lTJKzObGhk
wuqyvMPXhOcBXZ8IygHPWuWqVNs8MB1pJBQoiO9DPbmbXYLm6NrKW0FlkYRGlX3bSShRx6msDWLg
lilO8Gc0HLmHRz0nx1ol0xoraMhCHR/P9YSjqypJNgo8G85UnqK47OjWm6ZtM7+593tGVjqthvk7
dHNa6ns7eCtxNpQKfon1QLhCMXup5mHCzlm+xCNkAH1C5u589ny8Pbdbs+cJX8917hlfe2bAOiDd
d0xRJzXMSqbcU8GHIS4/IWb1uQsjIqBvDJr+iqq8VnY0NlddubRRlSwOS8WxsNZFEWtnUZ2JDwvf
MmjO35G4OlNESCF5KNytmCYYr5/c40pfn1gojtlGaJM2D3HhFAhz0lQ3nk2Ct0YHBDTi/WZIs02u
vkK3/qWd7Yek9ArM59p8ssnSwEW5yIUr9BYHT2FjBcMMmVB/6qVY37nPfkj/G48Sc2mvMm/ObM23
Mg3kfx/sdx/JWIZzB+MVwLgORKDvgo2RaoKzxE64mvaLvigRu9k7Cmt/NniquUqXmt+0nvQctKKw
2xxeK4f61oMlM1FzYtVks1FmpC3N75N4EKuZdttvB96omVtDXj3TWRm6DYJ5RK9OKs7lHUkdygg1
IE7ypCUTloM70NSqBy7+Y537604LhPoRWqB7FMpa4Ud8jy74rRLGfx2pZ8kbdxHyfSRb56e4dVkC
5xm4ehDWdW6ASCyAqDv5DuPG/REHfYhfZjRffQHUvg+a6macAYPrbpdW7rsk7dYWSnspFq+miiD/
uZ10etafClmm3SG0gwsXlg5rqi4GF0wXy86R0UbI2yiSanIgZdVI8hrazsG4G2lN9mJPxSaXURIg
8cXVH8x25Il17PXfgGwe265IbU4ys7OToQHvLYEzGfWkBxk0vc4dkVPERryhOtzZwemH28nAwrPm
urzmC4Z7fprp7b51pBaFfRJc94WMzibtnykWjtbZi6al9NX5Fk9XbBXaWKiTvcyRiPwtMwF0SETq
ngh6liO86+wsn42Elg0Pk/YH9yk7RjdCqW1McHwGixo/f/JGpk69DN2DKeXkQZ/DfNDTYWl+r7ia
J3Ij4owDoKZwYFi87NMILop3owCVdnUAp0jvSDu2skCUBx/cJK6jXVJ1zUpBgRTDK/xLa4VtqzI7
8jQoqbRQGVSfWpmcpd9i9STBhdUVI5DUrg0zfUZC9ZozqBInjDiXZUNIFjx12efF3L6YEu6zjAm3
QSAeVTx1sH3H26t+bH5pGh3iWDdumQGHtf6Cq2kzyCYC3EdB4FkLeimuK6+9ATY1MjPfECgEqj10
Y4weO0oQkUgVH8246+xu1bG4lbnIEgqjTndQn/UghOO736UnaQxT2tzgeEp+6uaci6dUs8/seUun
ISr01QmTRGX4aiRC+qEiYJKt9ur95HOEU7SyTBUFSFqkPfoVdxlzfDgSDzuK4GyEAz2gzjVp9T4X
HRmPTKdsClAajgi1lUnBsv+/8GPQkqnIcpn1Kan0LsJrYTrFYxwHPQdgZpZ5KTpCHbK7/INP7KJn
A/ERh5ZG5XDCtlk3UagVMzfktWtIrDnCYtigKZcyj8FlBfntXWSiZCoS1V25fWsUCxrSRQhUwX+v
sA5AG4tzjCZxT2BPjL7wg9Onjej4vQRYMBxQUACVZRFwbFyyBW0atFTTuPQMQwvbxGFpGbwGBbfK
FzdZDHp1MYjDVUQHIXONDzwjj6SafO9TGsynuNFlJFHOCS5bN+sSnFG7/0byDKZOE9y7na7tBxbm
aAUv9zul4KY62RA/XfKi2CN+alq2x1qLLQSXPwMj4d6WkqaN+yRYXg33cJrRTv6OQmVUofvzxC9q
egRCOfrZGLFlRFJXvu7QrRhU0184bCOlmLKc9ZOD/wqR4MQ8zVUCiiXmbLQJvxY1e3e+prSq3i0I
n4mmG72VRpV44KHesZ4sQeTMJS4YIgqmzzUED43+1A+ApvoE8k5owCyCLKsXkXE4F9PUtQBzp59m
MZOaU+2tonW8rJ9ETGXwJlQYaA9SYHLbIAuoU5PMmJWH39o+XG8xVYTEzJGOUM2jX4WL9N041Nu/
arljhXmV6e8dcfu2mjo5GOpPJoaFOVXgQ+72gUWOfEcW4m+9Wn8IkOm6JTU4pd3X1Uo7vexTnbhu
RVjo/H6SdIJCdfyH4zJ5MbCQHyxWViJ15RjDLya6nGhyd9lXCUffjqTSpVg4kaS7/gzKECrDFvHv
Eth/IGd8uPQorU4JKflrO85RH+7NJ/rsZy/sbrS5uhXv0pF4/RXEzM6k8s2J6g01/N9aAB7dhVsy
L049q2WYfS8D5WcvWUo6pwTHO7oTnTInO2aMBjrntYQnsw898FILRv9BNGQLaQzMqa8JbhpVyP1L
b42pPUzcts2boSChjAeFfmvmvBZ7tF6t1uqdddQeyT7F+34OvkaIUPpFiddgsqVl7UJPVAAX2Qy2
RZDd9t24RpyvY6Zi9COak0fD6zIWhhw+7WD6gw75qlZ2jM6Rzok81ED5l42hMJkMFe0FSuWlUYHb
azk4+dPY6+jrTN0BfZlUxSw6tY/Q1haibJOrt4jmU71qyRBZAetFVJ0rxWy+nsGPowKs86yE2r6B
WthDIlVsAhcs12hfBj871OsXKdzGmsdmKeooVTIJQluJGlfXp9776ztLypbnHuSoCt1zrxoXwykg
xU2axdKNg+IkD0YCutDUnv0kXgQZysTLJmtMSIj55pc3a+fWf6H3seH5fgCR7usNuIzo4cfZqcRw
FzxNlI3cO7IaqaS9nfWHBf4cgTsZEER/P0EOZK8u8oVXcP4oL10uozyPoyhlWc0oLP9n2xJgMNld
p1rKYBIMjz6ACKWFNfL1Ci4nm3F/xcMy5gQa2+Qq1wKDz/CLaKG79Tr0OnHz9/5h5SEilgW6FI0L
D81dBUzEzGk2aaVB+RGi9kGep/3ScOMSkZm2W8uA4Y9MM5fPexweQPmgHHicAhMzLg8xSihp5cGA
XhXOyA6zNQ8EW60RpnPhwpUM5zT7jtBJ1/uWEGiOMbOsBGGZ+ol3pa6FrMS/gMT3YnqFeW8sKiGO
eAdAiNPlvyvX1wTKnPdIuikPGSjPBT81JI/sKSCb2dTUhUK4ot++Y5ycOk1ftaGifCFyxB9GmIzS
PDRl2bgZiqFmDZVGixDRHaNobf49x8Y0iJxKQ0+R3cQydLyaO7eumkS0KBSW2uqNZxBlJUYHmZ5R
WrVUEgXL2XBEu+laBKzCHc9I0Zjr/WvnyvUJa+XZObLII8Q54lpG13SoBQIPDKuOlS0vx1q7Vlyr
0Gje7En0jhS990Uz0w/oenXpMAHRPXVHN32p/Ee01ewBoE1y9U+goSnbk0hxu7eXlOK/Yd1oO0b1
wSxaFAcP6BptNrmyJpJ2Qt4mBOYy37XNUmesP6zkYPIUn6u3VwN0m4HWEUuaQtq99d/sNqKF1qqW
u1hsT70KT9/NyISnfYXZb/6lgHl1Cry+zPPu8NAYGg/QdfG8eqCxiIPmjn7+4BniFIKnkg2xnFhQ
uyT7qrxhMPG9MhueA+ghPIwnzMVN2ZAbYFPscyP0RUHzyUFZ94WgQ39x/7y828WBdX2x4Wdi2kPb
wtWMVD3wlIItQv60yQJtvyeGYnbxPItU99TNYl+kkXdt6HJysYhpgZLfI9U8SOxVTwrqZBzrSQPp
O95lyXIsruusj1vW4sct6GIdI4g2UXw/6bBEF0wDU7REcb3Masx2oKiXW9apAgWZpCJaE8cISrc6
cpf3YXdBGel+FZI6Bs1E23kKGG2y/HYrqdCkpRCwbbQLNqfJ/DfmOagDnWq9z5OLClsI0RY1hiKy
eCsNPOTm1k21FlVtby6bpRLHLmPBrZGqSf1ibAOWVHklM4bkyPb9SQtRdzKVKULvcs6O0/5WtXZ4
7MSUp5jKttxsCAI2sO+KVQb3XHPcizBG4rXQSww0gBXdwZ2PsMLNJ756FXZWlTf/hnqZejEczVub
2B34O85w5JFsjPVJaImz6woREUzHIrICeXRHWBh0QdabDhpTtPkim8zTpEw1YbQAwgud9RLkqWN3
ex1QWxf2brFnLXaykCYxYWmbAmSy3ZsDmLeiqJTI5mA/aOGAgL/dAHN0TTnddY5NcMp1h3LjQAg8
Qg2CqfWsd2KEkHgFlgN2vpYbMI1ZvRSnQouep2SIX3y+uw1bwRKL8PQl77p0TxTuU1N3BBno0HDe
IJwydGv23sdE+Eb0gdRMS3dbN1NMYweng4zdd7e3LM3fML+x7Cb+lQsU42UFie/z4ysT60qy77Yr
VlpZWn87rwkniZdEwoS17GKJN8Mt82PrLvkeaf0E69vNkiuca3Sv3iqJCjqSTEchCTbZxYdaZoVQ
iIucPajFF76SUFtxja9bBETClGXcdzQzZ6+JT+fNF470HaPJauz8chd+wZGtiTshGSGVVBW5nHmQ
pOYWoZY5obVQkIw9SupwmhQYbq+xn1Umm5GukzfM/CLzY/TU7Cdst3JTowB6SMupId+NEKkL3PkP
4jRHxThVI7zTAhAfPTMI6gWBxWS3TqEfL8IxCUg8P93rRcB3JgMiElOwgRfmnvj641PoKsU9lO7n
n87Xky/fooAieci7bPYWlwXWqoXf/Z0c4YIMbYDqvwl3a9NXoMSuWS+GZBCpYnGT+08Cq7w4fr/B
sxJ1BXt3bWqNRfes7DkDcaLhmFTdqXAR8sXjP069wH1Qk6Mkn4HJIeHrB/nrs4+EFY+nH0wAJtqF
2I28XN9GYUMRF4eHbzR7slCAOLt0aSvUGJDsMJsZxFC47g8pMy3t+dkJ3Da+XT6ZN4aalW2DZ4AN
bXE8DNAMIDp67sr58d6praTtNbYyUjaWkv0DZ5osSqfB6R8Nr+1qjCj7M2vjputmzLNiPzpbLfKB
wRzBErFmsMmHT04HCcKE4jGo8U2SMzeD3SXIissZKQi7PRDk6ft8/oCkBjgNmgvlvJ27ducSgz1E
KE7P7DhlYNttNYUTWFVNXjDrrLG4on8l7R6AvuIIftKhjDGNf7EZVAtyOWob8R+FxDsHPXph4PJP
/Qp7A2LAgb4mG3KSl6VgBYdX3jSjM1729WRciTg6nKI/octRLJyeljNEiH1yoterFse5PUC792uT
GHnK1iwr4x+HmH2h9nGlS7W5rMlBigdcIz5C4W6fwYo7uHQaBYoa1I22vJyFCbC6iw6zErCkyWxh
0i+CSiBUy0uB49uciQ4R9vodnieIfBWp/IaufGnjTRgFspry7/xaHgYhZgivC6U2/OCh6qlrY8aE
Z8sS5tusc+qCuGQObBz2ZnapUzAwRpQQuxNjBLNURmN1v7u9k1VvugV2FJ6WPKz615qe4PU7isS3
fRDW4VUgMUgJ9DVOyVUxz328Wl+xEUx40Vap37L43WtE36TnnT/iwj26rP9ZMMzbNKqkfCCcASQR
uccFLNt/kR0qhf6I1CX+07/N2Ku7F2K9qt7YKzOpvhe2nCQSE6XLo342uOyIhUoWjQ3xzlmV3Oa9
EPoBfbfETr2WqZlf8JuQHRcnGt9QU3GJ8CbEueTJRMA9zH1CwGKVLW4FolV6ypney2+qiVFcs58l
3PABPlk+KSzl9Gh8ix5exWXYmeKCasl36RL3ysr8C7UVpD8j4y2ytLbpj22OchEGk/MZvvcaimC+
ToKiUPkaXIeYxcVgiCMz8vRsF1BZMku6S/MzUwMOmm6YPYHAJ4fgJ4N/2nnWk4p7zrBOEWX7VfKC
TveHoImC8gvHd1uENHJ8xGiL9KBD83f7k/j1bTIPJCmqzamuOl9Rvvjdjmn9AX0QPeFI/UCDu4ul
7spdYByTxMYA/XMvPazHCzxMrnV8a/FcTzWQoLVqevZvXTp+tEpNRDmE00fL5mxuHSsiYHVw1yt9
qE6XCTnV3mWu27gDxsofM/KfwDjT1OB9IWO5oSzFg4siV8XQhdLAZtn1PZm4vnBGHInd1/opqeBR
hxJvdP2Tv48/7x7rRvRTvEnlg7FBHsatdsLEPQjCtW2dvLKgwzeUDaGBdgA4srsI+mJcVr/3voil
VgVmghEqeeo+yCrF2wilin5hbx9OaOVwAbO28YYHO2nF4udMGTTNQgCChZgOp2Hm076GXhGkOleL
hqXjjjA+dBZKsyJHJnciUan2d4n4T5sIwJA1odIf31HkM4HY0EjnGS174phFsuQxxfK3mkkeCaYn
jqHbs95Yq7z3WilQHE052AgkyvMamLfC5EPsHsq9y3GpsmIV7HWO2U/UM8jlrac2DWJPwaM5Wzme
b3vpeb9qbh0SIH8UcJlDKN/Vmqe+hTR8O4yHLra5sTi9ZWT7y9Hph5rCxGjwY2GRyVkBZlvAqsh9
g4rhIzCxs/QSr9oJzzUCPgmv5cYyREebQlkuM6Y+I0Q4USCtzdc0Kedcc+MCd0jnFljMLX6SoY4R
AAG8Sj980oCC7h5nkHiQd76b2Px1Xhv2SY1E0c3rgvyyWn0uEwNHeHyQI/QRc8iWWD2Rbiha6YHW
dPNTpik8AfHCftRGhBdAuPyA1o0aes+X1LSvQ3ueZ+G+mTp7h8gTCVliykoZ6ng84mPl4QmbgmEx
ZnwcEtDASyKJOYWVb0loG5hbR/m8r/R71xilGI9IghRTC0QNoy6WIj4yI0bf7aB+vLWpXKyDbBBf
T3rO9jKCEH4EpRkUnDffNfqcnoOU221FtiOl7aseYOUpWGSLKzkzcH7vCpIDQjWb4GyyvBGsuy5L
cDmuSiNRKMM6r+/lreNZPdulCAALBJmGWp+dIZrqqiPDCSWVbc0ZST3M8AMWHBEs9uzUryOOK1iH
piYpN3h2zplVUKvFOfCTAMcmmxL1SiyKpBfuG1dOuofk1Xh4uQvbV6QIFnyLf3ye2lhhYaxSb8dq
rdFpjWRGEHds0YKrMkRTLox+mDAnkW0whE/DsJmsuKlrFLUARmyYh9tVf0GWVn64AQoNCQecbqig
ZoQXGPW0fTGiMKR7/2JOGwt9FUf2B1q5RQ6pYsaWlY9SxblYyEG/Nb7LoRT5ItdzUivDs1epUKCc
SMUusZfONG3jGpZtFywf/PAJPlEDSguIK3aOA5EOGLGmvWUDag4V6Cxlyt4rY63rpWZiDjyRRs64
HNvAR1KTnXhchI8xPbt5hpvDWIoEjENI2pL3/ZS3XAJaw5nQEs1VcQhvH60RRtSPqMbmB7DBPMYd
lw4IHp3fcOgwzki7grcHE7D/qwnY8j3EqJzqqnI/iYlxBySeklS+fTonFpiBYD1y8l6Pu7YCZMZD
unL4NPBMHSIxFcnp82Wgr8Bv4/qNgoY/Gs2322D4QxNM2GyNDkINo4QDt9+cCq3Q1a1UPEhl6nX4
p3TPoQr20DaVOftwAdmpXxHsByZAXlScDPVZe1uugfZbvh0drBBWl0egTK/5sdz4QlCAdQwsRJ5y
K3/FNZqsO8MCsn6y7Cg7TYmJtlst7Mhoi01wNlC7yZweCoY4KSQn70E1pD2tUu5LD3SpSs4QBoYk
QAQrNzSphs/6DqInfHgI5wIXYwshtnVkBU0A3KOl6zDzlojN8Cd0bQo+sfYVE2ndfC2VM7u/IGkA
FJ5quTN0omOLWfkzWUVWb2xljn29SkOGwFo/z03J5v+DS8xlwRsVf9CGiFvCdptN7ntcO8SwwonH
bnZsQbsxasV5vsXkNOx3VizasGDEYlRarZ3BEZ6LZQnlnZ7DYS+/bQerVHByE6hqezTv000/irx/
zq5Ytjxku7AIyqGviM60xJuOtQ8E86eI2ZZ1C04OpNB3JQK8TmrEmczg7LWc/qC/RiMKj6nLTH2N
DLwO/F8w6KIsS23O99q+RO6rgOmd0MsZPr7ZwxcJNaeEVo4g/0Jl1u7lXRlex8UJBS2SOF5AagK/
jVRAgxGtLzShEQDlceDmBSrx9sq+K3f+8fQD0HzS9JSNbjuC6zpIECi9St48mBXMwXaV/JhzL7+f
jXQ1hseuC77B5Afq8KdqMYWeUgcLjcaRpLSjlzt1m2WIQ1vOIbl4R6ljTBzakCSSrh2B69HrytNO
LnyMFeNsAF1v6+cdRHTJ82ww6Yfqfr+x6lCDrReTyY5ZvTCJAUAnEb0I9dom3o2PZZEKnANuvkqs
To9+K+8wxYotidY2vbUkyz8XQa+cy3UkzsWdr2n5ZRf4VNcFGkIRnB39Sp0VA1Msoe+XliczAi1D
lYLgdDbXJlS6z3S+EvHVAT7Jv0skJnky+mJGWhGbGw5NwECA7sbUnu3WwR/UhmYc6/L9qcfZsDix
GLVfpZmDTrITXM4cPFrA5JBF9XOPbh3PrME/9KMkPginj6GBdEzKYhSTikiw8xcmHtM9cv6/oOp0
BSOk9xZ06pbNAR3vefg8FqvXjVr4fAuu3eBgKMSCSEl/N4kJfARKrapdmvzvpj2CYuL/ZeV+O6jA
Mee15HaLQ1nFYktbKyD//8Qhnn1fsVEOuHxmaqIOrvCt7KO+j6IiLwwMjhPLQq54ZzJbFiU9URNr
Rt7knS6T8cyUk6UKgv2FdfsFEs7sPbu+HrOgiK+y/pPFxweHyh8omBHn3A1dAGDMRka9RUmmx8+E
StXYG99atY5MXjW61oI632EhDwCh3o5SAEzavD/c2KDB4deiXH68Ij7l8jskE7MiSAtKkdOG5e0b
skv5JDT5hmOsDtKuWYq59fvEoTVEUNGZeXrsz/uyc/fZGxAVfnLw921yex/Q7MuDAgi5mA9tldJF
5UPyrlOoJzvw5qvrQQHi6rTiN0nEa6rIeloRCapid8ScvQvw87f/FC55QqsQfc2AAV/HJ2hPORWS
lH8BIlG8dOvCQZMKDi5qETTQ/HCtg8BcN/1V6Dr1ehnvVpdz+5T0njqnhidJfgPztaVYu3sNo3Xh
GRK2TwjP6TLlWur6ccMsxyxY+FXFWmCgLVMC8FUaAu5EiCKzCAdIMsq7UamGJxBBewhvw0N3bNll
8GKb5vAVeQHJlcr7AzMpCx7bNn2b0W+4OIOA8xxooTQ3jhsqUkzpLVx0GTs4UJ2ny1jZrxkYSrbo
VoAW2Hoko9ql4+nc3h4uaC0lCprbzoSUD9lfgVsO25GKG/zLcf+CP81ZsVRsyY0EAIa37hE1MvZS
ItERhuG8vFADHJ+STpk53ACdoF9K6sr2/y3OhraabEYhJULBTOX+ahLUr/mwdtlE0LwDSbBQzuye
VOVrLPBiHXhb6MycgDbXKjiIs/cq5H9Nx2/sUvK5Kphy95DtOQRPspmntaWv7S1FLzI84FPL9h64
pJPNqFkeItznsaAf+QjPuDqTm+TqUYliV2W/Gjccxa5Nb6T9steslxZQKqozpTHyQLlBJhHLIN6k
VLSkRk31UWFbmwCNl0gKy6VcgLQ7KVHV4cigGDNiHwVygAoDGTtF6jHBdoXIYWIrEGiyJEQS+W/u
cPbpjxcMdnktcG4U0APvYAWLiF3i8+KUDqzrIzb/wfKSoJ29nC4/whH03mdFqBE4ClB49pF/9Oyy
Xuc+BGT0HlyasLHpsXHbUr8LonqB84G9xx7aSDEDMz3GeXcyOxiV/+qoBUkaCeZ1KJXCT57QxVjk
g+LqKjtVJwoYP1b8vjOZB9fo7Wqh7LouYpg3vzLxIXfUDGZc2KjterSGg23rBXop4tk4+HIHaXH7
ABSpRPTVMSAE0IFzZ5Je3AZ22zIRwS8Ye6O4HpoXhTSHjNqGk1ZIXwmuuFu6/sYls0egO4k6bART
7w+vY6UoO+150oAJ8gvTqRAjEnW+hdwaYOEoov9kEltZyDQATzIkCMD91Pdu+FIumYHoCEzVPf7N
/iCuZLbDxow139nU8rtr9A8B4hQoftiPPln66mamti35od1/fdDiu85tIuOTSv/eqgw6oMIz057y
oNAYSe7ee8sduZ0AJ5mNlEu8S/khWXeMpj5LkHHL4gez5cvXVnt2aRB/u0TjITVo53L5S5JOO47c
XdQ0yoMm/+9uvmrs2O7GtYNbOOH8PA+2UsJI1hWgxr+SvvgBn5n6o36BqwNFIMyldLXyoWKbq5sb
lgeAchlq4Z1zlM0ASnOhNAVrAznmaA8ejoqH4q9tMipCZ5j4O4HnjXtUT5eoZ4/Vsyq3z/8NHZZY
ZdXoqB7F5YvAejmlucEuohdn00F2GOeUiLDShfxWEQ+zJxaJrLDrskreyGsg/CiHN9xvu45fmjeo
3chK9K/ONLjmxQpIsr1Qx3tfgRvMXEe03KAyvl+PRdwTP4nmyZKAkcZFNopyOM3QVceEDXqvmy5T
9pZ1SYqcEgYMbkzH0F0eAGQOdAg/QI6RrXnG/cgjspUrPFH5Azt9AIjh1PP9K7IBOxfJ1MUvj3H+
+MLjEWwya08eNX2GK3O65NlYp5ayh1L/IGz4ghRYpES7yArdS80Ym6P91JDeRF1azr5r42IjPqB7
pRdFMbKHI7NwbouuOZQ0XlJr5Nwxr6j4Hj54Jt1LoWWEfSL5gsLi9UdrR9MvDdBGUFDYrTm8NvUK
t+wDsbKvax+Z8+jXPawBDh7CJVv41kBkl6l6vODV/K7zUccGLTSFSYERXWAMea6WplaWobnCV2m+
Zx2dAo8eMv2kLBvYnrLfQ2jMrtHfzvQnBbRbdX9LTxaCZQc7mQwfN9Bhale2ThsENit5ZBOHEtJm
jGNTQWKYfO+sfAuxwEmYfzXkh5vir87S6TkpkWnSLCdUAEF2IjLPlTJQwYnTXF93O7MdqdrxIYje
g2oTZEDwyOuurDQyWH0+ybS/FHX3hrcbhquikMBdEf5PrlxFjUIZ81h+ogVwcnOeb7GKE8V1fVFC
1YJzsIoz4Q1C2wLP81Ri5YhSHuSP7Jy73QEUX7AGidEzQiOfgA+bVB40lF4VfJh/8860MzwynP13
UG/sZUuryipzuTpxEpRHrtFQ6U/DU0WPUhNelMgzt6tptm6XbzpfJUDpE9fIMxF3CHyHo96pKw7S
Mwr1xIjCRNCGDkXgs6M+x81/4NdXJiLGdxHFqb6FnY3xYLe69BjmVGKadqIuNGUs+XPnWUQTMDzi
PTuA2DTY8MBt1zZ7jrw6M6n7na0PNd6DMCFlBOemDCldnWssLKatFy51VEkKN4sMTDq8oSyMsgJ5
pRiraLYId5F+US7uDrrJVv2oZk2uBF9YHKNe1ba8IFXzJs2kmxS9EhPMWoxsrX2KPt98eE5EE6dI
qdBJYVWNTP+ZUGl4tyWYkgFHx0qEuUu3blPCQdqJbpjx923WNPfG9D9r4uiJtqS/PBuZItTx8P2n
QbC+Wb8oWjg8QrN6eoOa2C4ayqW8Te8eW/KKUG4TGMhx27X+HkFR8mrQXLfQYVlLnekSlE36LrCl
POwqgOKWrepUEU7yKyqExkyK7LwY39qZXFmHnRDZITvxjbmFfkiP8r03NvpDrrG/nXyJSABM3mqb
2gRDNPdboIH0EQselPqFLHxNCNuOdqyiFxWikZHhcDaWiR1vBk8XdjEWCruXjRxqNXGDnq91LgGm
tDle05GoqbgH/pY+Ee3LhGX2GrRaGEPmRSL3wZiKJvxm9dnF7eGGf5JzkRkFhQSh3Y2jzglntxvd
uGnn7xKYqK7jqTI2bBlhuHcey1ULL8Nf5v/G5U58Ktw37XykOsF8lHBNK38aoIVLNlRHqlO5MTEc
0ZTCjM+rUg3j0Gink1efRSgDEu2KMdRAhlBpYh7ZIBsGY7Qp505oLiP69nq7IrXlSUIoQbKhDuQl
Nmzz0V1yyWn1bAQgPhFuHETSy8PoZQN24LjZ78oXmrlLlZ4ofId+ccvykC/xbIx+nZwYOcVeERQW
+knZmt93/wW39z28zXsHcBX1P8WOHag2XppY+457dJOLySlCd/dAB7bLR9PM7J+0Y5W6Eek1FzM2
yQbO+FMFvMX+MQfvOVdODCzgIHCtGzl9eXzmXm2morZxc1vOSX1hRP5fFCyj7T9/lI2LLk/R3rtq
aVmEb/QvcRukOWir7Dq8q8lE8AvicQSOxzh1koQLCo+yIAPuuf1gfckH4jtbBQDOkEjScwj5hGMr
tMHAC+Lu5X0VRRCL4tfqiwO63bbS5XPRpTau4UHoZQMUwaCzmRFmSJzPna4OZeMu/y2wlrWxZG2w
EnJgseJVnYQ08eI+cgItlw2SiTGM5TOJu/uhtQpV7qjkpV/2FTrUenADi5ipJ5r+/d7kVD7xrevT
uXMepwwjgR0OlR1e3istIydAk52knI99qJ+OfHdi3+Dm5z9m7FufwL9b98hlcpw4n9vCkSTdBI6g
4K5/TH4YAoSpVGm18GRH5qfTHGUoWZ3utShBVQuXHrqojhs9vOs/3k6jripP8D0Ld4F6tcU32P0t
8CqLeon+4+IRnILtpheEMWZeZyrGx+jp5GPDnQG8WVXBduzehgmSyUCNAmyEtGJctlX8mJroFolu
waesG4o92iuWhqAiEP4kzX4nTD3IdrUYAM690f21XrSlg3tXG4kaZM7CuOsiWbAnumbqhkKtcHxT
mMLD6fS2kEf72R++Db0I+bDH8HtSzLXCXt/gUldXou/9EY8luFbw0pvZJ+rJPSnDEDjFlbwJ5zL9
Awn0s/rEEQfzHOhYyyzHZPNxRF6A1o9c7+ozlESZ39XQllEMI/YDu2bJtkezIjuOv5LW+pHOd84R
Et+bWJdxXYY9ydHbNssx0QZMB9heGbqAyiZUBxVnNqfgvCWsZRHwaGnvS5S0JzEtb+Z7w63s00oF
bFlz4gDs3DbqXUCClQY9SXqepXPreZ5jA5GpZnLvlXzHyjvh/7PViDv0gtWm5cpcjVoO40Ae89/+
UjmAaDtz08tdtNfHjzcD/9qC5yc9eNI8ad1hxWOWmtaSowhUbXFia6RFJxoLqGEsg+bwOpjvjif2
uG/nu2A/+YCZu7WOUvJcq70MuQ/X8x1vVTPVpgiDq+UCedGxZOkww62hzs94jju1olI8u8PSCQR8
/xVhYHRE31NlKHyLf/sTg/SWjEd6DrFKnmYB5NyhEOWloNtntB/+4t9tnd5aEE4TYjZu813YDstk
P+oRjisjcn5R6B5DVxeyjwzuTYyslUeSphj4UOTyTIVMnWE5u2ckHb5o3N0JBY50M/yTUsH7evuI
D6spnF6fVFXreimVAzpGBf37h6D4bCOXZEBbeGRX3htn9MUGAn+ejNvyRnA5saZAHCmLlUHFWynb
OAVG+EfzopJJF/FJ94bEyyQOqpe3or3ZaRWhG63s4GPm6mPsoTi1v5JiwdQN9OGZ+EGVeWKNdwKc
n7CgI5Ki1kuE4rKuufUnbfMF15suwE1DiUZkuJH/GfBLtxc7rQqNZ4Yl4GTfINZVtoYFx4Op2Pl2
5ScpD+zIOUo7r7Ob1vs1ElxUze7HJ2McBZetJcqKcWftw7OE3F4qCDmKKYPbjNoIVm1gUkASM2YY
ldiCFWAGhQIu6aoWB/eIQdoXN1OXzGpuDtxLqkOgDSd1kmeleHTT0H8Nk5G0AYaHwc9ZHPweompy
OpHcv4w/tGjOPTrXxobCOO6WwPYDQBKorDaiuI9Wfv6i5Ek13NmccxQWBkwC8ppEzT8v+L6e4vb4
FSDOZB2stBC6md8MsxvUy2ht6YVFG9MkCk0yogMhQ3OwzDnlqwazK5kRoBSi1eSDQQCWzxWlCgkn
UhqE5nwFxI6D8fA4/9wel1hzG5vbsDrBN57IyXlr0IAmDOCiT3eABMH2zir61fphEAs7TT3SpjWK
mP3xn/3QAMVC+4DhcsgnPi6AwZ5kywg0szbnU+qwhFl64LHlxBGzO/8g1urhYUm1MshjiaFaPorn
6gw/dzDn5uQ78QtYK4Iz4VuDanWxybfjDPcMXPocyrVOuJ9Kemn5zEUhCKpH5It9fsoq04no1dLU
lajn5XZVawQ/F3bK8C3RLAOdEhND78ODhethMZlXUOHoLAP6VMBVw+uVDht0Uxo/2g/iaMhkjkBS
aPWhJ+WpIxYbnplpXsJ7Aa/q6qlSMNcNil8ieUcqC4godiZT474Eq2sUtfZBktdNO2ZWrQ5gGR/4
UaFEBjCEj0Di+qWXJgiws2xNDUEv4OvwgpiIQSf1DlENB2pu4ldka1VnyLqmMjomb+XeO6N6NNn4
rAXMwvNNq8d9eoHjE6I7tt2bzWteYnLtQflKT8cmcaOe06xsyBHira/n2knjk2A9Jsj+rvzDdsN/
u8fsuHvgONsvqPpjjIkTZUMsdrz0P3xfn0JYSlAkJAdoDFKYRdnlInbah38g4rEosYzVSVX1C79v
5VMEZB2m9FDoI+K8WMzZTl+rzYXrmp161MABdVO7f9PXs7rfVVjA9/dfeuNzz5RIbahbxSkGvBvC
s2DclaeqsmfzNHa6S1X952/yCXLm/KCmxN7l0RnObCfI9CJJLM0ZfJR8zZZUqttPH2xSyfgD8Rfr
aXlab25w8eFKhm7lhdbIPEqngDxSrV3Lm5g8Ph69bUsHUjJN09O5BiKTp1AcFquzm8b2mh1M4Kpu
p71wKpMjZgxlL0PI2ZYgmlUUk3AVNcql6uZ0DtW2dltHL0MXeaVeVx2UhVwPgvrDbgbJ+NT4tNYi
DHFIBDaqZr5Keq/k+2QuwAQpXCYuEJUft5m7I79zCca5T25+8wbWDxXorpZxKzbised+YeIqCe9f
rkatzePoZQktj99j/B8nOewrrqhpuWXk5sWwFY58Aamb0CTNfl9G6IViHet4HGbupud0NlkWvR1j
OZdsbtiZLFIn6syBrH4r3pgC+nsWw7/wIIJNv5Pgw3h09cdtbPzbBN9u2kv1VGWPLY7+qSav1ETW
K/Poj7IlwzZyG03V8ZJ/BD1udFebJiCYlbHYE9XP7/6QZ9NeEbdyfLcaneIPG9z+4YYJGw1IWJrj
/6xARhQMzYvm8U1D+xKMBxHfVgFdMWlqcie4Llz7lHcEAfIP1GVli9JEuEPEyanPm0s6GTSifh+J
VADgumYoRzL+Ga4AMJmeLD6F8Dckl3khx0DJ8QnxKq9MchodmXTxA0+UtGiscsW67UegX1vs0d+A
fd5/v2i1prPRjIdYLQnd+9u2gux1SBZjMXnO7PzXUYug1S68vvGpJDSCxDbeShICOzBKiXBN8XBb
j4kPglK1tDNLOPa6gZ6wQByTdGJp9dr4bFNXoTWeYp4IuYSyPkADYJzAnYvpna8LsRxaMbSBfjr2
KF+GhSf0x/OuuaGCGtOJDcT9pZE+oWfce7I2hqF+pIPCCqVJQ1koDj+1HWbFGrie3C8D9ffmmYuA
91IL3C/qtE+dfj2Nwk05CC65FwB553sybaC4neDs/1G8iCerAcsclqZcrpP9Ym/RvPgIkxohx5Xz
YLU4sJrrDO61IX6OwQlX5sPdZ9aB/NL5mK6ICsnNLdJc/5X4/iB0+pAeFnUAfrjjhQ+YJ1wBd6cE
ck46vylpHZI0MWzKlNlVNhvbN9XKVaRh6edl0HfeXpd9rpaNGAskfC5klvMem6ih9QnpbDF5Kq9e
PK/FyWF79kSB0SPqs8xfMHglJ00T9H2fVJcJnlES/EdbYfwEJZlFZYWDdV8tbP+B70GF7qz/QNGA
PJkELYXTm3jyo81conNTaDVeGIHtcXzSkr5Hbq/dr0OGBvqWcgkjXvhqd33tJaf+PA1B5Gtnq7Hp
Vps9Y4e9OvqVB3Jad3DS39OqRpzGeGgWsZH+IS/4Th8tuvzINwEDRDZA09xRr7cUw005pKrEXUcs
V421wJR4IU34a8sMAZCDtWIqxCcjcWNtUoW1bMZp0JzrsVZm5N2bpexwnihovdtS4lkORl1f/2Fg
JCdW8Ll3muyUF/u8dC7sJePo/gn15kPLDAodOe1JHWhc/6FzD+4hzZZc+z0yz0FDFk6gCqRGGXal
fQ06zzo6kJ63jVsUqAGQFB7QXnDZUTQINUU8U/HxEAmk2y7uNcguAigubTmaht3T0UPClB8aDI+7
N1z6Ifih5NGXsxyZro44g3LJDI8jmyxbC9Kw0QomUNkmxD5JJG9sz4gRD7Ry/9o0ZjZVDUalH85b
m06X8ietk+7uGa+tp74Ycta3v48wmnMl1S9VrybzLp0BwmcNMsZ8hnP+JAKzXUBgNSpmyi24I/yF
NPD2a3aP7kE9dUQP3o647cGh9kIEGbU0+ffy77+GrWb9cAWW7EQ3KYfQZ6vME16SL9m8bejOOR31
pSyjMHpGcx/Rqs7i7dMmEn1HH6R5urK8JPXFxQYDjUhZirqqPN9mXgf669xDkAzO1e3p1VVZgY7/
dZF7CMKMW0DKX1+tNvFBDoaUTZILBpWbNmzw3lTSo/9spk2dvdy/w+JxRSQ46j5jHzPx3lXM+7t0
ytvZzQb1Y1tfi01GsKmd+JRge4xwQTCcwZ5s/4otEGRUwfWkUua5BiN5RUsZAP1r2i8mNEaa6+2f
iSlgUc465ml38PWchGX72JugGj8SXtCbCilEVmCt3tMFU3JLjOAGU5Ujm9dbiN9JRVOQmCzK5QOk
gj0R6RnY4YbeDGMkpWzhoMoSLs0C+ELWsCX0Eb8NgeiCwDEZBycKXlMgluu/x6AWCNQgW4wjA0vR
dGNfO/2GFrnPishQsBmmHmEP7PaMsQfqolQWttHF+UAhm5SCgalLOo6n+Xj4VpNCNd1TbL8XJBBD
m544a3U+/ga6G+AEEioaoym16j7CTOsAyfAStrlZR/wfpOEode+rQXrgXKGFsrj1AFYqG9Gfchl3
PScJ2IWEWTcce9SiixewTSHjAc3c2xWXfzTeUtHaObiT00oLkyNAD2zEjO8NTdCHYuup2Q3bi4qs
hscEI4btPgJtjTz9Nn5brejBlkvF/dzDWkmd3k/EgCTkJWnEIwXmBl/ceW61JUq2Ys15sVfW46VS
ReNg8p309w5Tn7Cg1/yW2inZ2ZTalyPoL7ckaP3VmzoQY3dEdS1OFF4N7RlPzugnQ4I0M6aVOY4g
hGAHFgddok+uVLtrVe/DkEZ9mC1sdeiVbLoYSs4D8yEwCzTUj/EUg5hRWDtE4xbU/Otn9X8bEu8U
ZYNlL3K7gzbxTLwHMIBBl9n9jusZMIIvXSaGdl59C3gmhA02Edkm9qeTG6bb5ghfuKR5yG3zpiNu
PXx2Xo+nAGIHbeY49HAs4yQjjCwivDWDeY9Tdo6gxx4pr+1Yo4Sk6rZ3+hDCxVDo0ml3xG/Gicpg
sot0tBN9X5Igysa2vQtMp5gF17v/Jq5QS0cHYc21sinS3zCQowQ7SjYK55b/9ov+YGiPKvOFg9qF
gJhg6g8kG+K42rMzDW3oqF+vclj4bF1eXiMVomwB8irKVI10iWAnhJnhjQykMc2sIAzTZQnbRp6h
7ghT9otg04RFOIrQxhV95z3v2lR+pH0yrHYJpRAxgKNq4mvdfxiF9UE/hlsK55KHua0PtSrVM1p1
77OmpK/KRErjk090UK8h4Qbf5FdBChiyMG5+iIpujsw63LHBCZ7w+CP81CUvndJA94KEQHDJrS1P
/nf/hBqZiPEnVCgVVX3JyPbL9yoyALSFVjZPBQXQfE6XH/oIkHXOAfKckK2nieiiTipcRqk/d7aa
lyC5vx6cN+XyrvhlGYUQN8ZCM59tZtl1s46WXWvu0urQsOubgJtWsch6lJgRp5xC1zTSW0lpFqGJ
eeXBP+NdkRxHBnclsu5v2476tODH/uGngUdQlEKqswxjPSAx5VJLCw5UcIs/3EThXrNkWnTkfiWK
UaHOkjbQ69LsKYuS9jVGxwCS9JK45TJAngFRW4z1NMda8d2T+EEk+l7b1RCls5SaNuz1rdRB3Om7
JZL+ebC8H1trePB+l86TDWsIiTKcD/BiO55DOd5fznr+IZsmgFF8gdrUz7+nkwHOEsQVipsEbzlz
qtVFzq6pWhVpXoz/b4nEXDV9x4PF89yUtiovPcQIPIJxxFZZpIWRDxJLdHZksDKOBLt/UOa8kd4H
4LwTBRrJY25TYl7eTa3fmLwWKa0RjBFxiENXKspGJ28Ms1Bi/tMQ9c2YbBjWMK04ZJocGTL/ZsmS
/jR+dReXbMHdnqa5PRGtM3kLzBGmYQ2yvDCHSeEneQ8UGsfFEhInwv9IhcC30k5Fm7FI/UBRyNFe
AYchxYmeNe8ZOj/vObJq91tg7i9V2xBsLTJF6UYfEH0NwpALFTrL3tJo33v68HEufglzH5GcE0Ip
Ma7DZM+gHVyrzQOxtz6UR2B0T7+iP7NaN4fBJttmlTT30MOg0wuibAi7+RM0xgIzm2lc55sk8EhS
dd9Qmq6iSS5VP9hnt6UcXihb3vyZhlBbmzc9a7b/lLwwLfheEE07BEr552Yex1xVN8qRYZHbLdyR
KHPrSHaalJ21atVJbY6Lw/cS1tmzQvkeKyhVOD+bd3/HWOAXT49tvVDiDvYtsUM8xPFokJ1juN+y
KQpz34b5/J3oh2GBxdxf/CgZrdruKXqRIdNYtYMMig/AVU1Vr1sUuwJw3SGY7aJL9LWORCFR4E/3
ECFnUqW1O5GDZk/mBTomp4GUUiF94Rib6uo0Da1xs8IO7/QkZWE6Ud6BI9qLR+tn/7y1Mwif7drL
7ZIgiItYQFvp/gjo/ZoPOmBsHhjO3h+ILTleKjMvWD2vIi0m5ND2leZVb507FtkTFcbYwAukTUx1
VTfbXGM9bqhEd6wluzntlCJgsRZ7X52rFEjadaK2vqcT+bptW3dERZjScGAYlE+Uv2aRsORwNkk4
9lKktBvRsyhdYRXIheGrGldqm+X86HPL3FvvJ13DEPFlhPbeMVWkV0P4LQknlmFJA2iSUbsX02Vb
9JT8u4EK9u6K7VcXgeK7OaXh5jBd77i9YwlpLlVblWA+FzAD/a5mFr+D8hMFhbnKGgjkFKV+9CcY
7vdcB4BNQ5bm5NHDrAwV7s+h9fR2evgeOpqgT580WIvgq61EQRhhzXppAWE66aVRJ2O0w0Z9rBf8
D/Oz2UQjgRL5FdmSov8nE1iGpkJ2HwOLULxEKgtdTEHTeETqZLAKfEjVXKQi+1v41L7kDHBvu3rG
/h0pzjdqIhXefkGY9mpmR2CEBCeT0Z62EI5U8jMWrYcf5m7FDMZLxtAV9x3E3WWbm47vvOrupTrm
0f/crvs0fyzEHvZCr4WAYbD0EBSbdL689/z3DIbNsZOsecRz+UPOpK3iJhP+BmUOozneU5PmAUjf
uVmLLHifkLZxxVwV36+yFBXcQTOCWydTBa8zPRwIkNDbrzTmZVmq0TD4vHjxOsMM5GhYF7NH1jUG
0UbfyI5RSeIQ6i1FRixx+bjo5MB1sEjex5MNXArJQZezhzwTYS1OVg8QWYS1P/Jpw2fwYG1lBFGr
gGnseEq5JZJrvmZmehhFycsiz+w+BN1Iksny2G/uo+kACX7TQ1ql1qj10+GIB4MD+hCD7CTO9Q+L
kmp4wqI0M+mg6SkkKPL3g/u60hTmKrb8aekiev3kJHQ/gtTSNoQB1Rkj2hOJcOw+heajmHpnNIiC
1NuIu4m6nnhiJA3Hz0BUVjqp7Mg0vgm7g8qykTsNcxPJ0zEtViF+u0pAyMHNeMkucsjV2ijL0wPM
+g2SJ8Az/Po1k4g5rVscHu+ynNug9ohRRUWCDRf9cDV5uneOXtn3XOx9bOtTcGYiqeFPF0OD5cfn
8C9oOG3kE1+lMxoZiZN5XiMwLLuyfH8s0zn+2yGQdE2xR1Bjros2ejJUiyaNMiOmOunFLW7LvX1G
fDe9XwK61V/OxyFSmb3khXo6YRVcBhvPo7Bvj9IHZnveNf1NpEaLytG3mxHh/wj69QhFVE5WZwug
7JPkyWbKqZnA1JiULsVmhF31shq+4yqOSLrRt//e1bLBBag8ksxRJ20GbRSvU30SCufWaCnrTEuV
c16teDxTH51sR/ef1Cr6Fhh8qR50Nu4VUvwhyOD135RhkYy97eShGohwdtWFSccukmsPoNP/tsd6
WK35ny7Hg2xHv/k5027LMKHHCwlRs4/TuhmavARUbHjRPwCzmOvYZ3F8YmEEvt5ObcVPzkuiff/2
vMVIrTtIlC6fXUUuRRrpVHXXlm/d/PEGyorHKLTn94k5RD3QdxJQbrXfyXUg1IdAburLvcCfVK73
PLkGoPym08bKs80gekJ8/ZgI11ADnJS+HH7NEDppviGixkYzOLe58vRwGwY2BPbXCvrtsxEreLZk
pXDFHujAte9NVwsTG3SCLTizA0dvUFKs5QqRR7vjn7VN1zv5sZVDk//P0RwQSf5AmDX1+K9+xY5z
mGzvHO7rfI0mieX6UcnhZ6Cl9dXdTfw6EWNcEw2NBVw7AfEK6g0R6stBHWlp9RHkuFvMUbKZXhg0
vYkSaMwpDd5L25FBEvcbfJpa32H6cAe8nXWeLC1vpZZyOAHEQvmrlG6gVliAC6rgQdP9etWbJGQf
pLkvlfmHJkFO2Kh5XdeVCY4rtaYiDwNcpHoaAWj0n2P7Hf7418d45oLtdiJWtQgflj2HB01o6YFf
6niqOmjNct5ciTaP0U8vPb296G5UIIKhAtMsq5ZN0nKUPn612xI9yoqtazqbpbQGrRNo4THvk+bv
GfD+fDi6FtQcPJxIaY5Q/MLBSc42RcHxNkX7fTwoMqVzL9w6aic1UGHVUPTyaXqTxdO6cEDX/zv+
W67Bj9DGq38mRo59/Glc0oRCRd81Mljke31FO1/+hG59hx+OcK1nXe26O8262g3rJ4LFkWCY3TPs
KciKbqjqTVCZvcVIoRJxEKkeUgow9TBs/ik4oSSpmvnlGxTILwdZLKdYQTz0SwnKcqaX0VPoCysG
V/qXz7SsM+DZ3DNS9qdnzOhgIEFrHhZfQWq2z3NZS1lxMEYEkV5sfA0HRZml4O4vdykteFu0KGwv
Bvo/LthMJx1LuGVVZ9c+Rz3zodAWG+x3rs9aFyIJCdjFxTp0wnfRYMgo+6kxKSYdcJbxYOf5DCPP
mviSLRi3xHOQ5FoQxVW9YK34nNa0gxDWTMb6Ozbce/A9E8+W+azzec64JrlDUMKqIq4CcGwW7XMG
v1PfH23c8ODB4DktRGfllkfwNFtbVmmV6mUoMqfq8lP/ilepFaA+9Pwa1MZRXQLLhV0kcvLl3/gO
OpwZNZo3NWk/Y0OYws7dWPfE5A4OeiqYFkYVCJ5re0gO44VZDQoWmkR0om6x+57q0jQYrptZUAkb
Sw5wY0Xj4OwM/YePTtz6IF6xir5nPEgQylZ7h0ug3bcbyVAKEdnU2nAV4CcD4fOywuq59AOc1TJE
2G9/b+zweyW5LmDU9HklbAb7fdHQS9xVz82eBQf8ndcOA1SS1H6BWYwqDFT0mMGXd1ZrU13JJdWH
geGqmG6p0nzf0fJ8eboqmQxs1IFzynDsYoWfOPjfTFUrNibAGi+cv4Ct4AVVActyzq4xoMLKLLQ+
GcAFW8tbEcWPyh0Dwh3+VHvwmyU8W7vNuQhDhkrN0ksI/a4tGmtMWF5w2BUlBriV0p5MOvZdsFZr
2R9oyERMQ/3x51/H7E/p0/rLK9ZXNxhdAch0UgJha+kna+Y2Ga2eiK9rhJonREZoanSH3xtrw9YI
nC2hxkIYMSw/mQiaS2Oq9EbNva8FRlU4dGTO+FKGPl0QKkt0Wy+Co/1xcwwDB2LApetuooFUYDLa
x4kQn8YLDx+r51rKDm8rljk+vZPggjOPA8dli+385NVh9GQCy990H0sii4XqCa/6d+081FhJTYT5
WbKx0G/ZHqmxc6aGm5iiRnTr14uxauKGsfzN8U7CEF2ud9+RlS87jAzluMP2fgrPy/oV0Pf7E8Il
3QE3HGXxjFtxVN9UQMMRRDI/U9cegkn/js1A6zX6hEPmlsKxONAhCe9DmOFK/mMJNDuVPMVJ9i4p
rbZoyIGiwE4mGtm/EVGLj7f//juZNQFXCqzW89TK4lrMShMND5f9rxEIVQuAFUKxXz1gi4jzJex1
bz7eF/U42T+bAPWBoPehZykHH9LLhRZKAJKxPncVKVX8zPQjFYHZR5sPXnBE5AyVlDTdIilvC9+0
JZ/ZCIXZSTrpuDS/XM7bEs3mqxHpA/Zo+yaxcHzrEijTDMm7s1+vZXzANkDwmV8cH30XTXFBHW/W
fg2ep2emLgwlYJRshk0Ej/X3SoKX/uDMt7sUpc9w6kmk1wG1ldPg60O1tYQ5WcmUC7L5tOaAaF0m
c7G27+kkg4FUM7Kq7Q1+Cx+koDbI7W/pGaUobmfejpEkoPNJ1r+JbPbs5u3ed15lPOHOQ0pOWIlF
FHX50n06NjBPcTp+XHK4ykCFqyn6/8scTwiUTqtfmwL3jlcAX0lc3OskK53oUQkQN17kp53tU1qd
ZrQIqsSd7aHhIRShidY8P91SiCUN6lO3pn7dqK0Hq5/PzViXPOHtqrQn20Q13GH62DKeQ9/k1N8h
LezHRzDdlL+1GgkvaKujZ8HAo2OyOxpcS0EXI5ocvFAyGqKfaYkjcPPxIeHLJpbAYMsGEj6+ouxa
f/Cd0+ekW0cs5XnHtwS/Vp6Cj3RmikcQL44qyfOiaK5r2kpibhT/3Jmk8mpbSDZap4TGLufI8lsF
QG8l8CiZPb7x9z2YTB6Jcj/1J7tTax5PUTIMrO5jjnYL5b8O6mQadF5c7O8jQsA3qKNRemy/kZWw
nZeIfYWtfXOgNB2nVwZ/vUGOwner5DB2PytH59U12yH/8KEoaemHYKAc5TCWIM9TxCOnSwDcfpxN
zbq7NY96MptJIGW6m3lgL3zHV5K87rbzmBJTLmgBGYJJO+ypjffPrDDbY9hvEd5nMi7r7gC1hwtB
pzPnVNFQAENSzUyvVEwag3XkeGVBQBgLwXVLx9Txu9oKqblh80azTJl7MNhjhKUQ2vPiZCBVaEFR
hbykOIXuova9hbAkXN/d3IItIpo1843CtQMrNEpFuo7oXj98+YAEdG/5vmegCQHuztNBon5/HQVH
vHO3fS/QN7Hxp9376jyGF6zxvXn6uboepz03G/pih75dMv+MHHRPalGUyefcQLrukdx9VCJZ+oh7
2EzS6aHQ2zbH5Hhvs0xjv0yKwH2Y8M+wX4hIAJzGOsGbAZVeWSxQwI2gg9Rd6InerGmO/3MUTkdE
5vzvS3NBuokqEyT5Gkne3gaZqfC5kVln0HLj+k6QxQA9Ip6RCJ5XCzPeZZWb4LkQFG4Fe7EHPo8C
rcRc+2QfT5oXuWslGn94S2UMDzn5VKGc1u7wGOjGzR0EGq18216I/jpWNv7Rr5q8Ete+jWOOZjfH
m0X0RJ8Qj6IUUFZTineRADut32c9HMjJWeQzaQCpKNN0+GbfugReMsGHmgqsRvFmGoz+Ts5PHtqv
RRNBF9FBmC1EtLB4EsJdJIBqb+4ml2wWhv/IeRTv9L1Ux4HSuogBBDKgp0KdvfN6kZw8vo+4QSJo
+y/9rcGQpotQsCg+oa4ycjWEjXgkPDw6mzV+NKJ/isFMWrKta1NOk39jGxS6QLQIhAcrq+P2Rj5M
wZOOh7kpEAFM9UsotylvOyLfKsjr0RVgIGJFfX4/ut5nxacz7v+aHSI6W86adhgfXHROX4bi3k6t
X7IO0ZATc2nTaixg7vALvGLQrO+Kc/W08IN106L3JT+wfw1v5ErjxJzWKTeMZC4iclFPV2p41WpA
A0hYd1PQzZdeF1ssziO6wIn0CrXl3DV8KZykzcObXP+qDTUWVUq1KeKdQGx6kBNJ6qErfO8veOGU
VdfgLl9mPOTUZGyfifVnLEJBvomAkFejSqGxU2gzRWAAdPa5orFvCxJf/b/fllcjDg4KITZLLqnh
5DUaTkBUMkqxWgkmxVLPRuQex339eTfvTSIyu/pwTSkRdgs87sS9Qp0fAlFLbeZcQqDXmrpuiz0d
O0JFDdFss0hYaMOQLGr94xuKNSMSDADHQDGTFHNguRV/QhDJJTgPHs22pnHBcfN+XSZr7Uaujg5E
6RXF65FyGcLjawPEgR36Sr1NdUV7UxaWNJcRuId4Yx8aec1P2UnsCmzO2EDM5pmOYWVXIdSfFtf2
1ewMd81tmd3lo8K+7Yp1C2FFzf7DFIN96EKqS9p84jrppsD3qZllAYQs8aArZj6hjv37cVBUkDpP
LErZBg16mFOCE842cbk6Qv9fmHFQlZsbjhNocT3+CK9VDP/+oJ1wG+voLZTKmg2kbqm+GIUvXJpD
CelDSYJxn2G919aQdEyS8eFMdE8m7a7TMBcAzxwQSuggtcBbiQ3ZvV4182lR2BU6w4+W3l9C+Q0F
m9EUyIE4CpN4MZErki4den3q/GhaRN3dSQSyPr//5Fr2EyMUIp6G7rT2hqVieDeCLAbkI7RbueCl
p7UW0VWhuzZWwtEjdUVAjnQqoj7Vd3omXgpbPalIqK+7BHs987bhk1pCg317XXYJDUfKywzDUrAN
EpXDW26CvmHnxNA9pOXNw5bvGYrHgubOyeDwL1m2HsabLRjcTTgCYgqyq81aA9EOnqdrsaoPkbgt
UdFXR3vMRJxv6b63pZap7lhDPkp7qlieTn59Ujbn2sKog9ZNlqbsc2yjxQ7I27CTkET7CUlzVyNM
54yGB49J1VtkNjJQNU+gfV11Ou1DCgsLtVjRWaLTbaESRQnrVHM046HgZ9VMJSTdjg/Y+shV1k7+
9KThn+cnMfiW1PrFXxcEgIqCd2cEporv0vSzTkl06C67qdK2i81HoLZqFnWKfZaR3awOaXef33x1
weF8zT047a1pQOu5ElQFiSHw/kQRQlm36RbAw9EJek876+JjgLoE5r6IHPtGD21YMIUu2xfSlw8L
a1vKxyd+D2iav4yprTjnNS1Lh0DSVH4lov9MMK9/uPqmlD1EdRXCqxrAty+ZRq9yuJwPhbKXnLSn
aGusEoOPPTYkmH+a3zWZqG5SHAzz3Vov0JRroTj3txOY5q8rbtdk0yHHJxUa94QR/QWjDCS1yLkL
ZM4lQt/3Kh3efWyayqOQji1M+eeSVj1BTtGoP1pC6osMxtiVdpwSdb8htatI5+Jzm36b/Gtf3wh1
S95Dz3kIGWhjlNpilQmaKLw/WIm7fia+sDnAHnpY/QPShsNu9pH8FpWm6C6Ko6UN6iucTSxFiJak
0eNJb77Rz0JVN+epZ62W8mRvNf1qRMqSsy82qnHjqgw6j26KbK6ZlfxtpZForDfJNtOpWyb2a9aw
mR9Z89j2t+xIYNY4PqBhuBDEGtghq14XYF6Fsl9qmwWWJczloxGqtrkasrJQ8n5oq5haIPbcVbhF
9q+RdusvKnFZoeCunS+eBGQjYsA0FobJ5Y4Rb32GxPuguhSJMeHohrDs1GTicV9oRgnP1KvgKYPV
tgb9ZKyw4lHvHTn7zZoCaTOYWJrjnZGZOO6YCa9OzurDpICk9O91w2JD7/xck4VUGYfRsdFdYDlK
DcFr+cPxIT3TvaZIKcFZN6bivnN2SxLTHtP89ZLwYZSPi2Z57jhq3OUEnEeWJ1cbm4ve/2KUCjeI
wS2QCGBa7y2Hd6Xfb+trBlqMDn8CkwlLm4SgrLUUoGjr0GTQXAnhuLcsk562OhAtTX5RmUUaltdK
YP1fXQfYqd1M6r/gKLH032WIuPMnag2MeIwqVH9MZOp/KIIem90qxzb0c12fPY4jQ+3nwev0IY6q
Tx6JlAPGmuAqOFPqtSljgSnE+4WoJR8X4OY2aTMg+H/2dlQTPip1+QYFLvtLaEKJ84G+npStGJdX
8+hm0NJgVRdXbvXueeNmv0d/J+OddTFT7Bk0HkikmT6AVjWg+r9BmXmzy4BaRMJxew4m4uZtGgoT
2hCvMd0rnTwFt1CFhY7bKcr4Y05m7hyb2hraVl7C3pUbzGflXPQ5fK2r5RIY55W8WBi4dWZPE1jb
Uy/vFrkkmpveQQW00/kBIycephF1CT+P8FAhsvo/Gr/6VhbUzqKnBQ2I6Z5c4t3bXYZonhUb2CMn
RtUSIt8Z/xQpYjjCZ9E1kZmm/01AokebbOdtYtQZj8IAp7LWceYMjGGxTllowcSkEbfx5cARou4N
5kFbInqkTlVPyLzOlHJ/jvTDbxGAHZGrrnkcgagO2pDKK9caVlXE10b0GVlMwbnWOqdnGiozkqFr
WvYYnBiDGcGTJRFfeTzDD2DuKkgxXL53CtbRxWB8iKaQDJoASGZ2X3hZkgr8VdITpJeXcISwm921
lcMZKB0txw5lM8hDcigUlwkZ/1v5qVLaTuqNhonP6cc2Y9+dUeQ5icglCriOOxYcO6/Ay6bw9O3h
y3afbTQQgE8X3dE7Uj1F5Pgzr7klQkyMISwOVQD5/wAwKmP6cbAIRWkiMk+6SG12T0p3/VyScqhF
fIeqiw2oOB58xdkdQ3gnlvotQ0XYvzhGJlXyK4saF//8ycxF1SIZ8q3Q3MT3eGwuxsYp/m5WY8Xi
zZHEdIRKtrev1NP8VtaDV8f4Bk5ekF4pE6bpct3FFkWntFuz25cmrnPkI5gx6YQzTXbsN/mHX6wx
B9BKNU3Ki+Ihya9DOPNb2S5UBPku/OLJnZ33o020LGjABFbOph7SaZFZlOXGgJkI7QbSFhkQYnIj
mOuk5Pi/zEd9gGRL/RRHcJidvp7JMEcalJsHSEDSfnuVuhLQlw5qPGXDk4iGNVUlamitX0ZSdU0h
Pkkm1Zj8phJS8d/X778JCVb3BqXPnhgudS9Pb6PqDgSE/xL4S+L3w21gvzEqXI4MWiuPGEbAtmk/
LGV1UBB6ttaX+gCrXyCAgnTzJhPtuhqoCIbUc2pUJDJqZY1NeuFhbQL7uZM1ctUjx38GJpNXEv1c
u3M50mQD3/BCBeoVF2DksPqmsWUsXWZJTZDa01S9uwL6MNCUCgEANySVqLd5Oa/jtuFagLUZH0Qt
p5+kXhS22VZ5xATd2eEu1/KRMU6yTcIX7N6iyJ+D1O13BiR1AEHUqshPdw5tv1OIPI5buOv0ln/U
YAareksj92gvMvlzCG6NA4RmQUv+qX6IikGsnY6qzM0MK9vXqqyPK8Qs9qzRb3d2wHpkrz+7hP/1
B4U4Ymw3is0SW3vSboRApPH8LfrTVMIaVObUCY0GCxpotWoUpQC2vTZmPFt3YfaYTRjoBX/eFEs8
NklqP7jUNIkxj1Md2heTAMqUhjEMgPuGVHfH+jjTgNFkWeNIWlHy/XNknxom791OlrVcNTcDIM6w
JYIljJaOnJbblpRh84f1HArr1ses6RU48VCW/LlsY+QcJFbuiO7X9NRVsDPaWjXqVBnlp7sonaSS
C04sXxEKhJViojSNU80M/9WPugM823w7dXpeJP3v9rUgSMV5GXoKNfMS2gpMk9rgjZl4SExFNQte
IbO7vgZhJ/LG0fzaIQKIzdnjpn7Snl+zSVVYtIV6+dppKx3oW0ELvL6lacX+rPPjOTFv98xO6UM6
GFd53RljsaVnujPXE6IFSyTSqValK7jRZ8E8Mq6hI8UOZBeEQ/uKgT1+Fw/288VHvRh2t2E2VIrW
ZEKTeocom8c0L7PWR1yp5zp205OT2PB+ctHKNFaFd9jAlimoOkxSsz/LYcTrIh9s3iEkPEccvta3
UGFXoJK1kObnrzkG7bXW9RK4qVtEMyDMGFVBLCgC/Ktn5hfOUkpCNZpQqhYQYKUf1vF0elnMaQuK
Q3w4C1A/A0txiKtQ+5gqpiEDchzE2Q7mKWgRkpsrMnHTp8QxHan1Gt05DefPvV6X8NgwDR9Y+vHG
XkJRPqXT2J8i85Qe5S23NB10I7DUc8AbowTwcNEejRc5ukHBw3aGQNB8YT22UtXzZGJB1l3yiU0G
Ihxo6wxqewED+UlWpZ0xDS8nXloVMsXTMl8Iyzd8zrUS20F85qPkusNUxjwHcHA5iRqgFMyGWe6N
jANTPvDPEdAygTba0p7b4oJG8UN5XtCH+Upv/4liNgM4RoJSABLrvnYSQVwB1TE/PpSTrnx1UkzE
LNC5S6wyhuU3uvWJf2Jb5ck1giaJVRXzex5Y5+0uhTuF4DIkaIfZkd887rMqSAVj10A8juGs+8kg
YdWCjqily+Kx8/m+M1mAPQT4nkiBAKyA2XTfmIDYixHU3QzXfNq5x1hGzbZ/BBVRMkW+t9wJqamw
VW3zilXx1h9LLqdg4LQjsD6wTKo2BaMMop3jF5OeazkOmGL6AKj/ZjSI2yfOTkmkvLy7Hwq5gwPi
uHS8LuQ2UUMbFSGkGMaDzgCesNOyisCrlchy3qoF6CPeuqCCdFOVnY2gri4KeF5Os/Hw7aBPQVca
zFg15BRnBi/+6FHPbdxZ3KM97S5BYU/FLBIRbO/8PRfm9tPwtsfWRel3Mnw6SjtXph1wVjmaHXMf
X2l+8xqZtzVx+RJBzkqRQwTf+BSxki0zeZJB1ia01XhrSpREHpGkKdcKmz02focmallA2OTxZ+W3
rgpMjNlRmKmrEWFl/UCGxtE2wvYYpb9uBFQCsSCC6bu1AcO4XVwrRtiSkRrS/hnDpHEb8hzhXpI4
whqqgSo7lbLGvKXJH3gMOijTZwLlCphQrtHKIU62NZcmWu58/KgGDJowHsq/igbJtRmqmvpzf4KF
BskKYK1eYe6vLhjIZY/qpFyZf1EfL3CY84w41JGpYF2wg/iYMKd7fGXCHBCbtoN9LLPHjLhbRsml
uwWiqkU2AM5su44FQPzpi64FvSsvNtthVN1aD6i4XYQGOzZ5SC59WBaiXQvPbXGoOEqLdZ5VW8LD
e/bZH7jzE9HpFZu6Sd/d9AH5Y+kw9+aZl1raF+wCXFlZxmk9LPxAs7d1HtqkIfWGT2Ulh5cP2G6j
YM/qfl5JXzaYK6DJUwN7cWK+b59V3bMit78QqJ4kwp9eqVDwlP7TQV1CwsVp9NEduBeox0EaAQkK
PTWxEEbOGuktctEB7kNkyMrYgWS4jHBuvaPKNDtOThkNCB9S0/mcXvdoW8IvPCv2vi55hrllH3yJ
cKKzRmwFh8/gdB35mKKKAEsK9yr/7SqD1oLff0kKc/LKGVdkZWtXM6X+MbD8Auro+tg1JcytJYNs
RTy+KXscp7rkdsY+EUWMk5La7uAej9elpmS7jaRQmrPjAc58DTQkbdyNSiCwfJIvjtpqGdMpXMlt
MW182IEOJvq71E41FWkr8jpESE3DGpp2jtlmp1jhXu4oiHkbOekyxEO9PIdKc8+MvvOxnEF5JLDX
NYfDBLzjyAKrgig8gVHq0Sl6Zigy2cvTY7g76gSDyExElvKkFZFsgaaNVGzcaFADsLF7qT/eDy5G
0OefWXA3iFPTWpIOY5rbbefPiOXmQSDYaQ322JRmrhwvRmT1xVsVL7zbTIFQSFa5A8mjRSj1ul1Q
ByG0M/lEerYa8SsdIb9jRdgFG7D+MP3Er/2sEkOzmpSGTO7dg4kW9r3l1vM3TWJRuTAIUCAxomzI
RcAceq2FEtwhmcyA79IBbj2YQR0LZPTvSOacMMCfedJue9k4oRFuHow3OIwukK9p525l1PGH3Vq1
RUR1dxyQWtDQk700ZITBNh1FCbP00xvfFQxYTUIkCi4Ki1lJQUtgYD+xl2BDm3pJakg5UQdH1L9O
oMg1Jrj77S9S9qt4e746mhktxyhwRuKkshgvmSmc6CfTs7xVdtFDjt0KJxODJey5n/DsRmM59thF
Guv/SSZztaRXRI2BYxfKh2PtdhTG0J37PHVR1QpaiCpcXjDwpRhEXfNRwnCIrB9m/F4bvOCn+oqS
9zzKe5HqUtAqkBVph623EwvmGVQICMvxu0pnPvPhC8lFQOXQvr0a+eAVO/OlxcGMAWJbsOVXJxha
i6eSgU18gEevtAY6SDccMyPMYOfOuDkoq4Dbr1MQt5Lu35tmhRzOGy1zCrZigZTW8YFUy/Vk85tc
UqKa/evKkYQcaaV+R82xuYLeIzqfcO+wAajhgPX4xXETeesO/zvHznIvI+S6C3HZ37Rqu3J96tPK
13kybFYLYeLUDN9Ng6gkjYELBPoPtGQZ3DaO99I/9dtbQkAT96JfmAfIICMCYmoquTgec+vTpVTH
zxY1u8wZAvpgNfUOHbrQmjFA0e0zFbLc33Kuw6AC158zEuVNBT4TirV3aGWTCz/5KLS+aPRlDGo7
lj4Yw4ZcSrxZ/yv2ut++frPTrP6GGhfby7nlyRoo5GYD0pmC4rLVrId+JZt4rlILcBezJrFTvyts
kn706C0wFWFJWxWeBivKeHIcb7FerawBLZneX8z5Lufi58Wej4TrHLxDV+plFHgguVAoP6JXsZic
nzKxinN9d+MuprMTKOKMrh4fuJSRTp2H2vRnu/A4DVh1VufkYNxQ+6arvKBliSCJQeLr3O2oKEnB
REZvrL0NW+76ur4phJWGsvsMcAtrNBA8+m5pdsJkEVMtwf++gfXVTBwaFMXUoFVlBH/ROqX7RxFZ
frMvsrgo2lIL7Y0aOUSISOB8LJxNblyvbuzpE4jpDcnIrB/u6uPhEun2/VjZPHKJteCLshdOI6J2
Zk4HKpTPPSOkD0izXGxx35l2IJ0z37qm7t60NNfv3MRbutx2b26U5e2j4EVnSk8pV1sCRBy8d1dl
KOpax3Ic8Rf5pE/uXFrowc0iGbZ/Cs0vVtAN5+PeAV9a9Ywu6ZN47aHFoZwZYTErc5EAaf/NLYlo
wWHiREWjr42tnPGSjGChSNTTfsAHGxgm9gUY07W6TdlpavKhotGAHi4OviY5jyVjVL5q1HSq5u0g
cF2lYDIsZljSYXpxN0H8PfV7GKqyaFxwGbuNpmUy//QERaYUmEHj7MP8vh8aa7Mfh5R0urJPxCRd
eVD5bg8lMbocSKDYbIU0yN9RYH4DaBBEtTmnfToEGUMi4NMzVVN8NMt5+SsETsULDDcHFzDoWKuV
/pkm9ssqmLbdRmWyX2zn55qmOYAnE6wMOQ8jZyy7dD1oFRezq2LNYreotj/yUvdtodWZ/1t+/kG9
mUv98Yo1WGfdq68FAKDd7+53E/SguL1ipH870owzd1N7TzZAw/xQXPAwHKS6qs4WWx8A7nHjkfbU
VnU8FS2umgd33ctz+fLrV2ts4wzD3DE5WuaQx3VBts1Rhv+ZApRy5D/Fgf60vEUrUDxsjGAqED/n
iOHddeZ/5liQhWqd+3sLHGevPrYjEL0hNfeBaFgBJ5+4scVWFCIT1r7ZDRs3ojQMtnISdWMrXOAM
UOPbozLbyHBQ9CS00HnMpaaaI/96Rpf2HSVa7/UbBxHkJ2ozB13LzuMY3ZC8T/QFpLlQoDvKNtFK
KyW2JWdrN7/AiCqzuXtMUUShZ2LEbw0lvEQC/w2m67jYDHJ5v/OM8hTKs7X4Mqn9fty0xyWdGZ6X
Jqrg0JIBwhtjhXRa7208PtSBGskR6Naq2A8LRFOojMs4Jtd+org3FVfeIEeY6h8YAvz98CGsTQqb
GOPLqzV9f7xIN6FaxYJc2CmbyNVw0nrL4bnyn5lGkdXqqBuSV/IIWXm6c4kdJHRBN6lfmFdhcyx0
mRYwplFb7N9Xqi91hPPBNIeN0LjLcNSbgg9uhJinUVOSjT9UbQY8g71SZzxbZx6QV7ZK7tJH4Iq9
NL6E+91kKpOhiBCyHU7FcfPaEpeku6cuJ3twKO7p9u/ye6c21PIEmI6wpbil24rNeuq0C+qrI7P1
NelAVGEvCtguJ+tvohh+huf7a+YflID0AsRnjDYTdFi6hQCKN4FeZS16OzlCaunngltD82W7uQ/V
MsEjizS1Emmpp4IKT12w0MnPXJeN2suFB4Os+sojASiFLD1YW+PgilRHZi39ghwVyVjm/5Uijoje
iL4W0alpC/eo9pjfT39JbWTi6Ca1mUENmzH3UDRWQVMizU5i6HSwOXPnnBoTHo1kVYSAdJ0hfmZ1
V94SftdD86AddN5uzVo8zmoRNOEaMhnq4nuXDCPn4ROQRJsP4kMEaa2dzT8ioNmpptYqCoLE5IOP
tYUSzDjlGqJEkGYZ0+2gEDpdxKcPlafmjzy2Sp6jDaJFOXL4U6yU4oIFyQnbbx4fHi6HuCQXDMBa
w1tLc7vYokoMrlHinarCNY1/rNs4qhvh664ToMIwnGBr6+MOjKWwwym5QXEZubu6AJLWyiBzRQk6
/itgN0PbwRx18jN/w134u0Abe2pqxGd+twWwqvXghUC3fqhGgxyTMLQbFIq5x2PW1XOI+k2dTbpc
hUteBGjFjfBZCqjkF5mQwUTdo8KQqOQIn4jz7HjHs4F89u272vUJMCvzbnwqMo9F/2it2PKQ7zzG
sTbbeHB1UEkcmgTgQYcpPeJLQhB8yB55gCzRripTb/xGr6f9yX30ou5scKPVc1Lv57rU/wE7bII4
11BE4Tozh6cyDM1caVnon72MbBi4EqoHLqPFbVtRtibLcZA1iuDDOE0WbKMV6cJ7mRsGsVJv7zfi
gWfKYsOyonuT8L2dtjN/4NA8ZoyipNkL5Te//OTj04CM6ASIFG9E+qIGlIIDWFk2DGtAW4Tjb0UP
cIPZWwb2EaagHIbKT/yhDS8PqtTh+zKlSvExCL8VeRkkB2Mg8F6pFKYPInhZ3DXcUmP1aib5CrN7
Yg46YCrkKFuGETS/JjUHVUx57/9QxYEljgLADqV3S8cCZZTlBsrSLij5QYiSv8UNM4WjjIkWNe07
c0M3aAQ4lR1b6EigDwBKRUCZU/39oenD1z+dknk4M4tlOIqDON144/7JqRpySYP6GO1q/vZq1PSc
iltME+JlT6itLb647IyTFo4nKldMWGh8mloWpk4QjnLGlpY9NrYUPn/lPEMgJP2mby/db+aTtDrH
shuHIXjqwxxqgBYYajz7Njm9KLV0v21L9TWlffCTrU5fL0Pz7Q6BxDH2o/wxbQ1FgaWNV2ZM2P2W
HHHZaQis59I7TB8jPzuEj/2Nx5aarZGWeDa2sg2EvB9a4bVGh/3GRv8cyUPDidkXsFtKC6/TQFRH
80Q7/CUwGS4AYOrknxJHfqKXS6TTE68jMwKeyT1ldgvedT3nQNac7zaGb2yU91MnVuwTwHmKoGrb
zYgkD41rpyBXq7cGkBnUPplBEL46CdZl3pPUO6JeFnt7Oae17n4/8IJbbQpaSG3D3Bvm/rv2wQEq
T25kkWtGNkiirbynyZUMbqjzyeZQoKZ0+Ma10Hr20XFLRHQ1wM3iKW292ZsrSx7Q/MRoDhnr8tNN
90JJnHn2x/fLiuBS81bMpm/LsChNMdv6zqcapTiT5dW4eG/aoKXsFlWS/LdI/ZkUZ5wTFY1QIsXZ
jSYjejkV50Az0WUJvuF2Jbgk2dgdvTLY9S/nEM0JHTOmZ6znjZCDdQBej4oXAwbgC0GwwOdqqiNF
C8iA8qCYNAeKhOxABKXjhvHamWFGd+slDRAN68/1RdcqEn/f+nkloq+GObtfU6UQ47/qkvX+Byzy
KbuIBaF9REY9cWwYSuGfg2deF/HMrQMeAYjl3r/suP/LfrdBaM7S1jmju1yXbfgJ5qKmczuoXbnM
g8W6e1B4clDECcBiIdMTP3E10w8vtiGoQkdnWGJatlVVDOtb/iJfiYMQ6zGkJFCQTpmmP+E8QwDp
dJrMNuVfvV9rrhPRWfi2RW6kI2b7qL7qtFk6XKqO1wkX9UDwzjSkdfVN9/uwUgXa0rG8Yy+YaORF
Z47O2kRFzIlRBXBwBixak6delp1Ixx2TrynN18IpQyDmXgkALAKAobxM5pERQrGabT/CHdZRAWlJ
5iNH28CJgV/+hj7GGSZAHN6N+EOFRuNnVfa+d1dTptUKiueRa/OjUXY341Bq4Sd1T0xMgd5ykaNf
brkHGfXTGoQ+y7/3M7vUmwigiumgAqTy63d1oyz8UiiIx6XvLyaiiA2LwlVpa9sdKRgHi+IBEaum
kXGLA+SRQAFSPVJ2G6v/x6EP6uYkXZwUau0NorGYWWiCXN42Ttw5yufpvA3AkVuspPVn5Vn/aP12
S4XMlzFucIN2bIkbPjHg8xcXAFo+dh6htzrJJA4salWwQJYOy7OqQ+RWI6tEg1O5Y/88EOLWByiX
Ph9GS2qDa++qAhufoLQR2zpda9PRMwV9Z1kSSdA+5fEQS3QXpSZfk+shQbMkbZmW8jPOqmv2HCaO
o8mBCnKUihwod/KojuvTihc3Jm/CjIUto1Nu1rPIHllGXn2pkYmYL72nmRsnJrVkKdE3616MNbDd
+ZBR5vvfloPp1Qb+1sUabwxULYdWQ7BJb5qtFUYF5lIG6KX+6oM7QAGK9vDhkeCVjwuKb7exeS4H
e2iKtF5NtEwSCpV5GizNeiM4Oesyi0ny9o9fbVarvdqa3+Qyx2OW4ipMjIHnSZIYq+gGnB43huhP
bR78O187biyDc1tC5bbL57v9NeW9QeMEF5mp1hfolV2VQ+JcT4uowAvbnRpWZ4FsAN9ng3y9UVEz
dnQrk9RCATfmmNvD7NMnMfEBMlSk58oed/pszAQxXBxpkzTnSnHfcM4Lkb7RzwbTkHpN+7S/oPOx
8XQmf7KDFWaICLa+8foALX2+n4MUf1Wtu6vqCaDhuRL66sfPkF2FhNXVV2jSv7qmRkRL82kHm2gR
6V6usGXxlHz3kDWgIP38A/oTEzRpBDTQR2enOcU4a7zXYJy04TiSvTmIBSB6/H3q7ciO0MOBJkXe
0MY+2aGSgVjP7bVLUkRVAzfsLZFjI/UKSW6uSQdyusrd0mShbyiPPGUswU6M7b+PAeUyCUdopKSH
dueV80u8tan7cfWauMtgadjKZ1yvPH6+oTIiECVUvu1Nn8hqwihfPmFUiXuBHZrgFBLOBJhpwl84
3o0wPomCVJXFLnZmSWzO1O403xQqU7I2E1YYlLQqSHJum9TZ0lwfIzqp5FLulPOCCDAd/OWqOxR+
2XMpTWh2P7U3ZDiazAOHiD+6j5LoAOPA9D184oqlJvF3TtR2nWaGXggcbItmTpHi+bpzdlhNrc8Z
ILoqW2o+UM99K6SSY+TLJR8a3siQ6QhvWx30s+2OOARlgEWZPbVMp+lmuMfzS68tv62/57GRKoHe
ACne/nZ0hmCFvxC2UXaAV/VVfICMs+jT9qu3+8yRcFDaqC7iA4XqMhzxjQ/MUyGn5XiThEfqFfhQ
z4Dr7/bIZmm5o6fkajLyU3bG/4D5UsToMPHA2Djm25F9sm0wAkl6frIPICaCn6TdAX689+sU3FYZ
l4Lpy86PsjL/7ow4Zb/uB0NssfqQEJjiZ5gGNvU8qt3RdHKke36cr9H4r6RkXAML8D1XA5s1TT8j
5BxysWNhdadYWQM7oju0+4pEVMoZnzBilY7oleXPTMD2qOuIPVD5tzv316ZRIOx8bVGmj4jbKQ9g
A065bMNQj4CJSCr2mV8Zb/NoFtKoblnuZOkimN3b48PADabOg15pY4wusi5tn2g8SITAcKi+mN2s
KHoB4hKamiKBY9WmxJacP3vqRM60/uUpEpMcs2QmP3mKzO76LTHcLmIXkNX2u4y6DAgC+EVmt5ce
aoWiP/BTqdi72Bj1pUhdMw2issR04qs5NnxO6h1zRuNruWc9on9abBRc/fDjH6a83661omssIIFG
jF3FjVD3D3HODD1VVWgciLUpVJlfKVLhbWJehXmZyLw6IeWJLn9XxitUTeF7ZucQGxtZbgnz5KnS
fGcUWUH6PlbJ2iRyENNWDd9ynhQNPQcCdaFA7sIbVN7I2gUkpy5rVGVjrJiuibVdsRwnchxaW+OQ
wt4M/4fDcAlzBZ6b8HyEHKfH+0h++fUwF0WNiuMO8w+NgUTozGtrx587Zbsw6wLQ3O++xD+KwCit
6/g8iFZ5uPMQ/NRCGN5VJE+sQyEQQMxyGRzIumJg87O0V7+yJMqH7T/L4yUokRBzYjq0cc5GmFCn
++8qVo0qjXTWYO9/WL/6l56F4RgE4cdGw/d9y8u0qj66QNS6yUKNaXsTWMLI7HqO6uzQhWNLKa3b
nbPslVltcX7oaHrhjs2I5vZ7OjCznhxizagffIOBZVcBZrAZZcHaIla8hw2M2bzgD5eFdTT7YXnC
V3AdTqeyWGfeyY3DmO4j72zOIQxnwyjADwMwp86k+dySDsU8BuFcmzP9LC7Mb4+NQb0Kd8tQn6hv
zfznw7bT9yWB1hInSKNLlt4TstAdCDdhNkjZT7hhC/6Y1DGcwWbEXwIQNE36S6pCH04IxCTEBcNZ
w4ehv9Ym7XjLcyqSsD2i1h1wTl7/s2zpFEL/w6lcwyoqofTisC68PPS/OcWoLcd/n/AvZkfvc4Ht
V/b1ZAwzd5v2FI9/MXvlxh6Mo/ds/NUoFVqUqpwxV5mJrknzDzr4I8Irvv2fkNgxic0/mnEZ7lyr
RZPJpAT0CSUxwCBSjwV3vVVgFUWHKcArJeKxBG/fmB3zR9FA3yJso/NRAva5+T+JjeXnsaVrI5sN
NW0Dt6L4vOqZrSRuRUTxq0dy75KkAi2PpH0RYMTteuwwum1IfUQD7W/lnLrzT38k4iZI771+dwUr
iIEKHm8yHyL6gcwUudEbO3yV2li9yIKO2O5FpzL/MoPaydAwtI0TAQCM9PmsgJ55cp/yYBeforCF
XOMwWSjs7nD/jD19+IV1vTGH84jfArktDs7yjqoWRJKhMQ0840RMbIQn32jHfLE+pAhHxwuI855E
HkXx7Xo3m4xGwOcAlB0ZTEE/r2OnabGcOYtYkHKxkklt6jTKGgAuhD2we7UeJ0d1vsUoxLUZE6Gi
uYcvOcFN2H5SK62730OiUX9wCqSrbRoolo3tVUfFh1UZu+4ok6Y8f7NXi/DLe49qHW3AKcBqozKT
LOyJ39KV0gScI13w8Z8fhO5gfuSHJ/oyTfxFqXmwxtJDtW5r6XhsrxGnzmWYYZXSljjEAMoTrSfi
nzHisbr6hW48Y/pE0cYsdh+uWW0KDpQigZ5oDE6sHF156FyYiKylvsJX+gwgFsjLyYagvb9taNne
yA7SLo2CJT1lSkFF1tQCFCZDdcCUCAcpg8AZaQeEGWccxvrsPiR+gwKLbSQZTsa3Cs+7fsMXRyvk
3LCYgM8JVJGFk+h25wnbEHA3YjgStH9QB1vckJ3Fd+AZyk9RYppp2SL/qEFoPIXk0wk1dBlE/8UZ
SQfoLriyugsIwctN3r5+lNDsqWUyQ6ZSwFUaWZSWtoFqSWTvnemLVgCAOjnA8IaGZ81Da6JOAIOg
MXvaumbdoaAhysWkAzqoYA0k0AigkBgeUN5hYRxLyMtrAkdlE+s7abUgT+XxE5bJz/j9fosY2Uk0
9pziX0RUa+iicUaEuz28SNagdIBgti0xzF59ZodwpmfnA1C7mLL2Ie3dtqz2tR88P/hIIt3wXXeK
uv6jp3YySgMGNpUAwVCqQRKD14eFX34vf625rX/VEGTufSgjnasucsu/rN7Qsi6B3WPGo8a0EcWM
VJ2mLjdU+jf8jWp/qAyvc6/kKwBJAay3kZoDGtb0JuugzBy9R4tSzdbf9sAkhgfWmFPWGE4Dz3Az
Q8zwirtWLmgeqlgGW6Dv9xkpv5G6jx3/3dHgVgukmTAqu572bKqbzUCEKR4LOeg56HHjyCKQ4Srj
e+x2wTBFE3bpC/dqH+jFD//UnZyEhXVf6HpIA1XLpLbu4sw7xau8v5YEl9XgMUPZKkcPsSlRxQd6
VBKk8pQYbWsaV88EC2XByG9fOlGq1Vff9GO8NnsnCgVxzab1wYyI+lAFJx8bHLQq1RM4OUQfpkIN
L5RWWalkHY1Yuc6YGjpiuLsLEG9mWefjCLrXSWTguTBgA2mejyD9M1xczP+A3O4/l8styZUh3Sug
2dHQxIIBvWbCJ9Aa4g3I0skCzvofVIrgK2zQ+Vl/J/K59FcA4tteluKORooBUmPx76XeALF3vnsd
eITfnE/C3n+Ir3YB24dwjryJd9pwYWcos6jb87RRwhSrHkxrM5PSbo0k9F1Gg+p2TDxF8efmzcMo
RWUwTyRxQtsuVAuVeC2tOD9PVRg/GqVfN/ARHfVs13aFDRPRLh6mdyTDG4XVfLAX1exo3oO4s12r
5hZDG14gPVLHoZTXWg72eO7Cll8eD4qckwNoaeagIbW+9o/S1QcLK8zzTTZynRz4mdcSOS4ySbRv
QOx6Q8lJ+nvMO2YSPTRWYOdjedNYiZwey+A/xPFAARHphOaO5BVEi3+m+Sy5kubkIwnBVYu4nYp2
bs5fQyDsD6zgM9IrXqQUyoBP5/8MFcbYa/iHW1admRNNhQ6xXOh81/aNXkDkpnTRBMRrDPynMbdx
hLPWHipg+5Ee9DGhropoIvbx9TPOX7Jn5BC02diYpBf8rc8+Izb8EBAfYkIY+LxIxfkIWn6mAojx
8n7tW2SQR0VsuFqd8m1TNq6OVawz1SzSbJpoW6WQTIkZS73j9e19SgSr+HK3slguDSMYWbmkGSBf
O9BsHDqElKM8WQHBI98iwebAL0QHJ72BmcBJVQCwAufTekXwHglVmUO9YkDSGF7QYffJFralQW/y
LXuLmRIxBxYhWLaZ+HpcIpaz94/4qeXWIE+gC/q6qZ1eHbuY0IKy8btyhIwCdceIQZq6hnKMfNNY
m5STz+Zslq9JxOTpk51wp50OjHny1SA9It7pxN6SQYg31wYdPugl3qfU+YaXvsHBR9FEoyi57DjE
dhmTkN56/KPaXYxphtGiBWk8sriCrqVqK9f97Xix71SLMZ00HfnY4F2KgRhPPVrxvhAac8MX0Gin
BHdRFy1Ecmztko/vQvJkq5Z2nktQn/r/Xkw2ztqk32Qb9hZOYvK5ybrvsvEaxyy5Snf0b/lpmOel
6lZR84/SY7lssC511rNu5EMiZC+7neNrZ6uFgfDc9IKBNiGKaqZxvAoOFMsZTH6NQ/YlJc+Fbb1D
ofSHto/kb9dGFuT2x4EZAoePAwnHSK9F2HC3ZD7JYZQi6O6eSvNOO2rE6sm87W/ghCIJEtRI8CSO
Iqn+Gbn4lNQEoLgn/Q25eaKhwoWeeWNEFgz5stybd+hkhW0hI+FhQRTLRZWqKnouMXqZBN0LgYXg
76aUkQGgD7dvgyl6U8IkRHsxHntP3PjgRxWsXABKfIRyIu9S8r3oLqmqmLi6VGnXeVQwnO+TFy9r
b1bbikXAzyKsSkN0ENfbUloMAwr3rEefeXib9LhugKD/qRCCDcXkARLyCLTMx+50m9Xncu9UsC2t
7rUD1wdaO+g2IylZ8CIlP4Cc99uoNDc/Mlib+QQ4vMvp0H4/teqjswCHMecKyAbXw98zzth88Umg
iX4eeg4Di9rEefSmKdysMCNiux0suMKyIjZzC8G9DGegFMw9e9RsdVKzMu0+u+xhCajwte4kcGvw
9pfdR62LooMuS0wbvyu48QtGNpuYURmQMus15jFvvyFd/uq88TU4T6/8sc16HnV5RMwhThC94jfL
2M19QQJIxh9BMArfrACK0dS8+l5hBimLstR4MGv32weXD645HJJfA6tixnloQszfhpD+FaYpU6OI
zpr1yXRQ4sHujfCMmTtDC3hXzfmXmmHzE3SYpuVCJ5YcyqRujNOnIxtpEFgHtHBQc++VbaTiUIG5
OUv04jlqqFDQ16iDtYxNlHTwlBqMvLp/qx5vfQFuAsHIEhRH7QNgLkfiXnjEpdi01p2BkDVbGhGx
uPzHHuvp1IiOQkKty/NLab0B+h/jpREZzt7WvwFEF2spoq5K/9FYeHC2Jn6DWJNHTYz1tshvRul9
ncFFTpAIN3TKu56mv8qjGGbjCx/apTu9bXgf4pNtW3Fg6ojESD3kTgnemxJdS21NWgYDvmcF5f8d
P9sC8rUULORwKNH1yyGg7ktYyUfyo2W1ka4/8CGJPlFSfV8DVy+tCSROySRp1uSGgURN52s3IBqk
kgBw3BiKAhBJkbH3vFclZ1PMmArePygq8zd6AswGaVqlVqjm0OCFArB6prJn7iXDMX9tCJM7fwTg
1gyUwbnvgmdQDYTBBPJBhMo913sWdj+78/SRvyg839lAcmIQkpRbp4Fr/I5Jnao8gcVgE4rpzh1f
gXUZ/Ydi/fADj4aZvtEB75VEjga3rearncSdrWjV3xusq4fQHeGVU242o1zDAX3IsvrBE0J7BPaI
sVdhmh4Xj+L39JE7ucgeUrganEpLCuakTtiWoy3Wc1psnBgEkNSpzTi7KR7vzt6PjOhXkOcQB4Vk
CXEF1kKLDpp6LMBivwcxmMWIXpYYv3wuDjuydV+fnnlfKI00R7ILdQUubBtTHjAfLzgrRK3GN9V2
wE/8fQUj4Mxf1inJzgL9B9Yhk+Zf4/IVaIcQAA2h29S6qyQ5nS2c00urxld2YMk0ERJTc4h8GGGs
yJIalyg9Spi65Qn8RHdvMhB672cWPxPGJbbBmaKx0Bp0dAnb3vqx9B4ljiXOPNOyYi/ucbbdOOp+
1q+XiZZsc0I1A9tj6GQfB8HBp18LJS65ZJ8mcD3XA4AjSagO/9eRVknLF8Q/gDYYSH/ShVegNs2N
3SjNbz3/x6IQNFMTOYbyv5BtN9sChrQwWl5OtU216VFk64Y+RgQM29ldkAjqlE/+mEl43Gg1af7u
/ZW+cHKgJ5Gdx2ZNRZqjQFuC+mailo3WiH1C3FQGTWojRd2DCOXSiJVz9GwQcJSOCzaqSKU1XGDk
rWBFTt4GqU8+1ufIjs4Cr1YsdnImMA+RX1P55bgia3LlTywCijDNLczXBkLyakSDe0pNMALNY7tZ
dkx3FqesWHxNPt7XEy1MdTpNcY4hGPabSDm1zWGwMWAjQheE5yWehzPs9Lil30MmMSHn9jgL2nvJ
G3mC+6waEXRVjxPaIQVCpmudtayKATnObvQWH7GD5cBhJRcVncrE1eRX+PjoNlEmdOSSPzCjvX/h
0c3BxHNPwTwTpYuMzmo6j/ztnXI1aQCTEbPdpu0BCJy7ZbIeNEbMnkMc7IOStpMM1EAseJUXmOk7
q+YzPluo0jHA18lyb90LesU1jyQuFvYwX2LFhkiZlps/6MoJWET0u5JQrmMbk9p7YaQJCb9QrH2o
1LrpJ/sQmTJ3ed8r6LB3YDHRsefx//8OTs3ibqOfY2/NXVnauzy77oYAQ1F7W+ONnoE1bOPs+c2E
mPN/S11yPyKZyUg0/mFFaU/vYsfo5kMBk9U78GeCYdqyyZGqBBNhsOWrdzc9MHF1RmwzqbRzu4iX
4ThTDORt7sD1R1+rjXIylgScFbVNJ7GhbJVocmj/3sv3DEI4Pd6aLQA1snquo0mSRql/ntPpEkyO
gk6yFOtRNkdCU/lmhrItsYsvoZY6F7TgVwfxlgbHJO2Asj/Qg5POHMCIl/wxsZKWNjQBzgQutAl5
rmWPmutS/abQm0CLb5VGOfQcgoxoTg29q/jCYAofvlIm1aBF5zrzennpOWp2DWGtcXJsMPCtf8Eb
7AxpCtvWczGS9M8+INC/rKAJUTjguduD6mUERyHcvj9BwudyNKju9yYU/sQBfdQtN2vF8KNXMFV4
4wFr4u3DT1aaib6pHoJxtsKCarY6iWYa50OMg3dKzGuWgvlJ5PcL5tm4yUn7VCm0kiJKc1iLno/o
nNZ4Gruolrnwfz1LtyQccSc4JDRhag9fwLnDploZcQzMXTfBKJx/Lh56IH2o6I+pYvesSWtk6qcm
2xI97J6KMzU6J8+1qLFtBeED7M4XMQPmUg1wimq5I8sOY1pNCXnuKXnpuj5lGVixDJ/OtbV/XjAq
eOnFiLGzMd+cnZE0/CmeBxocSXddCmEaDKAhq8TZlAL+BfIBSkTss+/QC04NejRT+FWtbXYDupmW
hP/Iqf8KihepisepWFKqgb/N37PONQ3FX954O+PhOI19z3NhCe2ZkyiachkJy3PboEhfdzMHMKHf
TWTEUShi0sBlfFKIlSE1r0C/5m4k7+abEeoPD3XgKZFuYtonYfTNqFpv6eJXWAr3/0zWzg5qbMw7
qqwJDhEgMi4FT0GnLOoKF6x5iyqO7HJzWvtAef/R4k6LD68c5v1EadaLu1RSrormqYETD+7E1fgP
fnRYkgZ+pzXGZF6WhdGt08yW5j6RT9CcVJEh3w6MomzelajMTnRo3EAzldnrmsu6S2u+pg6ENQq4
OQwRcVIlmGow3O4vFYZUNYw3fRBdcMer/UC59QnA6AEgStempXBHryyBiKU3y+/X6l9MdhLPHXt9
6Ig/neB91N9KwUc8GZ9xsDO3I0ZrDm8LGGU4fWnBxhjOyFDgp2I243Iu24MW/MuSV4ma5x3zyg5h
5iodJ7HAEwStD2cGQoSgAePyB0+/tfxjVlpM/ipR63DonedS/LQnQnddwkn0Z8Z/6dN/XbzjF0Nn
3FHYy/FTN7RXD2/7EWBavOqdjRrXLhwQJ4oJvvZTUZnm7uxGRUwlzUYU/13NF0RnDwzuftaRmO0a
wE8ZOeFXn8tW5MRbaNISVTkNtSglRsImlbs3tAr04jsXo/B2vardBrq8TVReiz/iRsq9zw2tPWV8
jkigbLAUQC3yLTNYl7i/WmKGQCeFlh37I4L/LT5yH3MYN10waKcQ8OXLnRomUTODtbF71JqmhOsT
0fYAiQg0g/79pn23cPuXKp9GTmjaveBkmLalmA08zouI56ug/23cWn+DztveDHfd3ERGk092HD0y
u3UeuUg7IHZt4FZveeBTgKT5Mhn3v0bFwm+H5kIv8EtoISIdeTNB2nKcqcmNZcPku0Gvp/CYcU+T
h7ADcBMYt22fnkgUbvTz+pB7crnbbVbHet74eCiH/o6gq9IV8VmLWJH4gKEdJN+EzsQBfsvnTZQa
TrDFQLNgjAqxJem7k231j/xzbPudvsSwr2MQCqMFkusv0pzzTR67WPUjVb6g7soV2OfB//zCjffE
k2+dJjwK3e6vbU2dXqYjfAznw4jeaLSn5QVK+Uv6aIeqiPHf4cew6W0Ttukm9fvFUzdnhQrpy1RD
NDHz0VJUuBs34hu3uddI/Sz3IuRX5FNzL2boSNgW/sWbfIFt5S6ziafzlUjM6vNvnUTA1wSPfVlP
LgePjmYipowjnhNkeP1FidysmuMuEEL0Z7m+O7hfshkCKM++4GmC59y6cCdf2xeR/qPhRm7Pc7vy
EVwlMFfZwKueTToWG0ce+SFzDVLqr1NSp8wzGRXYfrmyqMwi1qGLHGKams1zIvRTGSBsLiy02ttI
R5VVXQ31H50MGpAiXSh6NIgKb945jhhXeB2fg/ClxG6OKX1ssaPcHycH+PhaDMe71jKY6ilQKKAt
pan8wEj7x22MWbxrPPnggYvVlwTQbO5knGLSisxx9f8kMfGK4y0gBRqs/QLrNeuiAHExyUTYrpVl
q3978ylXDzZhlQ3IYoZRzcL0fU4uvq49PvSPy53zfKWY8jaEIkmLl9WexQbu+VMj98td1wX0Z4iX
5Zs7mkmbntgbaqMSbj7PH0tpL87OcUsL+lzbmmCh93he+zbXYlUfNDVe1Tis6z+P2sZaYJpQ8B25
gBj1WR592z99n/pAZZdaLQVzHE+gnhYiORssBH1jLzQD0onKjDdvEhrsUMI6SgqXRDl6Y6wUfQwe
CdUkXZ12eWAyKtZmowiWFjG7QS8IrSJOQgyykmwto9V/NmeX1rdozCXCZjvYepJGR7T6HanrtAmk
AJKHc3f0RJKDjT8W4iRsLG/rr271BlCiTxz2e+iblw2GADOV/ew5ZKe2DFCIkv7Hul+9sGGwkYbG
9fbNfkg5nHI+Z2RGi5RJy8X5HK1TaNif17c/oQNuZooCZHQKrlDICXqgZb7XgOtQZaxJyYdRZfRC
IVVubHv8tR9ODbjUTWBWhmvOdimLcnDkSz7jabO5LaeQeWd2s9s1ZKmSqLvBmpFTney1mYrNjEYl
CCojycmAFOUfYbJpZawqg3D5LPIYDbNo6pJdUXls1zqle8LEQOxQdYlfhZ/vRgCNgWo1SsxzmFXV
5fg+SYDEfM45V3XZpNPIzjJuMp9QpkNwtlljuqZ5S1AdYLPRxerJeY1b+lggOaIBS7gNf6FJ1Mrv
s245P78EGX50MkQgqzxdQdd4IPmpSXtkEFU/PhTn/Exfh14htzOzscZmeaKJ7UdiPxH0NN6b5QW8
BlKMcwUYVWtYO0aqd/W6K/Veou/PJdp4dWrR5Ggy1ss7UHnj18Nbbl0MAvJYRKkY0wNbg+Oemq2F
CXfb052hAS9A18MYxWoJlNQPAp8dYbl4d1P6u/5J684HYny8du+7W83qRM2uqsNVgDW7fB0pdGpB
9JepPeMM4a07IdHGw7QjI6EqKvQ/EVKVhA7RqIb9rz6bw3J05qk3wuBSvfioIheNY9QXUYmUvhYG
Uvo2K3E/52h6r7Sd/GhtYXwhGVfqcC7g4HRhtmQrRwHj83Y0CNrNyoNFwYlQxE0A4hQWq65xoBIC
x+GsIEewUE/b5X+kkR56k9KSMpP++FolSv15gyIIRtLA5LGMRhdk/PcIDAdwUT/QSERlz4YelBL9
MJhTi+5a84uzEPBlsEupqtepUXItYHcI4SFb0/MK3eu8tcI551AyqtkbyKhUreRQAYqWflJSzqbU
9v9EKP/vqgBQpyyFbd68N0ZqlyZcOMWQN8ovYOif76F3MNWmZa8WWJsIeXfl2jUQmcDiNAPXItij
s4TRAnFvsx3SsVLug3kshsFxBVBPK9XUKDFtXBLfJEkz1K1t0LlYNs4rbSMxnxf6zRmTt9OxMlHS
Z+EICeyon9cMK0g37nvEwxnXo/uKZ3MsHIpQ+BxUzQOqEK4FEhaTxESJlFEoKv7vRnxJBgBPqknh
E4UETq8pmhKJmaB0Dokb8rELIAcqtYOuItTizRErxuG0l95HC4Rk/gykWacTmzuoPexQi+NtheKM
D2ltszZHIfiwp3VTGnNOAAdl39VOdRQpkdaLhGD/lAw2XzW4dLpD5Dx/r22hQQ274S2W5Ei4orra
wz5DVCuUh0Hjf8YLE5SGo1i1lWruR6Hcc65RvcmdxxsIRRnKKlgRss7m+eQmuNMNgxOyiymgnqff
V2fE5StRBiARaGiKoQ5xKi1/+RoE3InVZVwXKIvU2sqtMffFyqXZgKb2BJMOzOA9jivTf7itYUEI
KAImz/tn81d5SaKrV8Q/ev3T2PyApeC6E0pEl6QDPkCNZBfKWWKlOLTFug6WfVXXI/FO1Wjf7yS1
pvk3B1NpJOpYAa2T0cCCzVbhREzPm8en0Epl29HxWlWlj8fNEmxzZFQJASPaOEzOiV6xTHpVC/y3
rFUpoDNQFwRnIRWcT6ILNJaLBQLrJadrtkdPUMArbtOMHpKLjSxFKCe4TDhaHQL4no9F7vcmXI6f
fRi5g7vmxlUllpr/Gc+G2UbKNlreR9bdf/gO7MNeOzt6DEyvOd0xu3siDTHok/9Wkrxy0XX+CM/h
auGOnAYZQFtQeXgWMBS9FAKFvV5yDOiWtnuq1PWUxv8NbdQaWvhIfh2qBIzcg/Fra5Ct3Y4iWlBE
i19S/9VC/LI7Lfz5aA5fRVB7j06v0tatUyoP0wEljNV/jrOvbfChEzDyqz2vvBRI2etOScJ6wRnr
pCsdf8ACQAV1HV+gMjLWsHnq56w16Q8ZMqerxYv1hdEOGlnW9C1u6iPxL6J/jzQssJWExZaDOkKx
nPkrgC7C/kTYPfroOSRN2lvJ0cN3FwgqRcHVbGfWJoJEiflb+fwrjndgsbnSIfRdM/GyjO77TRcu
c9F95zkMLsXWNP0HFKqI6aK4wnDwftLM3SDjOK2BVXF10l21RAc9cbS5vTlXCnyZCYnHrvWYE6xo
5GvU79UAiSIMz/qyWodJo8SzGRsHvB4iATqmrepEFk2TkdG7DemYQ8BS9l/u5zIPwQqY4SV9J0jA
zpuEjW6ERMzuWZfa4EoEanA5hZJFpe/xP+SgJ+XVnCrR5K9vwRMrZM2wzfQq2hAf4geBmQVkLGIY
/Yw1kOIx+1T1EbI8Im/GpxHWMsH1E0joxADcHFRt/+pJEcZ1PIMRf25Ijj3BnESIEnTuD7/G4Tvn
/Bsxf8LHyUGu2f5/+qPOrmk92NRY5mswUadYOLgFycx+sFNpg6lB+Ma0W+HeZVXVslDAIBBTIauV
Vu1+87jKf6/tielsPOY9lNSiUDHOl7FRgFmNXkIJo0h7VM4EdwY4+zIeOG//LUqxwhAsX4OY2VPk
Y5m9OFno4OhRmHdyf1YKTz1qRjuTKNo+6B1eyvu5+n/ID4t8J3k51MP5Uxbr6DEQE4nv5ZT9oBKs
XVK9EuA14WluBfOB3PtY6jMAL+T12KNs7/8ZwLLK7FwMDhnb2Lk6ILyIBIXk/Ax0AxDjY5g+Wf6E
bVYGfrsgGF0uAw0D62XfkdGiCsyZw+EVEXC6hngt216ecCHSTWQsKUpTns3dYyi7A4vP/yH3tTyh
3GFavJeBK8zvgC5WyBQHlTVvTWo2AILeDE+Zxp01+zsrhaZDqsihXQe1AE5d03dfTXAo0hz/eAGL
JuAUJcRQDTQueZX9wSawT5tK2e7oFEPgfXrKaovMFKVTco7X+4rBbQeF46/dzLHbHCWovyGcJlaP
1/kT2i1mPVb+fHLFn+1fJ01TP37KvhbJW8Vch/o5ZU2MiJsJnq7B65OD6ffFSggtS6JE/qXLfyaZ
Z66yCV9IyJWYLzX7hTQAr+X5R25zgBfusd/hrO84bQ7Bfxd/+RvK19nbWNlONOEAYpamc6Fo9LvG
8uGGaEZRM/jpjtleU1+zjugnEbsmdXEtO5t1mMsQ1Rqy7UwDMSaX8Sd58rUrpqd3xBrGBUs41xf7
UlUxX++UawpR5JL0iKqcRowBx5bUKvvTIJ3qSkrteL3LRPbnJhMkxvfWqAiBEDFctc8JAMHaU2AK
Cb2UzUtVj4RtyABkN9yDWxcDQHhvEUIPSkUrLw3PfdFesuEC0KHnXe8YSQJk3S2wD14mD+zy827O
x3EJFu5/+HAGM/3X7SPUodOt2uba/GcXY8+B2t40n8Id9H3tX+xyzJa66allKHeNnRkmhsQC5vYa
9rk5MyiB9nPJf1H8xK5CbatxmC0l6/PFJszhWVys5N70Do4wfOZhjyIx1mB+fTY708P//U5Ptf0t
3t/Mui4C4FHHhgrwkPb78YcLQMsX013L7JcS6Z/XmzRpaUOrheHkiGclgUrL84T1TEPnSW5CRrmN
phNJ4wKJzMUf9VT0dTcNi+5iJpKcJ7WvQr9VUE6rcAGuqehQEACnAAy/8jcJD2MfpwK9u+mCsxeN
IfKwodJ+rU/AydZne4CJHtB/UM6OsOn/UxBA57NOyBmrH1QhuKLM3a7S4B7r7llpqNlgyTfd2HUI
tVpUPN0e1sbl25hDomN4ApzHqehbGyZzSe9megtCNsFdJGGOgxXSsussQuWtjlVKjElzYpGwQD2K
LQ3Ngqwj5t+h16zZGByj4vSNAnthnG2XHxkiisB2XaK9YQVB9ZjpLH9d7nUhwbQkFRgHOYPwdkHm
DiaeaEgsvqo5i7Ctze/xcFheptvJjvB/NALwdv3YLZ2zCA6TzigPdxvbL7pZzjKoqy9OXS8xCTVZ
qey+IaKgWxF0eRNf/Zf8/A12i6B2VExeHWFwOZ4cquh61B5RKnMvyl+lvKaIqdc8dz3+iX7u+aPn
7sNwS2rlQUZm9RLm/9PYJZcuwDll/d5UPFN0Oxkv9zxMpCPmPYZ8d/MI16ufwgu+6D3kD0ZAUz1N
3grbqpbGrK2vCqIJw5nFTVt6jDnm6SZUzizEtQY8NGrgKioh7xWDuYrd61D7g0Zo1UCHU2MlhLyK
N7ZKJmTwNh36kTVBnfeePU/iPN6h2Unajj8obBHCZ355JyQ45u277tQirTXIm+GZTxSCTY0tmpdp
UKNeFBzrLOg0sUJRbpsE3drxDoMaQsrSTKy8r6YCcdKsHm9Vg2PfsXoloNXR/fOoCN9O4U6ad34O
EI3rvuazDKyoxNdOV8eZAKlqh3z771Z2mjveJ7+HD9HeJs4Gfzmv7aKoZfCnyaikJ12eR4auH9LJ
Xiyxndhcgv4uKdrWVkQuC+6HCdgusmUzWyaSt7R6z+ZFrccSnvelHpb+ckp3SREUMWnR97OYQXB+
/9icgmzILYkV4UqjyVAGqYAm/dhzZ8e81gndKarD74OYldkGt/taL6jPll/5tym3I+FHnhOFC8zR
hvBwK4gS8iIQU09drIzVpOluttVgCHt+RMhvuBDFThGtDaUucRkQCbNCAGXS6UCS2mgg5+ayXv6y
6HUyDLPHMpxjO6H/9ayfLN2oJiI9UrFTJDSarK+DGQUuWxAjWJ9v+Jy3Vgs6bJaOrowljC1uDx5N
C5LmCC5+znnK2jALwiflomhb5Nrp/sw5gUHl4IwXFbhQS1qF+pKEGmD++bsx0oR3cWcZ6cZa4vrv
EIeyzqPXFDI3KdQVqmbnXys3r+s+CjEeB94Tbn4GMiEAUNg5hNk3KJt2rx2R6UYAYRE2+SpG5gPZ
m3de3tgvO0Jb/Kjsp0tGrxIBo0k1Fe0SFcwqmp03kNEso8juP9ciBcg/nz+Wr7qXVqki6xSU40VW
iigM8sZiaXjuB3v5wGBUvV29n60wrQZITvoCI8KWF+d9zpHpnKGgujjROKbYrfUtL/kDyjigCtlT
DrOgp0Abd0MrH3iyBfLPCyLJCmChvl7LN2653FC91OO+6Wu6/a3UU3CFGWpHtnbkoG4nTYR8yW1h
a4m7WvyZJzxExRsVEAOuMhgunjU6iVLskNsoAmEtoZoTcAZ227V006GmDj/Ncdmni50fyf2CSzWK
eXWHrndFEfd/5TYA3aTjlf93/MRpnYEOHUu6YF2T/dkQ4fKUGik9TumAcWW8hiaNtGcFoR21aBq9
Yatx+Cl7J62SawY1gnN9VatzKGIWtNYX1/FE+v/CKbtjUnZBuvNW4yZcq8iQh/B4hrDf6WwAiSCI
Bk7oBcRUU/fN6yONX2JldIjSmfXuTXaHQtxsag9pX9VnwAWW0DaGKQEBD4FevD548k7pCM3rdInQ
77hTDj4tZiJ8AA0QGjOOfpszNGYghYnk1ECrVO31XoB9na1rSpEZGaVBN2MjMGWdoKZIcDrr7fSP
Ul/LwrG065JUTgStAAKaVNaWFfan/chEjXpjqah8Z24yv43v2jPvG7u0D6p9MO12MTj+Hdunym1D
lzo1883zRsa03J5Vg/7+ec73lrtE8IgUJgHXzRnbDTADceI6VVTdpYXuomeA+8XJzmD8pp6M64os
JfihvB4rIoS58boWIw/nwALyr9vhLK0TdqdHscX2uy8l9zRZj02hu4Mf6mJwbGTi6XJ4Pj1nVQf7
UszdN1MI0G+MkEEdm1goTwF827QZTFexg0mPviTNcJoQl/lQwzvbtaan8upMRG+aiaG/TXeIrvs5
wRKpzzPpMxNX1Zd3bQjmi3cGInRvlBrBGLwFJ4dZRLj6ZtaY3Tgl7d1WglL+Tf+o7yBN3gc3MAwf
zzANRZm+8mcgDuZlGRaHPPT0xqlUdCw07fKfPk0VgyZKpvlGZM+5g1w7okmZIQnHv5wWuuhByfkj
P3JFI4N7Rr/taDGsWC8wDgc3eqJTJhNJEBzesTL0WOYkib3U50aL5FA96M5CJwC0oEItjFHIr4rX
7ir+K6jIFMHGBcDHTj0AqGMWof1+XRKdRNxKMha2aH3cHl12mCuzx/voudy8Yq9joEoiUeMZtPnx
rzz/zyn/KORX9cFHTHnDTQiNxRJbhJMBBRjveEpardU9V6PSDdtUv91/iPKX3shxacoQJiJ/QwRZ
Prtru6w1bNFNRYyOFKYl8VpGZ1VFYhGZVZD+nM+9Nfl1Bb9ZEj1z4UkWEvxu1PhFvzi1kC5/1N8v
0ZXOXtirzDuAluH9vYfDwV1RLfmrS+cZs0aaFCBHWjkK/5x6OP3xI3rOP5PAQ/84HTtkmXqCKxrH
nEprV8yV5447MRoqU5b9rE9woMa71wP0uKmp1DN4gpqFLMuFGSNDT+C+fd+Pw+fmzvFaMPQXZ13J
MwyWluZX2Ig0mlvvy3OPImQtLSKJRmsC3ZN8Mm0y91wENeZsnFLZVISwCNXV90ZEvHS8FXDgE5oK
v6RyqO4qpZDYv0kzeXi4z0KZWRWRKsFqYG5HkRZeQwpE8YigWjos9YpZFZ++sicyUCVfn6a+dDEQ
ia6nqjiflsBWjPrZlh+8nJmASOc03coHAi3TWf3ieGR52l8wWparK7VtATT7Bd9jH5eYU9GHHmzY
k4motaNF55ZHu6AU2kbWpKTIgHnuZuzMInBm4oESF6Vo7VJm5cTCYLG5qD86SvTOMR8dEH1ZTp0a
epJfbxJG+3+VEMRZkX5HLdZ/LUJFsKfhz4VPkAPJCiaSc/4reC/Y3ktmcIZbbH49aX6FBoLwdfCk
EYPO+g4c3wm4/XQAhnhdHjDzqORe8rK8wwq5QsO7GYhYzaUNav6rXjaLjgFKZiGbFYfh1wnAA2vK
LOHDR60DCfjqE92Lld2sKf4ST0Z2ms8qoIa2XAnAmeR/WKvTeADMLb2h0ofVWSTP8zc4bcsnaxNb
ChvZ4Zg7afRzMucWRi67FzRhE9DUsXRqaHr3+H4VhoucByttfcA3U4Lm8BKDhk2tti3hsToaaZYl
uzmN6I/myXYIwAXs3g852/ywgxNMOb4To2sTkxQ2NL0BQFfd6mL7yl1mxgKA6MtRgWFf/zwnOyeR
TcnWQxkUiBWOIo+x2uHXzBQwuXHb4Ml1/gR499SDZf8hJl6DTkbXc4nTnZi+CjfJRG3W0qZGJNFx
zSYf+uuM6fWibbhqVkoI+VOfnEfgQZ8zq2zM0xe9YuQIBQbJa7BtSumDmlDBI5HGlgFeRBWRxouQ
HWbu2MxiAkWWBHxq7ztRwyP4+4KlcEhRmJfkajKRcMkqED62Mr1o3uq9nUBUS3CBWjqqQ+TzZS4m
36SvfHN0p+rRF2bcDTGqIO/DjErp+U/EG3n+A4iLKAtMO3Tnpqiiw058wBkrtzTVYZ9cmoQg9U0n
1t0y0ckbLD1Q3fQqoTylil3gEqEops/JRUuHLkj7ZaXcfPV/E4GlFPHJrtwpSdQixFHMRYMiR5W7
4KmCp3hxjRgjsF5ZuIaa/cvc4rCO3ElccNl48TYWtBzdownKgJH+u796yDoSrf+QWviMp3fZ8o9C
sOm68AjW/rbh+z1hc32L/nS1e2alNgiKFz06B1xuwofJxMenH/R8CyU0+dvYdPoB2dkajWKohLWx
3iuhVjf2+JmTziCMJkiaEMgo0R2PULEm6qk1S85i9MAko4g7CxRcmrPjcjJ6JeNnfZ+trc+gIeip
xqL6t1i6CVLwFCgnp4MSnpHPOlNI5YTsF9IKJdlp5d/YVCjs3srBFXcs8PS39qOR40FGqFCmKFGV
u2bvdFChFcukgB5PN2X5lOdKqOoJCVsf+BYFXsckPWqJUHUjcaIaeVm7VnOhlVKQKesZzVgs6u6a
GVrFXwuAkFruN0AlRyH3q1fy+MpS7dXRQ65SI5DJiE8YP+oT1i5lS7gVrk+8iMMoJcPxNWcCeGZ7
PLn9G0dxM4AeqfXIeJ98t2tlkyT2hNqNRsnGeeIp6UAzZpbrpDsByezxo1tKQKITChP43WG1OfxP
1lX6uYTHetDHMdTtkH+AyV/ZeRAjmDxNT0+2ncdYkr2CUlEqhhNnjO5X2iHoENYBpIJkls4vNMzq
wdVCage3BBbX7vlQmt0Fuaxl2Pb5ruULrP71njebngtl7KUMd1WogPlaa0dKzdtHKeXzbrIOUioB
GryIaL0O73/SBnqkCaXhxYzpQtM/8fSzqzKwBuBMnOPbUfPCwIaXFWEwy63sXo9Sr9C3vgyehx3A
6xAfzWFDra1O4h7Yx5rOrki12kabSYvdJUoGQXmqmaF994jIFm4oQM2T41//d14JkLNXoJTYSNRv
EdAgcNNjNudmK9Q5rSp+/3hqVWo/mmkj7ckqejyQoDBQOu+CuGYwwNEZkwxaDtgchzpLRY1NXy7N
BqYM/749y9uEm8Xd59vRQr4IfoeGVn40ZpiWZWq3uDW+SFhO9P6HVmOndauJUpiP9I9xNyRtk9r3
QfB5/qy33yK38zxF09IJsLgQZpQlMXws6iunK6LD5BI5UgwJRhUUWgLQ/J8i7zxgnROR2cMo5qi4
Jfe7zeGxvIX4gWu7YkIjhz8ylq+NpCnh7cNsnMlGJkIsnMR3j58ZrV0egLcbFWfA4byqCl3KR+vp
ZOD+uzTTPECsA5IeRLJpySwb3O26vAh6fQ2jLN/KNFm6vdmouT1aJQVWi2x5w14UAKS2MZzEVUuh
xAj3PWiAKWUJkcc7RC5l+DpSmtka7ir3TeGDfKvl1yudzxnYIhHrsBrG2iyyEkA1qvqQUiq1/CMc
XlP/lFpw4HhxrRanLu5ZqECsxp96EvTww1K1PxkOiqyeuXGfDO0EpH2SUhRiSwkRF3wPhoZEFAbH
+Hnjr4DtiBl9VYercdkOWPgqOIAl0v5YG7ojHQvcgRu8nDpvgQma5DDHwzP34HrP9RpwdigSs0U0
88fQu7WbSBl8Ie62x9myzmN0PPDjhwyOQ9f/Tq9zR2OxB6WlrsFjwv1SSy0n2xjCTqlKqb34E+nA
POGdq2YHQpg4lCtS/zHCACGHwRdeMPxyhtPx4mZ/6mQGp6/WFABNf5N4NqeqMP4HqQ+8gWiZ7JDL
OUmoUuHgdfeSXaWYSq0SeEI8H+m8ujqWF97IcYcQ3uWpBTCSIGpMyzdXdYtW5rAj9U0gxNib4VrM
VGWaI/RBNb3VRX8SSSiLHAFC6CfUSxKeYVEReLFDS7+m91WYKGf1hZeWtgNaYLxaCypqsgAadx5E
61mk1wFwlcoQ4xqswugmJ69OBpZvMMMSRTPLcch/kZD+TleiNbkUipldDM7EilYfv1fiX9JuJv0U
F30OisA2Q3nUmePtyjI46+a4ro7FpphLtnrdf3M5zqKp0P2d/azJT/APU+4g8Sam87y9zY7VsXmY
sMnXcGQ6Nz5vpa7nxcLHacrVV4L4Kcc9IrigJ5fJLv/8QGT4WpF7IY2jHGKojjG/9SL21N0/dSCP
LTE88//hmC+y7+qyvb1pnZBfynpxv9NUbrW3BDTmG3ZVugVYuSp6z/xZNiLXdtGZYZP1HbxKeMrE
hZz79XGtg/tMldZPGyYWBX+BeBbz9K3v1cWCrD+iyJJ5k90Rff9Tv1EANfHLtBiLJO33fluOHgOB
mPKQTzU6ubaJErU9Gla27eCnv64skRTzNgFg6mthVAXqD+2HMTfFUVQvFkg1pgEZWSuoLJL/OPGp
RZakT9Wspj2bZeMX0P/wQ7Z0EJ3Jts9rYX2+ZhDLqHrGt5Re6/mv7Q2FIJQ2WduvaH+e5f/1a+zO
Z3NL1/DZH7MEWtpEH15vE120aBWR4+DZ4jBMJUnC4quso0VV/kgV3m4AXPHUS4q9xCF8D2C/I0Ih
spJPLq7n01s/5E/IPavdtwq2D9hcKZugFcA99G1Xt/2dUWCXn803r5FAH23illj/zp1xk7r7eIqh
e9kGeCCJKg+Z01DORcLS3OUXaQL74TNuMjEHooEbSuf9QefQCPEOxHN4T6cUct5PPOi5m4EFm6Ci
EjG8MZiV7MWtnwwxZm+54aWNgfmB5qlO7s0/hP6I32PE9wbToeef76SJ+9ZjYP1VakdRFpFuBt29
6W+sQtrz3KWtzAwHI2bbiJ7XBZ3qiJZtLwKuUSeLZlmtlygojCvPkBOvTGJ3nIbWQ0CcBEOwJuRO
1hmgzBzQ4/voFgg7d1rKicIaDpREJzz9AA4wMq806Lpd4M1OBMFyAwgqAI6aNuk/LhNFokLA9kzB
i+J2Kh58lVTYCvswfWh8xKf8gYZD6pCpBvFLjONP+DYzT4GkxTy50a4WnArGMAHj5FOqU6GIV2ze
vnlBjvc7yYRlsxXBnx3FyMDHNPKj+VOVymgfxLzBS3dq10ADcfvCsYg6bFS//4UqiA3GzFcUFZ3L
oZEjb0SN+dyBH1enkCXy5kp/NGdz1kUU2UCQNJYlzF69YHLTRe1d/SH+3VAoRFgAXhaU6UBiLp5+
SiP8t3Un17s3AhMCa83VaSWGTVJwxukPI1u1YtyjKwDDYavXAIr8N3ftnp0JZ96Xw2dAn3oB4F3+
umIySl6li61tMcaoUni8MnIvmZghbeCy8bVShJUyzobubKblpVYTOuYGnp245frbyHHpzUzIhbSi
LaAhpZlftKVlHaBxtdvRiFENqEydqj+ZCvYiGp9TqfwE+RLs8h1VB+o+QEKnhzBMLaCeOxRlv2n7
O3rWf6nWXCYgkss4vEMKfQOKwawQPrF2JHqAMkbUADlYtMIMq5NJfYXWEjjVhizGHkDqxzlnR+2o
w3W6VjWaqeA7knIwQay07XgmUWA4i/SphDwSniY2hVtypF9eKF4RxgOYzX44KeO+Nu02h6WfsZcb
V/DdKYcQ6m8HeOg3YYkonIF47jBJZFUhEpyh7U96xdAAZnTjMk96vJL3PnT0x9XsiFLftGGe7KhH
zh3vg9lfb8wXaXqMTzzJ2Zso+PyArKR3mLsuY58tsXeTJ3BiDuD170dWThujtIrpP/38f83DIRK2
1wU5xMRScIWQPjhFxtL/VhVgDDln0zmL/rmp9trt1AUKpj99xZHtXwx+1pDv/QVabU2st/kapnb/
mrkbbAZS0Ud7/5OpEcrenMjsGPXZP7IO7UsNdz1HRe3MS7aWIK8Ed/u9lzhB9gV71CcKF8Mf1Uq+
pqmPKeR9FN+9c0YzyvHftXkz9Ol+hMSp8c3KPtNUo80GJubPTOmdRskCnHzu5Kp03lVOXhygOWkm
GxotKZ3VdDtFKoETqf0kSqnIBtzILlzHJgDKHPkn5yRm1H4jrOJlmhpG5J+gIG7T9f4Bt3Kmbfg0
CjC05H0DCjCL6XQTs8Lia0KaPw6vjo+iIwZa8d6BnD7p1gIshQiixb1WBvazdAZmskWI3uAnf1ap
zXuAvkp4nf3cjGSGyGVlkRTghxErH4nOENSm7yzPRTt9AXpbY+xG8Z4XSljENeynZC+Dsvy5XD6d
nSZa5lNdRm92n8Z6HCPh8iB1LUHoYh51VzD1W+4RATPsH9Hvjhcv0i3w17JLkZPiaqou96jiDxxa
Tu9p0h3B7e2pZk2KiPaTwkelZHpaUrj3mAwMCuWnzPf8QPor/XAinzXSbLu5BrV/kOOYal+iZzv1
5Y1ZXWcy99gfgwLCd8K90PoKb5e4SMkqjQOlTpdqkqFLUi2eBzrtyvYERGcYONUpOOLm5rmee989
Vll3SSidsJIaMQdC9U1qZDr0Jh1uiVKE5epJ/1DW83A+6M3P3d7HBnwDlkEdJxzYgwB9/NG7ynTm
Wvg0H9w0i0WSLvj6EY5DRz1urlaKvhz2n7AFdCKuib46cVsxrPZ6BEDCSUkoq7l8B+qskot1Q6Uq
1tKY5v30e7OSWF0BZUjM9JRz3k6BMlFSmKIdlaQERNm1/NjFmmzsau9kcn5M5ZoO0SFSoG+DjBfx
l34dTdbd/ILfXEkXt54rhkwpxRlCaQvY70osFj1NswgUeEArkt6kPVygGQ9GxLN9wa9/GwcOx2jo
4kAvZoVmqWBZ7FuJTc09iNbNBMHqAnAz5j2Fo4SSq/gKZFypxrJsYuHaYHCeXjtzxrlCUSa3Hfmp
cUThjRShPaMVGI6DwXQKyZqLqpUyVPe7EwsInZMbeZC6V3Tv8zgVy6ez5tConYjMN4BqW2IorlFR
dwDNrWLFH/AIrzqddfcoAFetEl7084I5qzUCcghRg5L31kaxYdrDxie7gsnoggYjIFEZVxWK33P1
WCgsjIAk1Ej/yOh/Q3MOfRzLcFGsx5+/X/eTLOnzMYR9QxP1WlKKQrwN3Qi3o3rJYQEYHgR2kyas
UL1yB24D1m546g8DHZblwbVSj0UcWXZwP9Lvv9CrAalcGwoedmo1oCc+aAknc/lVi/7+9PPh5X/a
A57l//qKL3A3eoj8ml4HVNBxtkJ9pvXJ00L1k4vzG5FPTDkHuxAdgm7SaiteIlu7azJKhFWXdE0c
IXQl2bYRKcTzs5tEd1hpBBq0dl/EaYOe1L9cioTeNIaa+AdP51EDESkAQUGzKZPSakAepRpiBYof
SSZzPTyLEflPaGSWmJ9FKOtVlFwlFPXRia6jPSuPwtGGBCDbtsh/CwM2JUEGTwtqHI2/+YtRwMyA
T+lpPeSTsizdE78BAQc1Gm2RTTAjRJPwFoFif/mri4fhcSJv6gqlzYOSDPbYHmm5aNtBHjzQT7Jo
vaiBLjQBPGtgy/F8TPfIQ0fK2lq2Ua6slf9IjY7obRrQISGgyMTgdjZRauDv2A6lBe2WGsnMSGNv
Y9YlHW2FITN0YTQuNiM2c+aV8wA2sr+vbBKMnLcZbXEuB+/ZdxYq87f2U5G9HS9jCVIoVsDAF+w4
p7IMIZkMhKqL9BGcihYe1uR/rk3Tjn2kHJj3p4BKpWG8rGhwaNkuL/R0XhlZjrOMxTS/q8TIfU0p
nuGraDMOxWAH22bujkORfe6I4UZ5efFD58yfWSmRNhfaZGTAWM9pDGjgfQKY4w7RvnefTsb6mJNa
uSsGbKWx0hOEA9PaO4JJHvKJQma1vB2AmefIQcyW/s8tcTtNwSCb9033kat6UVFZXmOH6M+jNpBR
gawRHwg2ScQSlr4mGieXKnxw0W+/EMma7t6qjHEYKyxJ+jBDlxf+4JpB/nVHHjMQFN9g7s61WbEE
pvXV6xH4w6jTztLnGydYNJN37ajebjWYKvOU9kV8uHYSDwXfZG+pdWj6lYY4/Hnj0rc3u6xElNIG
pEgYCyYigQb/LNI/biLOBEyfED6KbYJ2AiI8cu4mXhjrRQ+9VWg0WypeQ3aUwmv9IBbjjHjzvnPu
yrK3iqpRYIIFPTAxFVDvk4w8+Cg4sPgN4lByXkux1pjL1zbtqULkC8JIUqXRN0LojqiTxR2XLwJ2
tdzkNaAvdwzChDW5f6n/QAwOfaFUV6iuEbWzSyskOovfXbgfbJlZWwcck/yY6PmGRr8davhR/2FK
fHsy1ngHNiBzOASW/WM4NoVFanWGl7McMNyoQxr14OWQlU6rqb8jCaDucsYsjb+Ymy5QPjPqtIGi
Efp5unRWSo+2QAo26koYRh7uf4ZULx6uTQVRCTWuWPXaQIoEczb5idPZMhO/VL6Ah1HW1cQbn99v
7GAP9/rGa3a/66cc+m4I9jcuofuQyOfu+qSPB76eS7B3YOb0qw3gkx6smEfpLo34n1ZSNg/GjG3/
Wpg/hr7yBKtsIxK56RW0QcJMONMl76co1kCs234cIIZgJAhYEj3cH6/jAN3mIpquI0EBDJbV8w9v
7Lip667zFOBAtxmJlqxoUvyLsGkyShG8DFXuhcZ3luH+Vo6yNd0xpNHHsbrnL5lG/WeWkvSpobMB
M5jEzTqiTFv2RjtXSRbFH39Q8fo0ZVxRx9zjZquF2BETZq28L/OLyTu3ZQy3B0YGUppqBbVdF89Y
5/GNk8rHpyuLF3+Pdz8RJ1beewiAxOQ1/eGIpzZ5+x8q7b9OUG5gfjneVhdsMNZ4D1tMmYQH5dUd
GetBa9fdlQk4TooNIqgLva6WPGixYECCymuXzhaaAq7gOCNz8GT7lsWQ5VioT3ActoFj7dcU4i5E
aMN+1S3roZWf8FjY29f5W/znsO8rac0hr5GkFXfjrezk1l+A38X/9BZ7ShduRmAe7ZPS3U67r3Uf
vCbO7S6HxJEqZcVLRJKZtBO2Hc7TOEh7tRtXVqsG0ZIV6QKsxoDTqbU5x4vmd79vTBYmxvqvEHIj
r0hZq9POkF6CE1URNa+pQbhoQyJgxU32+/6+oQEw+CyVAyu37xxD7svFPeWjfQlhZcA3tVLiRGIp
KoYUwtrRa/d6htTn9X4feD6CKqlsMam8LZmly/Ppihn+4xQBBLCVCgBL8TgKezVCn1GvUm6xp/aE
4wmENAbTO2D0J0Q13ftzra41Zeh9DwIgtJS0kC3NfINGxYDHmHgVt0UxKAqazL+E10YJgKCtwFKR
qo+oIparDl5ZSqmDV/yTx8YUUKtsJxtNGCcFTqc0/901HHO+tiOYGmTmntJ7ORwO7hYuTBd1q9MY
ww19FlXrBgdQ+v3YDOkXz1h3PU9ZhNv+AJhbsrI3cAProltcRSIiu9LkCXSYFS9eolMdl4+Z8urS
Gu1zI18HGrBWgm30NiCtQ0o5ZyVidmyPz/mQ+cZdzc9g3CAenzFfUKwBTGMxDP/7m0bzDUwDjHBY
QK38XwIgAitY2pPuQvjHb4tCYwOQUnQNErYB7IhXnqX899ag4C9YDqj+9DSiD53Bb/ZQE6Q0BRrk
HVCn+Ux1yMU1oTyS7ET49SkWkKyrBIcokJBHx0DtxV/Vyv3K7WTc0qMk/doWhTO3uQw8lgUK0EKo
DC1Ho9ZZT3+0bQldfklFsLISnZBGmeGKryZX0sSsu+wz6QRFePzby2Js/L3rcbwkq4AJZnYbWvBB
oAbcjhi4+e1Xfn7AUfiuyvKadpu/2CkKO70yXz54KJi+jz2f9J4vnWNghYU+2zPwEnE3Gj4hmXHZ
xNj0qJSzGeW5lxkZHOX3rFgps034CKd9/MNJAXEIU5tItRgYkLoZm2svxQMN/m8ys1Y+2ye3E+tI
UjxTNpVoYQrpmV+yY7wMLg8P1AbpAk+AQE/d/8cGSRf37qTT3AoQxOnM8FipfILPx4yHAKXdpRg9
cQz5Z2K6NDD66CEepoPxDUN+uOjGjGjOaa0V39CJ4ryExwa0yAI2TY1LEzIkrgKodz2GVHmIfi2b
TJf2WVAgDIxax1kwc0uFywa6CWwI2YgETIPQkYMp6w3XT+OEvX8lqp1EZp26yYs+eZ2MLYK8Hlw5
pPz/Re/fUD8jTJOtJ15H3hBT5O4sI5OfH8fDoV8aHyoSjtFA4lukdCiY90QSjnPjJKs0l7KCaAEI
mRGGawVyEW/fGEk2C9UPajRxEAXD0ZFyw/dVyvGg2MWu5aH1y2Oz3cc/aIpdDHtRz2hWWBTwdkrC
P8puhikTCgdq8zIyd2tmwDq+hmLUiFCEgNLkonBhmA0xnKXloSDrNHYn37I6ZDlIOlqRFkXaZyxo
MIKVgZA2HNh8bqvu+bzscwwO9waQKnPev53ngyC7vrXKcee2wzxsbZpuHrzx2zkJIagvrlYhfWRw
gDomS73HWTO5CPKgTBUYtUrbXnmuotVM6hRJCItSdNnqQEn0TKPuNANunpzc3ol/u29J+hwXu6LK
f9uFgI0lhG3x+SNALseB/oBGyT8ap1iJL45zuBqQJF9uJan6R3yAayddRnYBVDwReVz0EPfawWzk
m2x6ojmTCeF/ZRjrZpjnabH+klGIQHZZIO2r6GrpHwFpR424HoxVkE1fKz3yq1AJtlAYEIm6kWoS
1JMw0klgE783vDm6M2SNhJAU/aYzLJjr7wGC/ktcu9GCpRb4UwrPyPF4uMKWcRjWdevjsJAwxObL
hd+55WdrP6WMdPw4jA8UfYwybPEDrul0P8AGigTey9BfiqtOj+8v4b5Xzysw0jlOH0z8UQrBOZ1b
ooZOTDJ91LDsZOlWVdILaZTsXnEqE5NQXXhj/tfHhOwgHNg/JTWqEh8TCHklqBuPRI7qQe+WwqdL
jjqlK1UXTRi0PtyGf4aA0rmGckHkckTfW9VTroFqwG83NvI4HC3zJzcJIbhLe37Zek7n4M8a0BXS
jm091TUd/lP6Ufb/iBwTqpNl+ouQNBxb43dERrYbqUyxwTCXGKxWjrmvcorh8IRxLT6icfaYwZic
B7PAaFbLzUaA9u/gL+SpXpYO+ewP9G6/weU9ug+QJDSVIPdsnXvIssZE2dSHGvy96rjebC6Eo5bO
X5BjSH0OqmHYJKR3t/i1QYEYQwZzVQQdrapC6qRS5+hcSrZX1Cpg+iCM00BPfxyqqvIi5F3jV3wy
69ukjaoyYVs96N/YO0xA0IL1PlQmZdeOKE/F40JC5NzY7haCoz/oUGK0IvvECdfelKLjoWfH9L3D
Zm2Yd+TV61IYg9YbEW8TuZFxkfKeikE0u2EVPkewdxc5zJd2ljnPNNGpqW8i/tTgMN5Vh4dda7Ya
N0toAXcJu9/YbyOexA0VVIhJkmdsi2TEML0I4SR2ZgjYE2MKZ9w49joweItwLYUXGnWCypvvzNZN
hqeCPzHp6oT5rp/MEKsigekcPPrAOoyQu04xjIKk3dJ1biE5+gZJHQnTBFny0ZWe3F1hGeLBe7qo
KXnWXlExATVNXK8y82zag592dAPP3QwdFnL5NKWDZDQtaCIntXxsuv2n8lN7HtXSj+52mA4aCFP1
eX0bi5KGZcreJCet9HEWedjNECBmDz4S+JlqRp0yqGTOJYdhdeG5gIofDCOgNfM35yzKZkTd8gbt
ajvxNj1fte24zXXBnDQ9XEm1P1Sh+iWZ1KKp22mF4ypwzY1NJyjVhoYZ0Bn5Zwt2/yOiBbQx7Wqx
1Us5EXEP2+EN0IcmIt95Nk3vX6XOj41BKLh6FeAbEJ7xX06wU9FUdmBMHRS+ZulvZvKPccwA27V+
psljFZsPfeCT7GKqEfRh6tjmqM2ysosRBhiDM/t5zigR71K2fZjqKPMjc73wxQas3bqhLNSJyRwK
qL3cB/Y/igRpbJGSbXhlno4WVat3OXa1Lx0RdWh1ZurAEKzwH3b/WXrbJgD7dDrV6DldIJyVg9de
LFP8nfL0sh2P8K84HGyMqe5uheVke8Nrct8c2FpQ0/gefvt7fIVJVp4UX+Qif5xUlfgka6h8Rnxq
PO9KStLH7yDXZKV4ujxvjs8C8A+w5j0OfC9hY2aJyJSXwurTQ3YM2+uhxfmpN5jSS40dbS+8wGqn
a8VSLf7/E0JSZZtQgYRDgwOiFpiBx5UeIWzYi2nEFRl/WQGi37tXkB9ARwomQBmt0wzRz+NyCCMR
ezQQeuyvjaOASwPTgqoEMzIGN3FMKUrKWAJNeAqaFJNa4N/GvztszqgmaLOrjFvRVvFaa9jAuSLO
XAeISIutLxIElOvlATsNC9cqO5pFSzxBxxFGgIJD1sroa0SDswnZsKPbUjOj0a5i35AwCI1JpsEt
rOXmda8htIBwJznWRViztqzT+s/qhz72i9Wik3TnpmQSH+z2Dffq4uBDKAUUdQZ/JDTsAQJEsCLG
qdFeEGUEYcXQWkn4jjUSJgSb938+aC8VyY5b7Cnvv+kEHj+MwKtIGkK2f/0AspGc+8bHJhi3mKZp
TidAqvaKo/9gnbA4UNSPJYB9318zUMsN87dkQSQUGmo60IMNG4sIsXwEvzS4c6e0BXJ5Jhg0lmSl
7oBvsYZBIdnMwoglTHTICo0W2TdphSicWHM6vp2BxiYp53ZhmJ1L+qmWtxzCIvaF5kDyNVjO3xdk
ICpk9H+MwKzdezCFK0jdYI9hSbfLFgePQs5TtQgzJsVSXfmfX+ToApy0DVKxPr+fgXNDxNiszjFZ
BHs1ZEhjASlcSa6EqJSzprH21o9sWSIE2J7gm1wW1onKIfCDoDKNGTcld2BcD0e80deqPV17n0PU
/oodNEcM5qCwWLY4jcxW1bUfjklYq4HzowudpxSdpsKOChtfj2LvKwCuu6Ifb3n/U80nUiz2cedB
hK7PBR5/LqZKBnkM+VQN8npUecqVm0fHL8AI+8CqH7UgTCjbuNOw/ZU0Azjf3qe+CRunO5/XWXbm
velxwnVLbFwU6mm1ho5CTeJSysTFw0REO5bcE+150jjjK4ikEbJ80Z9yMcb0IN3czH/e93pl9Bqw
eFfxNaqdWLRPx2rfn/2A5/AQ3qN/5z1ZD+YEdiYzAOYu68GR3vvWmhWHQDPOgxrfMKbmrBSvKQSo
T6ZfFfU78XBPxWS+rzYei8hg6eG5BGskcWV1IsokvkqbIMq9fAdzK3AXD0blotS/+eV/3e0fEYUY
qs3cSRq+C/z6gNgAYR3Ykg1GQ1ZiCCpTX2iaXuVpRaLVkhAJM+SxJgu2EnKS5s/ES6qG2AKaH0Wx
lwsKRK2LN8QGmxEvInXnyy42WBBGkSAeBWChBY0WrD9hBJYYay9rElg6OG2odMmych3rllzK32J5
+/Nyo2WUmV8Y5NMdV5Zkb8GZM0VCSo3ycOvWBqoac9qA97j5XTIBuxoUDbn75t8JDXBpRlYlHIPm
xYiUiB0SjagjFY9TlpOeYbrU8JWQInTb3lz8vtYtVJu9RZTbV9hPHY8xpQsVyH8kL8O626D9LzWW
ypNIEUijKoy6KIV4eVt2EhGcZ8oGTyBwlJaWwqlmvE7TWWlY1GFHfuurNuniQGqh7vkcQeOkJRlq
6oAHhbct+6pLneWb7uWWZ+gw7ZTk5RR53rEtFQ2XfKiKg4qYAS5PlFBNNkZJJuK8XD0ulqA01f/5
Zlsnaind+gDUTfcGvAEILIqnxvpk1oyl82l+gV6aGkmA2MAQroPUv8K42P7VFuU2Ur1OTKMsgKew
+1jgLuHVswXfS9bIfeQpl2P0WHulHIz53JXrHwHrfTqk6RPwl4Mnsd+/N/4sHFt6ITK6fzfeBzdO
h8ljY9VcQZAGUrNUFX/7A1NrUVr7e3r3FF+pjYzj8RXmnb/PXA3abVLs9+bma/j6su2gjsNQGflr
NpVL49zH9zO567uILfacsBRJQXayCd55mySZYK1nyEI9mRwwcSOehg/qTMbBU3kvfJF2VWd0txey
R1L3XWODau3rWzIS3pju1pMREa7KndaCSyR0Vyq83jIYoSA4RUopIwlY4e6d6SuSaRHeMtOQMSmK
TRqpGIepZJvQE/DK4bLB2nhYFNq4jHaJ3Fa6LopfvFhskL1LibQ+vYKnr6QaBfP3SrnJlCrshRcb
OIGsoEh8QZFx+PhPvOw8HKu3r0nUdQhbFXjMlBLqZ6igfMkcLuwgkC8lvCA1XPX/HaBRmRUgREZD
p4u8jlkwDXjNWTe4QNY1NQ4slIiqsXExXgbUaSc+tUV0XJoPm3HMn7yiPjEOX3UE0loTJQO7cYCP
d5rBP+krlBRok7Iyk7cDDZsnnr/GoDfUbNJv7xd1HFTWPQ2E8p0syNTQ9wX0haZYpVhQ5CQmHUes
fORJJoMiGLxsHfcSccy2a/BIm3xJy5Jg+UH399m93lDuqaBrL8MIBf5A07Kn8w6JBmHeF8nXlHfY
vJo1ne7WWGVM1EcjxISij2sY3/7Qfw92zmVNXo5IQbq/06h6iBaoKNnS/gDqJGVj3s2jiiwiLa5n
7S8MmxktmZsLpDoeaWKdu5iExhyS2QKRidKUlGTEWUSRWjUtL2SEE71p78Wy5D3XrmsSv518JxBY
fEznmNf6HH6YpQiaciALBtb/oE4f+L+IloDiwSzwQJEFKAU4zuyz0bTdiQ7SdoUDsEU6Av5ORhzn
DiOerFkqCNYLXy87SurlmXIoHp7JkGkSMEP8ISOIEigke58dXTAt1MMAAm56+koZAleyuiV9jKDe
1ArqPXCDP22smXZEWdKBSFtRHq7QB0ZYOh/C5OGr/sgBBTkTqySAU8yUwIxonNgtZ0uqaGkQljl7
ddyrbm3K1ktUur3iTCqP5PUqMZy0BW6SSfqX2BfIkDqH982lP+Qj+orU6j9oS4pwpug5Oh18UoLa
0VDedh+BEDmvDUs9EUmSEDAEI8fTZWVGEMLBQwIxtOzyKzBdN7v9+MQH7eyF9LyKnpahjjD0tEoP
kRPswx2yMAYLKJA7KdtCcQ/11m4bwdxGhBX7A6s6hVbYxOrXo1B9X+V1g/wuMjDjVrFZCHJsZdlN
uzUWQRA73cz0ovEOm29iTGTMwXg7pfrIhtHAJgVP/Z3+oe0dBcZPq/qO3QJJsZyPDS8j7yzTOKkB
0xvu8pxjYYqNN3Qatl473oq4f0Dm8MlmVTN0xd8CKmbbBObv+lqv1uZosfdianbXSElEJne2o2R3
5DooAD/jgoqzXG0BdLLhJJZHImDgJ3lwlcGA1IAC6Fe3YelXiXEit6Vqoxvy56MWBsn65HFahQ2o
yvLT0hu8ic/LnwlGVMuWHHjaCQUT6GFu0FKiD3AYBtmdFBXHbxzFpvja972dHEaPziCYqsRr4AeB
ZBIAJK+HdzA+Vyl+PbQG4NZK6YzHH7zJDDlXAIVMAGRBrjOBYMRMSEuDAJ+MnWOFv00nhyBWa2Gr
8dKbpTB5oJNvEieFzT2CSRZThGyE0JOErUwyCZwYalH9B66Wo1vP2sG0fAIhdHX48PMSCYq4q6hj
mv9DUDmzsH2jKUMY9WsNsUCFhIPAzbo7b5HdR9TJob89YmZ/lXu/oxtUVC/MLxKiB0B18q7PZigJ
MLjRMiUPaZsiRFGhVfw9tAGD2VVDNO6L8geLf+KBS4Zda0CKH3Q3/dpdF+HKzp+DrOjLfVZ4fvzo
F3joGQBaDYZ+1b1McPa8SnvBeSssp9nOcPmlDDcNlYnZk6Qwa8u8uPqyDHSI8vdN2353XJxrL3mX
I/vNckD2asxsylVLlC2FpoiC5dsL+bNI1j4KvaRUlkps+j7fGU7N9Orwa/cdYTEoB5wc4gJiBd63
eCepdZ0K4+8WeG2IuCAdZCcbMjJV1Zg0GZ5wLqlgD293RIDL1GN95c2t8UfuXLh4FXwzf7t9Zxz2
a+5weQl43L3Zvqdq24i/1XAAv+FqpEmLDBNeLz4aE72q3APgGcNihsXXYdgOe703dss+u4cGFgbn
5RAi+//ueaXYm9J1HSBSKm1DbFGUpuW5Kr7ymtuzyKYcIVsSd9Nk60fzJA9b4VPoQMdOQCqP7Xns
JeVFYYqE5f4LL/W/GO/PVTZoqRzWJFjpOjvQIZzcxjaMrYCij2iqEvKeZtH1K2+DKwn3cnew4eUD
uKTYS5+zvLKgiorC6waV4xwxP/XGa5oJrmpmwkBOY9dwp1QPpB8yIHK+8IWi6Md0P2EUN4OJXZuR
+IieechUIo4BZ+cCywmCyJjKcRpP+2WRABt0OvUTUJ3xYz1xYJyaig5GWGPg4BShEGYBReXNBfAQ
cOof2Emc9uhrAVWERJqlEjR4C57UvlIutMnOcrqSUizmoWS8XXDnPs37W0YiaMw/nrLocBjO3jpe
qKePTcI39VzlYy7kV+Rn6ikMinMm1DjHB6sFvsKi1mi5KYss3NBiscXU/FmYcpKoAzUnOdoRPknh
1SXhrvG7SNMl3C8fzQ9CVgssR4/IJHid6dsvChPOvnYL3qcx540J9LpDmEpfe78xTFqCuze35CGs
nG5e1n8wzn3q6RYocMdp5IWvalAeR3wIH96CDPIeZgaIUEK1hrq/Pe57LZiYCeYCBO5X2onzIS8h
6V5ugJwbmfB7rPkuZT4TM5ROZLdlmRIpY2DzxkToiQzST9K8tGGEUqPiPMn7vnD03ooFcj8ro/Cm
a11FCYbzskkoMNv6GQd2iCdthdsUw3bDRh4rEgw1mFba5JyfKw4vZ2XjrbBPSq+EZAIc8sIwMIpv
+Kr2yB3TSySXTi6aetO/ODv3d8iA6MV7uyd05meQxgP9fXSsbVn60v0bKwDTg13hvRM06IUsbQGE
q5tUQJ89SP7UrAO/T7EveE8xDk0MUXUEs6ASmruxg+V3rXopq/8D3iSP8fNYuRcaUa8nK1PuKAFY
PBzSQ6/uW6hOfyFz/sH4AmLiYg7jBQCTELplG+8p/xGj7v+Wl5JV3RPVIy7bEFSSwJu5IxGUZEKM
CgQBzi+gdnKmXcD8n/G7AUeahQLe03XtGGpV/GjWjLKQ2qrBDExnzjlsR4a5OfrdMWuyc2UPau7s
erC6DmCfFx0/+EWywOGnyvRSiDCI9F3zjryuPj9WhRF4ioQqsEQ/ZsU3gN5GHVC6k6ok+nfpzli9
0scmpY2WJp4hh2WnyX3ZK74GFaZY4QXgsbXPSuuEW60nsX+VRDbEGpMqLxgMtUSDZbwKjbbSeNvM
wOoPSIyfSdvvfpiWFfxBd+QpGZFc0FD+JLgpCYeHGt3KHo78COwOokJq6b5XQfLyx8/g6QOxNZKl
3bIzR47GkPWyQ6X9VNZKyLGNtRhvNurJqZAIX6wy5xSSVMtAL+LYWnYkx+TYCOiR2X1pguI4Uuny
i51POqh6wFPQNpX4qNH1896IIOFnMsgZ++ozbDJsxKy2hoDmEP+Ew1Tb//+SS9jDfsieEjd/jBwq
cz/oKRpZFpqshLrwFpJZmm0ehklpUPcKD3gJ9+HkBrCo787zwgveRHuqp7iU/3UJEjyucT8A5sYr
dwA3FODUOexx3ZwGFcatTGKDRqRXDh7m9P/EuU+LKtigU8F7txc787EnTqgTjZvZR/4+/+58t9dG
iR6NMc1o9dKrlzewntvcWvkmLWE2PZmuXvWwgKWRaffWW7HR1wqfGDt8Orbf5eqvf1GQFLrAYDhI
CnGTrECTZJYred1Ct7fGj23xxPsgVkVx/jpDscyUWh9qW8jFqfbdD6qZc0k47Zlja22zcEVEPulF
JgtlIIt90A4BgGUs230G6ZMBWzNKmUYqUFbHBbwvNkug9fJ2GdA0aYPZ/W4oHukcjaMy+BmJz9IG
/phUv52cc76E9D+EuFmABJ3eONo3xqcsLgrtLsqlWERj+EanJx6eJnmZa4YOH8NVMovr6568U2eH
ulprlRpeyzTqCNY9D0nCsF53smx7gN4VdS3h0xxePfblbEXtGokETsD/nZUgaJUezW2aEZA/CpxW
ltUtGGRmhSiTLJB+gbckrX9OoIPlc14k3tJrt2k2QpwLXM6IZTrSMUuEYgxqrp4Fm76x9eFcYY5W
JJjSh0/BcsywwDZ5p9+1qH7RqvqUvK4mmFAFeAkw3hfMc1Sx4xqnD/lcZ1igJntIL3fw0kSLed4v
crzcyta3MDzNwHG/IDa0sIQ9LpoFEELu1qtaCUXCtVPBhpAkzz7r821nBgXIiJ6Bfd7gnScVCzJm
Zt/oW4snoUGHc0C2H6WEayJrjd2Uy/LfBcQW328aojg94FlZaFZAzSYb5LDnS9TNnG4uVfcb3jk2
D5c0CalPD4ohcrIS12s6IxZ/iQpZ7p9ennMzNEBN8INAlOsRaGwkkqdZCLHdMuLdQkpBL1xTuKDm
T1LhShFvyS0h1Ddv2oaWrYt6WaQwpHWpjlbFeY+r9PvwSPWCdyj3k6KDJ+QG3Eh/bynXlKC3734V
2j+gRuUOjenlsbg3rCfF4WUSdSB61cSFHQ4ARraTfBSr4nGAvCElV78IPAnytTIKFHXITJrj4byF
oc94OiHNyptWp0TZZ6zJY1Jpxf1RvYp6SV63IGIaa2n8rf7RIbCOvx9j92WoHu/s8mF0McbIqSCM
XupQ+yMyVr/R7gKQlQIFT6CzZ1ZqC7m28ihdjOkpkcaDWpN/Q3tjh5Fuj5nE/c714940Inf2EvjR
kqBCzmbIyU0YZSG6hWBLNQUFckXrtmT45nQwhWaYYMKv6y/gI0X6bspzO2SlUwm4Lh0n5kuAVpMP
q6TTAhGYiQuWlWeWn/AUva4TEVCy/94BJuP0WxU3VC/TUI03+W1zB2m9K3QD1dZL4s85CEPQ8zKk
hxhg7yhUYEKhlKNamT4K27fetDDANu4O6GoU5PWDTviab4LtnY3Q8JCVyqvXgsJTLEU4BnUFNe0z
uGCE6pIveWr3KRl13GNN2NmdQA0Op1uLV562t4YtoN8xCibeljDF6wNRYhfU1Yoweov6wi2uaVzY
ZKVTRMkWTkTre1aRzDOdYS57v6h3tY3uuw2USR12vth8TinnepjDA/HaBKSoP+ts28H73D64+X12
8HUeyZmVWppdHsjeyMQDBivgZuGNbyNUsrjEOuyXSGCns8URhAx12IGguSM1rc0lnUfyVZoGKQ2B
AnVb3ogHhOX4M+9XyPaUVTJnfiuEpHeFg7XGTcEHBx/rwJ4eBDdg1/5kMgDM+FMUikaNHvO1gf/z
sxIgb95TSjqrsNX9qn5NT+qu/HgkhDZdIFVQKW2E/uDewGmjl4rYJqPUWp0hffseaOi2Vfichy3D
N3r/xqH6Eh/BMfgy2zxrPIHuwUmH1WnKao5eVGNnQ2NR1WfpYd1bCOAqRYysJXoXE7gRVP9cwD+8
1NWyQBuXc2taoOXT7o5Wg62SMMNJbOwy+jY0Eq5kV0oPWW2H3CfFy8I1DobTqwkhSKkhCaeE20y8
/kFM/6SJBNWV4Ce9E3W683N0zuyZQAnrRA+OAmA3vIRC0aB7UjUIfWpYZJrO715zB6FNXPSFTFuU
58nHs3ZezjlKwsZ1qTmCO+A3zNSfuDPt+tOJlRZWTqx937K1GJit44+V4+JoPqz9ug6zOeC3eJHT
U/jlC0DkStJejNT1ElYa9lLwGU6Ef/BMk787N9rXCh31nWrbHR3OlhJuKKZB84SsTnqehsTiHRVc
6xJ7fqgF9zENj1Kmcfb/+ijWdfOZ2vk9O1CK/CxP0caSG9FjkQmtPHfhPU9EtoX3n+ZYoOKtEMbZ
uZA9v14QWpVKRhJZ4faj5RWMu4KIh2agcfXaEjGPuUnAc0Whwoq+ezN4mSCSBKY9iHWFGFrvDKsL
2fCUKlpDEWr7BTnWT4i5z3b1hFXNAHDmX73yOlaOdV1skoEenNT70+ZabzX7PWP3KW02AkXbQtUI
Y0htsPwuAVqOVRM6ZxPHtAq5JzbOXY77fCndCJ35akaewYOsdnCObvwv3/FDVwb1PoBjMwjxHRYK
vtm9uPZNA9PSf2AHwacGgFF39C4f/J1dgPGFQtVyZ3NzcfQX/6jESlL11vUO8eevUT2l5anu88WT
Zt8N72BC1M9eeC/eK3RsmUaYVPqmffsE5jeR/1UXor1qwSU0XIZbIjfl80Ky0Iw2UA2NbK0y1zt8
j/1hDWgj/2Sh9brJXZ5qMx+ZAVoY8P7HM8JLZIAYPeUa4U7QVSm6yBWXf/BoJ/79g0uTXOS5pQbi
eTmEnfErcl9dTRJfNlbeqo3nPVIAtY3FVan+Ao09fpsYngn0HZszFgzMY9aKW9PRtTh9J4jnDg6E
6EqoXPj4RFSAObfp7OgBB6QGJ9HqcWz/YSHbwpO+KyJb1pYTfv+VnCblxubOLnDn6rhXNXKhYSbW
IgJ+UEB6tUQ5BbA27q5KzLC03VDVW1T00dD+4oNON9G5ElOe1UtM+cQMf7oWMQkeSuXk+N1NquLH
95ePEylDZxsxG8F6MPSDE1tKoaKFgiGR6wNJiAZmvfKryohJIaruODO+1sPpM6Lp2fRzmpMJpXYn
UA4DWJrXA9vnoJe2jVGzlDKSgfF5Zr0k9Syrc1KIS3I+mT0ZNYuVE7awlE4Mw+LLVjWUtm+5kRtD
VFtmAZIN+P4InKlTMltrmbem3j3svMapqRenpygpooLvoXJ5jEZ46HWYoo06CsyLlLomk5WACotD
Irn/Irm4W87vW4p9TJu3FSOAiE1eznKi1uCMB8oQmBoKizwMLNW0abuOWK6RpM0hKAc8oHh8OGRG
iWxqy5KSYaiPAQsBjcUJPt4G9k7xEq6E7PwGOATrgAgnsDpdd+yRwB35QgIC2Xijj4NV7QzCx3tD
anh+QxSnTiUzpA0/zXf0Tap4nmLFJcYH04h22SgTgovhQUWfNRznc18ZTeYl55mVDQjr2WHXh2dr
yleQIykrY1wN377Je7MZW0pNjMN6TmeB1UBcWimYL6X58ZgzcGjeFG1iNdca5PM7UJqQSOLBON/t
ywSPTPV+ncQ+34ZS+T/4lbLT7Rv/0ijJV7yI+gWz56Ziy+Lc9jqYwvjqaD/bW/jKyCUZHYgsAuuU
qF7AhIt6WToTm5Bv51GIBOXDRTlycITCosSVjj6UlLrMTRkSrv5FH8jv+42s5PbP1QF87HxIq2L1
wgVlczmh811Dprbyf1wbnjCPIw+h1GLWNy0llNxUy6c6Byac6yBEq1dKHUEFSlA/3o2KohfzmwIf
TJrrn7J6vwPWK7SVjLfQ7uIFHKmIpWV8u9eDRdn8oYTdY6iVKDQwB7GWwBm+sS+FTmwOihOkfXOt
Vpcxc9YWUs7s+aX4aAsEZIQWHXMd4oaSOCZiFFtmkl1S4I6AIk4tX4N42DFZwFPhLf9Mpp4BGSJB
6R8EsTw20cPZJI1qb16x1k1f+/ewpJiCsv7uPgo2s8WvnZyBubb4BosXojr39IpZ6rfy/g/5U92Y
trLgNMeSzKLApmoheTTeVdeu7rjwOx5ldiAjKZLWd/x0Yv2xLvws1OqHb3y4LYoLKXm4UvRTfHsS
shsEjd6S1u10lAmrFGlgj2cymizGLdbW0xbRmMdMXC0KyZqoXsXAc66eJVgN1mcepH/DypKX1OXZ
lfhSP9AYBqCMrSswjctp/vxvOCmGRVQi7AyR4EURHIczUd9hocKEZIncTrO0tA8Wjz4egljGPxeY
n3i1Trc+HS2fDOurrIfxzsUKNgUJ9KMbswfJgyNwvSfN6xKWP9FiOsHEu7X5kfk3ISHFCTgPziNm
V/b2HVxlCMcYYzxsYaxi1QexNna/E6DN6cDOzL9sKWczNal3/uXc5H3bh8UqktjH8ObywhJEQIib
BNAjFxogZz7mYrdTS7KhDbwsvM3kNBfxQS4RrMrNQAk9b+ABkydg2lBwC59aPonlG06TtZPaTDAs
mP9X1oWcuH+xYvkVlHVLVsX9EBPuocNKRVqNPm6VlnjZG3ap3rffjXVKdjdXMWYOJTO4zncHoF3z
Z5vLL/CCuRreBq5yJtUZ0feDOq6q1Z274kBhP8JoqQoR8B/IhGtBQwXWhDpJYrfdKlnrx2seTCoK
Uv62tHPHX20sIzramNP6Vo+jpNJxwXybfb2bpvw8LEnCICqkOp4dRCfhEMJ3Cy6RJjsvzwpHeCNf
6fHW8vKfVhub36k082TjbKldqH0Salu3m+u6z1S66g7iWm1N7PNAjNKp91W12LYgfuBgadZOhEPG
Nln6mpxFrdaJJuJ30d9X2LQUjz2WazE7T0zi0lb1l0mVxq/tWtwJEZtvzIBRKOinWbLJ1jmm+fQK
q9igCtFBl3+yaWBrE2V9seikZDaBtpCmT2gZJvRNSjlPL5viUz8YcZc3iLkUeFpGMQHziUa5QAJE
pTbQ9/fdqGHeDnh+5qyp5lh6M/7neciVnJXAjFGoRjhNwIvZ5S3dctiJuf0nP4hJ42SEuNEhFfIM
E+AFOoK1mmXZQmyVQ5C+osgwDQSXyL9utCO9iLN/dZ1HXqu+2LFHGIAMKSi1RCd30xyR1T7UZBiS
aLmITfBychWIck2S1Atfa+1s689926kALG5xiQpMbJOmhCfR2zzPZktf7JQe4EEr+7cxMe8//l0l
w94ZWQ/vLps0hQTl6zMvxZMlfLA/MMa7Ar5MPpWhBJ5jSGv2Z81+7p+/f56FziGzYT1DmKUwF+2O
jb233FsGtsBmM5kGaSPDRqVxsEeRpGl50abBT2v+R9yrLAfvQmLQnZ01rAqcJQdWlPu9tQLyOW16
Ozzz4gjCYaUMSOTdR36perJM5HHJvZs3m+OgPnHWMBtg/6eYhmbsVmAKVe7im3c9TlH0lYM3ch4o
XZyB1sWI64E3ku7om+Ujau/uPVbrd3kpjSR+/7OstMXVqMtUpGP9lqZuMMEh8/ay0WhMXNWZhDM4
NxSNs9+Crq0veEbmoXW4EoPCTBmWvpd/J9IGxQAZqsGpHSa4iJPEHpl73r1o44isHX4WH4HFywwq
/huGVIHY5/1mhypdA0BXkJZqaCC5Nyt30fEhvFew1tsr3oaO3whCHh63IuSGIxKuv3AmFZXwb/u3
C4kgJOHatDp1u922rutUOiUKuXjLvjGBHh95C64e1tgHNZPFVB1+yry1h3WprAGreKs069LnZq3y
SIGXskIqSEuDieNYOD8vk3E4ym/EAri8qBTdS/gi/jYOxjkpI2adOln57rcRPrm/RSDcyKGrmEZh
swMbO+ZK2ERUfJa4B2WXb7oOyWjJQGNp24q4DlcGlxNrUwOEnqUM/+pusL6b1I7cfnO6K8j6mK1c
xLrm0kgOcy4ADZlFJGFTcFfU8hsxTchlj5kuIZVSkR9xYdRt5a3Xk+Nh3RwGJkOsraJOXdCyEG4t
Ek+45yzLLpIV6lCfmR99YRHXA7y//AiMTMIBRUlbQiEhFwCqjItWBba0A8OslvDS+IQhTqY2GWKD
Jv2QOE8GvPKK1JumPJLffiz7MW5d9Mzskf0gVrfmRbyq+3L/4yOD5Cah7kiBQVjG+fLsZT2YwJRZ
Xh2cpMXw5rJkUsxBA9QBK5LBKJguYLOMoU0B4YAwQP/EygKp8akxPWl8cOCP2nrHqbqwaFzwCBeS
Db36G9jZsiOWDuVHA/pV9+4KRSVoCQkYghVxcNPUC9RJzkuvFX3sbsFpetxzL/g3FN2D6AynTfa3
vn/XyEXMoWvN60YvlILeSICJ4M1E0WyoMT8ZgosF614MzU6tFNlzqaophzqqBHh0VAfOKJNqoGvT
vHgnnyLjBKER7/1Ei4HbX4YX4cMLeG5OLcFzjLMDLKymivn6jkPTDiBfwrJqXVKFB/RNIUIY9XIe
wWceUwUbP9GYlUv7PnDhw/jieO93vajnBHChohp/Kh7yfUcpNu34SVMNi4pAJWP1Js3oz9tHIz2s
o+ZIOCHxTDvBTuy3DyRuG79dIAGriuq7qL0MIFPJQQalONpqOvBuKmzF49Tp2Gjb4P7YGv2v7Rda
HHM4LSfpIszmUHUAJFTOkygPDEXPmgzUyqMmGk+fMOcLyb3lWzox0E/DLo/EuZ8BNxHoLWoxlOGJ
ON+NLo5YLujbGGuSsPbbXix7lrEaFXB+sjnJ7stldeeiVfPKq8DcNsl8EHlL1mBPWHuDsDtczfm+
RFzjtVtfWXrSTvCayGYiAlz5ahgdj7oobaCA4heahcIPulLv9c9nu6J/72Nnw+GnMgWiKawAEyjG
d34vyPBWOimBidVCFxD+NMzHVqlsx5DET/XH3ouQ6t2nXqBAAuHVYoi3UortlJwB4clJYlBx0zEs
AsOIgoxD2qbYP2XcFKZhS0nju78L5bcmpAhO4SBx9DWXt4C9an5mNvFNt5jLMiPqlQHeHs7K1L+x
So6NFPNzgpiKcpbzmlGxVcspV+EjegwF0LsZ1U6Dkgaf1Nj4kZAq8eicS2XkiHwl47u/kFD2kceS
jnYxfXm93YsjfuMoRLOxq9rP+LpNvZX3LBwniNMdnfpSxdwyYHb5LmA7ozGIwFH3BF6/K/CXslVn
v3po/n+ZJ7XFurOCgOOImch/rwF9jOoJUaMKMPR9y/ePdsZQlxe+EUav49pwl9NInML9MPAX4BaC
XfWoOyAZ7YWumqe51fu5Nj6kG3MV6KAh8fkNrzZk+p6igHSYdN+eply3uXIU0ZX1AXqEHZmEuT+s
WI6VXyVWciAe64ODnMM3eZjFi2Y8AxbA2UodBo1+R+OoxvxcYOGkpQQ6wPUfGea5muIVeQ4oDHHj
AcLM4KDXE+aihKl4YM0nt6uT3Qcr+m0o9iQcL9+8mSzMU1+Qqecv0xeQEW9zU1UnSaizUfC0m4aT
U2IFrdLHxT6N5gkeVvdq5BxYucpwL97CiiBzfg2Hq1+blf5Fpf+RLQnCGhZKNiYJsBjHvLlT37SW
kQD34guy3+MJ7SiFFP++WemLNYUipWQtrQ9Np0koDPiPL4JRecamnEA+n1tvFGz0Olqvmy5srBix
V55UIx2CzwNBZveP2LE8CRH1IwhXUrchI3P1HOgnI1QlsxtFMKkNSC5wilDxWb4xnLv1gGkTt+XV
0O5y4xMHfiFGKnKfckWadMYkvrbzGR0vGnVI1xE2gRJ/oGSRzabazZR+RC/v5YSzs2owCpNz5uiS
AWPktl65Evkn72nBinERkYAk4yePirXHLMePHmaitjqz/pP+7RT36S7yVGOJHsuIoR+whwaqk1B3
F7gagwdBHNkdXAoQkGb4b1ioFXx03hcXQKMqP+EKtxwhHW5rxfqy7KMUMYsFp+8ThOmLz9d2pP/E
3O2Q7aBy4kNidXdQEnv8n/YZqCYLUBASMkmBlCWgb2DMuWiRjAWnHFnozg2PJBQisH4Y5phJ3B4g
ke/c5lf8Eq4tAMc814UE7YJgRF+dfCxkFKjPd3HmgVyRbxhwgNoGLI9B23k3uXsaMtaO7Hn+urmC
ZW4z+FYbs16TWq0Pbq/ihipRTRi6xHs7nY2sjRF+hEMzVIvhJpT91OhUaFZQJImux+florHgmpOc
4Cd5tEIjtz2PvNDJAokFBGYy5epGrQ284oRsKIdHmesN003i0xB3AfJgRiCsXx30In7OyybBG1nt
Lwf/pEV60sgRMSxL/oiIWJTlKoG/1gj6i6adeLBLKQ3TQzOTCCxLV9HejtH4Wx5hk30hm0++XV3M
8VkpIwzoX8Db6iLOSpkAh2oI+PHCUUXbpFJG5lxjtQ7oSIFENkP7fn0gQy4+kBUQyinti13xCj3+
caQQdS6sb1NXr9o8jC5Bav4fxjHmBml9rWUqoHM6UcJbOT0BHX/+j/SD/RfX9WQLIBD0oMGEllfi
lZvLTLin3A235xmrv8v03+XcjqtEdAhPlLdqtPXEtXaa1eyhW1xK2NTvMx2wqkbFHaKQdiILnYXx
vIB5ih9Tb8FVZeJK6CdSgLHBXmSuex08j3C6K4ixkdyy9ncZl07AZ2rK59uVDQmFwthOYD6AeFSL
ZXTc05tJKUeHpk5AerNTQ07cISwMT6D2Q6ACN//85pj9CfojONSJzp6nS7REOHWGYHNefkHoMCdS
SDu8kT++AyCCXi5Yl/Rw3LbcSUliYLz8opQnLW9zt3X16QBRL332u7KO+11olFAM5oFINY2bcPsA
uv7YpFLDS+KT94X9UHoNI9z92TUbxCOwJHSwIvbJdpwlDM01DqTBpaCJ7VU5v33FHZLLYOGkvpmx
u1yRG01AxI/9/TqH8sAW9PR0hSUro1SCX83Wc81WLgc52saVvunrMTk7quCwU0DrQLlizj7DUvCr
DbW8JO5MQXiHcjamZ3o7ACnHm2+S2khDfoUbmNU0bmIN+0AxyPqrb9A20CTuRkiBWKJ2rcOP5uPp
TzUA3EFfG0sqT+jFU47zXfNY6Vz/nVd3SOUGc719CFF2dYYjbwh07nNSSewRop2J/8f6gStN13yn
wmG8UrejuheveWZv1CUTHE5UDM2fS9CjB03L8gfhrx1XMTHKfQ+Qvz+GFdrK291FsR4GXvCIeZZZ
WW1EEV82kpq9JnNbskYnD2yyU1oVgcay9TQiQpd6DEHqkUv9fVYzSX3G7QMHhB/aSb168pziwgpN
76t9oCAIVBrnAB1+vOswwSujZHNScBbpIvFbunZwy/181rN35ylrxSblgAARLzjlBnEdcajizYx8
T3YNQlzz3nKrqNrTI1Myu3pWbz/uu7DkaIPf7PVM6GrbFTAut0ILZkMcjo/0Y/JM3xLC5/kXVa4k
H2Hun3zj8t2jEEOxATsamBWO634uNwfQGTjgJidqzOwYuhCPhrkZICzGVtOdtWA/Ir5CNcThy+qs
/fSTf3tUn0Hzu35X7BYOEWYXZOnROcK9OsrZ8oAzbZfk9BOhG99RISi22dFUW1OED5U6MnIGdwO+
BTTKGDodTU0pkXFoYBMr4rTkJ+1u3XnJZx4YM5sI1OUcqB5yfan8iKJ2E8dq/deRNkAuJ9slLA3C
RHrp2joyWa6OTfAH1Ps8crST3ZtPeeb2mIhSoEjLu/HuP2sOWLxUUXd7scok/rkmoc4NCvzKPGi7
TO0w3EA51wY+uEs2+c9RkddPM/EX14klxLG7wcH2un+gcy9ttB8uKUVC73nceOdCKVAotkCWZIq/
n7wk8cZcFh7r1479e/g3XZDwusk57CHRCongexLBIYF15rS/J9WNzinjOwsZaAx903NJDHDstYaM
f9lTtH6A5qo+FGdwgpLx0B+N/PF4APXqWphNoI43w74B5Rq6b8AQ9S0kFn+HeIe4DbugTTnklW8W
GnupBo2CRPQWwlYHWQYrhGQsNtMknDWlX8axAM/LgqwM4rbAABprcoPg7bmTroQVaUU8QSJRWUEW
53hkqcOwmzmh4rj6Vzw/MgE3YKbRjC2eNeSHb1n6X4+ALKz09P8X1KRnYFDdj9wroRwdmDpb5bfX
zlsF2UhEH8ihowEQAZ1wl47NSFET/RqAYd7hwvjOqbt0o4vNlWw+w1MFQgSgJ7BmH6U1Wr9Fn9WK
pWHdL4mJjtyPwVoI1DYIuflhfx0gQkOQqTilEBEnbUiVc4eyay9kP+YK5dLVb+HGRSkftySGeJsk
EB4iAYtvkuNHTnWAneZgXhmZmcr81DQtiab68vjwicHcB0ksOmv7gadn4pEX8MuSYWJbwFY/NMyc
kF3FOssXy69ERGncngO5rtBN1+hxRA06SUZxYwf+8r9epWXNes1dSkvUV3/3EqBLXF/8yKJQn/NF
JupGq8Lr4eph9z6pbiaoXOr8IhwS5BCsyhCxdY3eaLHped0gzxmOGSXer4xOPTqvp9FdleT/u6oq
2MwqD9mI96YN63l973xRBw5AcziQ/AKVA+vgjZ+Ze9o+Eonj0hofGSGg+lYm0yONmE2cq9/LH7aW
kHwPh3UCB1qwZM38IQe8wz7b7iBiQ5DeSHEkmjQNmmMKAu0rm9aCumLi9VyJFxJ4mgyEIhrdo7ah
gTt5Eg0Ok292lgj0nYcjD49kVFNIkH5AuvZk3lAQ4ZPjBShIOXywoq+WpU5VRIMZukxUnko3Rc04
JUx64FWQ1eBWXRk2BMxMXvlVvZVU5UU9eLsloVxZf5DKP6GEEkYD3yAYShpo60Pa0wxO5TAmCE5T
rS6dU75c7ru3ygdzAl0F1laNwmc4qDwC0SNMJFOFLMZJYn7r5UmT2IlGMd0LW8laVRM6rUsrjaRo
kGyRjdM6Q8Z/BGd6b6uAxeARtMP9SIO8Nh7ANtyaQSEw56pK6gSvC4NYDiiKAJy2I/+xwNronaUu
vsc4nS2YojVzzfc1XrAwEOSQtsaFt1G30ySd6vYLRWwzvC60X8KTIv7MUiIHM5OM1qBLxoBQu4nH
6q11uCD2pcKJhff3WKrEUkSQRBTqCD08+rVQFRhdt7Xc1c4rLnnkbejyNMExjt9pU2ydmdBzHMgk
12ScNG37BKSk3Z3JHnBAIuka1Zn4Z5OzrTGlsGtpkB+LmrWJk8iApir6TnM/6q4dO6wykTO0SCF5
wBibnYvxB8CD+p8zaYQqeYm1sBHLxJuR6fkW5YkWnk2JpzSR0ECLGELD9FwrnBokqcs810hq+Gym
P0KMjjHNsKReog3/6Fs4lVs7Gke6vuTjFvjrOhT08MyQtdClIiDNYbtUrj+heh9nO/UzUs+ZeEXJ
u2vb5aFh35IGmSgwVNAadi69R8lhuLdrJOTZNbUL00s3DYmhZkNEi0dDasLwaSWAQi89XVmuJwiM
fusMm7Z3pHGyPS32T5XM821CFalcRGxgjRXo6mMCqBUt5+FAd7yCbeFeDxQh4RGgZwWgUpb5YA28
Xq7Y0Iuk6mKITy7C0osuDd4PSyuc1ukj7L6fik8Z+fbT5t3o12KFl7CDwhT8AjBS7e5z82cuQFZ0
4fC8TCcL0UDyJ/JMNC4oPtmmqEj5imePWGKbsczD2PnDKpk8JWJNTvQLx9/TJvAY3r16Lr4TDf6p
mCKmwO5lpGsIGxu1wIjC+2We5RuNdJt1W8so2KNtb57r5QHr6Er9+quwMKCgJJiHxXRidBBin6+1
fTm7OliySiRPzmfbHj0Wj1qZGxLd3WX2epYJrZHoIrlE+hW18Smv0Z3D+bn/NuytlaP8xBW4GmQ0
Zd9rUhng98VSfRsNnoS7c5Ie8EHS3sFYbB7pqAL2TF9dCyrTjXUa9M+oHLCZzq66Wi7Ez+3YTSAp
gQQYqDTTY02YsJpimdJTmP15qbXD81FGRQ+qhpbqX8ckgop/Z9S38YZXQIcXZkAzn2c/uNkBbdcq
2wTMD5+dqmIprKKTe305cEpgwmP13T/waDBu1GPZzur97KXahZ/VDa/ErnHK7XFkc6e7pIA0FZS2
giFd2H0d7S/DRwZ4ueP8xvjem3bBhYjN42rS3scf/pi+3zzhzJVaflGuF0n98Bz3BmVgLIiTk26/
eS5s2zkVcV/3hz3fTDCh0ITi80wm7UiZSmcEkkVDcPQT6IwVYOf/g0Jp8zscTP3ueIN9A4Mqjc4/
DBaYDXTBs6EZHFBfRs8UDpzvIm8rvGMJofUihWoxZZQ8QrvqoHti01nHfSnvG/5Brp/JV1vHgRPC
Up9V360dusv8hBNac7fzrekPoUzSZgwszeZ/7YjA2SLG+K+VoSo95XLB4E70e5gD0dUZ200vciMv
DK+qLMrbTIc2AK2OJnfoVUF86PK5gQmrXi3sEpP0iruIiFMHdSuOm/byhK4dtCCeQ/kTQ6FPqfz9
z0hl8UL1cFA8+sFqNxCAJKTuCJje4GvOQ+KtdyqbQefwYxILloBYqx06x/L4szEZ5xZOvkmVnZMj
bcBoDJHne2QcRcVUrULV0clxR+JJ89qO9I7if3CaR+bkOwBnSO+DKp4N/mtpverjxKxOvBhCdrZE
sq5gUvodzNb+0BeiaI20ORYBQQKTL38iGHBwzjoJKMTPTfP/sJ+LMylGmC+cCrBPq6Mb3wzNqRwM
+75easT1cnAz7bW/r+bGkBW4OtN6kXt1NgavX1MvBO+q288ZNsJBgojMzO6v+jQTx+glWpA56gr3
kCuFeADnavPttrpos/1i7cC3K/XL6UKlJkkwUecGI+BDmpiv/DrEtmNEcJLpZMGOCvUPMJfRexOq
neNFdYGUu+Gkuziw9Le9WjDuI+KD/4w12FzomoFA7Q21ObGUlCgfJBGuDXNvrwhPyezh48XnpyFq
hqKTlJkf5R1FjJGZ0RCj5lSn53+gi7SgMMngPYbFQf8a8nNZPhXQlVCmD3SsBYMTOBHnf63r6hOc
gTCvgFgUosb7QNgTQAkzEKbKmPZQkU2BPa6Hdcb2ByiCJQx96I9I3rd3Y7N90Eu0YBZAgIFXgexx
75ag53TXItR8+SmH0clrMFafDSeILbQeZ6ijPOfA6bwS/703VfzE9+zGJcOt+iXJR3X81eOEg6j3
u0EJb16kLTIcJi/1jApTZ1pyQk5WUeP0sP7k4biOVu5VhhdYu6IlwcMWpAiauI99WpKOgNw6glz8
Jy4d6FDs+SZdX1hJSFmWcDHdsAzniWoWSW9XPZzTx6FGUSbvSCj40uaYZxFWqGidPeFmMbTI6Lbc
ATFSoAes3rijF8NL3bGTMRt/6C8f2S6cXaI05fWnn8h939xbJ/TelEoI1cQ41fha7YB7ArejMcm0
8i33bwVak1b84HPxlthRkhbHwKBJdQ4VfRLCzH9vNZAI9RyKoSiKGBZmfiHYFlE4s+3jJxQ27KHo
zrkhvaJkyHoexEC9FebVvdrIRSPNRWomN5prK4OUI0Amp1y1kdSfRgl0k1r+yBEDqglPsPYkXe/D
w+yxTOO1Sr+S3el/Y3qrfJj4dDNNZHzjvGrYW7pGT2jlOytUQHr/mztswk+8UCg9owSHpy1dSpfk
B735le5G3fTlkvdtOc3BtJR/c6cYmVTHDdKLcM48joYFJ8cDeej3wvtffhUkE/a0ewPegY0i0ZB+
zAxaH1S8d3otHBEsyK9F/OFmFmp5H547wuquzsmyXzkRdMPKSw4xxg9GS43wQQLkBFKwWpA9C2wK
pjek7WAfUidrbiF2aYab42+tkaax7IrQcFGBd6wydEU2aJKdrV2HLy3oDFr7jmYR0mrVoc1pZtbU
Dm50kUU5DwhJQCxA0RckbtuKZe2UY0oKxjRD2UMkuXa+jJMzJVOMEMP288EB1CJXH/Nz7v6Hs3Yi
iDuW+nE0h6ZWM3sZogDFfJIWgbhBm405gSh+wiFGsnyz7Ff9vX3G8KIAvfZM1E9ssUa7vKPyT5dx
fQXL1SaQG++YaXLM+pPPbhzF+YLqBr0xKA/V61lhU4vYtB2I4YpToxtaCp/u8YGSwaK9JX+HCeAf
mjDvWnRg9Dd/EcaJoi+LJgFdCCq/fKlBKE6ClQmVLb2vCvkZvSgmQwQ0ta7SMPbiecdplqWOkSvB
yltvxa1e0LiV3kSa27BRIxNUeEpIf6y7HbIBRVmS5LtMO8ksLgVXOtHVuJ61doRUDcE2+PuNvvTD
zgB56+q31KhTQb41xRmxEdf3p4v2vTvee7WCn/iN9C1m2PcFx8JDEIzCgbg8ZvHcLn1PAolF4Nlj
IKspKXTWavJGiYZumFEJDmMVvFNMbo8ArGIYHHfFBjDSYaoFcaZNow3YFw/YQG3GafikUFqoqgZb
tqtJD9G8BHpnld6/NZ4OD4PlVgGqCTSETLLIjoAdPp3pn6ZGdQCx/BuQPURQPK2FxxuxUb0Do2zr
mcesLhhXomiQNPc5HrJAmt7KDob1otgWPpzk9eTzBa5ds81HQ3DWJecpyUcNTZR5ejajGUz5+r8L
wfQd+nynqgRmRhnPxM+Ope5loyJ8G5en2siuG+c0Bs9cz6EF+NXDo+MFabwrr2yZbwtJQxe5RDHU
U53ZEDNrxAVEoZE6H61xgvs2mttmp8WLs6+auyymruZ2iJE+m/buc4rCwCg91Bd5Qk56fSHnTNYZ
UKYDbaOhI3ugLAFPaI3xs6sYw4zTmMKzpAPhAVB1vkcC5a9juDHo/HwdWe83KIqiegJf62SuenhJ
Q1E2BC2BKrYTevnjhnC4nBpMD5KD4/w0QcpyrXnnp0OJaBUYS2PVS72wN6hpD6Ksz1L31FYUufoB
rmICboLcqf+LG4wKKjgQPQajACyVzZVrY8kgPmwQXsvDaK0HiMQlupq4uBaBQtxR2F8CFbprjMAy
lJPmmBnG9CyQfBwe0cADxHfFnJT5Erpsm44HOVsJeZTN79rntBwwWuq/Tc034hPtSB4JqGRivOgQ
YOjk0PGHyz7n892Ap9FAZtsrOgpH5hkp1qRsGlwjN95gXB1jzWrFhGmDJeWJTot1BmoAbG6EhF4J
IO4Aj7NgK+XiOl/zzhf3nW8qo8ujW+k5pRQFuuc2EEmBtWc6HYSnwSvVjkUuL9Ki/YPuqnRMHt44
3q3KBuhXtzDpUuhTzBjghbicjOun8t3GtQwBxKh+jcwBQ8UJNLu0vfjzBrZWyaply26fAuyCwiQd
ti2E53pnLqApci9X1qDwM5ZtXQu8xxCRqU5ki85kbvU2R4CKvdoAj25thL0w5HkPl6l+UwOOmc/p
ikC8qTTorTXwvQ21KQ/QkqnsRP3tYqUgDDNIEKHlhtBMn/zTTOviymU+iauLmA3R9UDWL73O8l6Y
J0vHBLbbSzxQ2euiXBMcVYEsrn9MhGct8Q+3+wJsiNpK2tb2zhWSqZ8nYvRavRnfj21myH7/uH55
dO1UwuhraN8Uksg5GpEG79Ylv5v8SNOKDU3pPirg55N5EuDIBpSdJBBQlsMToMxKQ1Z6soM8iDCH
CeOi8xcjMSxF8/+Iqqhs6CJ21bwjbdvUJikvv2KtNAY0ZQ/WjpE/0HQv3R86IKBEvdiGRsomI/+U
dka1AYprmismBsvSQ0rNKZ/zumX35PqaXS25c3gRxL83vDxBeserPbXyyUgL5qmIdVgFIcVbZCPF
WYUSNW35G0OI/LXloG7ZLerQ1dwRm/sbpzA7UHWHdHEqo+6eZZz1YL+Gvcoe6RYEFHzjyUJd4pk4
pD4TJaZlI3hOkrqFHtenoumJegJlLCoR20lfdnf/7jFK+d8tBRcnSZe1h+NZ/8FZ/1cq4GjCj7vP
kpog13L/CRGqzNc9QHzBSsnMxD3ABYMX+mBXjoaJMPhbZYqb7WVyHsUVQ3R7bnR1UzSuukn2KxVj
MflCLP2o2Fyji2ZjgRvfCrsXXg1hdZnMlQK18Mv04q3MHhietnzYxq2n92iStzgUPoVIiKHVSOJV
xI8RWqseyreC3tl/awYaywNwQk7X0WhrNTgiOux3zz4i94pJTdkwHJ693uPc72Sd84hBxVsTPfFI
yt9RKfDiTQI7yPhLElWYCEsKvZK984iA0MCjW5ZCKGltiuAgqIkT11RbDwzqxwaKn7nitB0i8K6K
RMSqpEJ+TtwvYX2Yc4w8XCWeaIKA8nemutM7NE5bn4pd4/8++QDEyeYtJkBwY5BD8666e/iqpiLQ
CRt7TLVjkKWLX1j8uLdpozd48zPv4+EArNgjBN4VfnXt1QTIyl9y7vyi4pQhkqPMZS6SqqcWyKWh
bLaDzd5EpFKZsLYLB4n9Deg/sN+MbuGTw0Zip/q/qLlqU+FqnMXDQifOAHoEzMaw0vKDcut6QY6K
6bbW77mtGj3fvGsb1+lsHjTjDGhQnHLpP2m1wLolzF3Q7rANAhj9ikYHFxOVhIXacCWECNEVpG/D
x6U2DGZ91ssq2QI87aMnV/heZLdPIC2kDzWPHHuteWiPxFIggADVKHXFxydEkTV23TtN5hWWjUHI
689oGk4GgYbVVCNRsTK8R7XRdCZwlw02QLjdl+o3cPneS3vDbJaO2HFgf5qeX+h6ezW0DHt4HNkt
wRRg1C9IYDKpK2MD52gGfPzMM/t8zlpJRIZkO4g8NQ5vQGniYWCy0Uy9lJGenufPkqoTxlyzpcA3
AkQxARfeIrc1FtwXkiVSZDP31QohU2NE6HiMGe9wcGh9t1fItYHQXnCOZbjpI+L/39MxfknZiBwX
LjSZi0g6SiHMqT1L1pbNntB5+DAy4SCh1jYI663XwTI8ZMsop2ePmBkYrBTF45JrkYvAUoOHRraL
4J2PwWN78O7N0gjKjw0LHROD5xVwZhCYns0hoOPumUluWdPWusS/uji/57x4bCzTo8FpgkCbabmb
9t9vp0Qv5ubo5riBxEQ6QVMrk54WWfFKLaZ21PIHvrzRrHBePZ3FDEnEDqdUKWqmmsB+Tw/mBaMY
dZzhiVj6I4L/jUdFQwx6GB5zbgE1+IVXlA7RnOORpQY4Tx5ie9hGMdAf1g39neilJomZ18GT8xhU
L2S3QosgboO5NMzv9th2+L+aYvHUcy7PmEOFSQBcrHcOKA49Ua0JtRqXzn+wp8602u2tS9NVnbGR
8ihFQTYwQBanfmiwN/ocgcfoIaR+g6EXvY7silaa4TEn0w6h6yXzzh6dyKYEmhbQGSNLtDz68EDk
SQa1jR2FQ5HkYH3JkRD/16tftOzbddbEQNEbagathbNl1LgDa4cxwR85TA3+0uyCIboieHhT+8Hp
ykBOQ/0Pb/m141KQO721SRTayrG2Ek/l+JDw5GiC8GLa7hpxp4VYaEHZ3hecw3EOgrkBHMpUnF0u
t0my2j8qFdBlT4ofUf+dB4iYuGqMOuWHhF42ymrQKyf6Chc9HhYuCzs6WeKNC+PPMaamPGVHxoSU
g2twt1QLrBZ73Vcbh024fNVsRjQqGkLWKbszjde3PEYcARBqNh7DsMcpdsVtdVn7VMG51nCCmtoC
PfDd8jNNA32AGz8lhKuyu9jwfcAhFQvvtkqK/Hy/VmfptIP/+LP4Gh7Y1M6l1wtOS1ER/2xD5Li9
RC9k992BIPMaSjBCle1sMHFsSAf1/aynoj9JdtosA4wwCRkqrSaUFwmSfJniv22Sjp4u8Dy3tIrQ
2lKBJUz8yP2IN1czBGjPZXr7gccB4bOYxoQx/3+eTGZJiMZJstciXb4SFpzx60yv8hH23JmO9dHm
tGQFdS1mxg0NpsjbKvA3SbYhU3NtZEg4WZpRRzHuMWsEEG+PtTgHBsp+Y5GYAbDDT44T/3wD3qIX
tG7PtXMvV2s4/xcUrvYh6ItTdbM+ZLsfzs73Us/5MhS+4dm2g24LpMg1JDi3OEu1K3jtrSfapHAO
qf5yVq+YYJmw2Sy51Ivpzi/jkkltnpdl9bciz6e8MsD/ei1A7QcUk8kB9lVqmCachE374mXqRskt
yVgme7kBb88ANJq4Gxn90C/sC/gm0M00Ogl7KXvbkiMOUZ2oIJJ4gXGcCWWieqyTogiHwjwHD0Ap
1XGiKPU6JRT15xjJozEgTBvvuwJbrSHB1wlnoKXmrlfKT75aZYYCSlQlkSnduRKvkx6ikrlfOWJz
mYUjtf7DpGYFI3dqtvT1jcP61DGZUPrd9ktI57LMJygppWtNSAVhTLYAI97FhXOfp4hgZgyGskYo
LWNkomSmJfLB+5xyrsse8JLBa/0ATn+McE1r3vQKgPntwJ7InUpDSZjN1K5MqoxRoCiMxhpU3MpI
c9MPnlFrIKa1lwlme3waoxhOnQCOeJTy24JO5yHa+LPqpNUwUNHsNrjNH0JplYCZTOaAvV+KV44V
kNLK9aYx5FJ52Uq+Y5QYMqIYMNf1mYgVu2ZbtAals3KBoXBHwLFjfNfDCnmOTbayKU+nsDDIW19W
mwRBEt7RGBr4e8DD8zWM2UuyxUT/ng8rLDumYm/Xadqru3eAVuSdl0DM1Q4mdqkS9GlJXG77X7Jt
nmERF647PZv8b8fNneWur+mXBaQM8Sva6dNn/rO13rVuWlvhY7cJj2N6sCihi/xds3FpyX1Y32H3
vzOtlWhYO+KZ7+kWpQrpHt0XD6NmohyAubm9Z4ByAV2ogWlYC1KXZAlE7gaRd83vnVltSaTF9zxU
6stg0Aikdth21YtrKkMozwVkGgkMBSNJ6PiJbl4B16cD/fV1+0afgEhLkmoqKqrwSH+VZ3X+U2MP
OvZVX95UlNSlkhKmkG7fJdpIAxKAX4tYSJtS+iMjQcu9D9RgWPX6e5eCJan+ErbwcMkTj5Xbaudi
r5EpT8XXyuGBgWzULpDwRhtxoMxKNpK9LJcSrRdgds4KyXRkaUdkzgV4JAJu0CJ40iNwGrFitjgS
9qqurKcgNvfn/ZaPyonU3x6XKMP9uJrZNK4Mz5CxqeuLgwC7rB5D1m/LuKxo8AUe0o6qC7m9fLEs
OoPOlx7dKIpYaJl2Aq+wAA8xQvsY4HLJJGfCSd3uF2FCu8pGFYAWkBM8m8w5bWxeu20+Z/4j1lti
r3B14HLY2XeHsfF+gfJM8iU7ZnHj5I54dc5YIkcmXXkHM8GPycbOM49djhMFwanLpvt4osW6im2n
NrHOhsZ3e9JUpDfT9mZdZ0OfHCX4g2PxhTeJBHVcZSfLDzJ0PjnZGqjGfaMw6ZpwjeAo/XoSfhsh
v143vZ00V+SvPY8pbCVFNuot/zT0SUR6T4dQN57Ep+fYhEloonpwF4jzA+lSQKNf+WhQl8wsMaUI
irEohRAWqmSzS/EW40T9V1uT4y8OP5+nIDo3vZ6iyyGl5gnbdN1aLHYsRMTb1gxndZbngsnsIIYz
ka/eQcwH54MUPo91lSZsBa5vOj+nKN9BBvsAQZf4XQ46DN0CNhIM9DChWENgpOoPMgSHj0tYLtyH
doQJ6JEW9uO7T49rE0JsCur4irCjkd5PlC0wS7nAPiiJrkHhbUER1qcMUy5nX5YliIqKHJtLGDRx
I6sT42KfhLQShtls1HDgLofk8ULdpmYGxfux32ts68YVJjcirvORdxy7z2FGaD52jQ/uey0V9rgn
8Y0/ArExN9xTgU3AdXb/no9Ue/n9QrdLacNIXQZODrqJItLF94Jp1KZbJpCz0z8Bw9THswWRsH2G
L/3Flfw1XJP2aS3RQglNuDhI3FxiP/7tHwCOXEK4eOJQ1No57uLxTFkT7QVQl0sGBuNaWJkH4NXi
k1DKnswZRped4UTcQ0cCY2ycJCmPPdL7R2C79ZM89aVx0vGEV1wdhkbw0hgyfHk8tgo27giKtbbE
t9mvzhQKrCgwAykgXkheIrbvoiBdhTc7YYp/BbZpoP2EP5blxpv78ku7HDmg68sRI8MUDhFkL4dE
bUiZMbBMoW403qw5fStUYEXc+XSG0l2MBvPaeLVchlJDGGC0W8ZH+opF7wVJUce6DdyPlS9SjCBM
TqDYYfUqWJGvbJaOQHjMfcGIxK1phC6T7kuM30YYO9g/6/7WzIY2VBZiul0QAv6T+v1R/vO6IStX
efHGOQNHCKWLMlvtfxf/31sXAwxdzqytQN7wX5xfoXoab6KNH9GZkOT6O3GzFG1yhWl+9VH/CxpB
P7LYq2gVxlNnFEwypgPcWBNCbG7HrGzetlDGhEfWf5VuOgwK7YriS/j0FdYjROUbiq8a9IJrtrt6
VfCe1b09iL2vKFD9Hbq1aYBRZrsmdDMRnNs4SAKKl/wKtKHgEbCiawfj0U1HV4FuS1XCrrzavTSj
D3kIPKY3izPklli0eDbacgbBQeUjC7BY/4tWpXUR4s/JqgyBYisT+B2D7/miUwZ/aEB5fkd1owxJ
xyfWWCrqHl+A/SHjo7GC3RnL73dcyZrGWLRLDZZj2cLm8i5A5N9ZR6tslzc5Hbd4rJax/jpQN67+
KRlnRvJd/3rdq/TZZiXAGQyDVcRqZ/GeJc7mFNy11Dy5ce1mIFHkjtnN3Mk3eAbMj9xr89k0zQii
qOynzUXJCBGsZEs8DhHD5o2QBK9EKul8Mm6C8XVsCcHXl+ogBQwUXP2YPEJyOVO4uVkQMUv8oaoQ
ykbp1rLj+y9a4Hc1Pz/NomOgKAefV7G5OnKV3R4DogltKmxjstvl2WFmuWITBZ5Ne93WiLksq9Z/
o5qG5eD9GpAuiHEqRYHrjiRloFOL9WLqjEvSuBcjIl3Qr3cEvY5iryt/x8s8LAleVAwwTekzlPtG
gewYBLAq5kVaDUu/6EsgvuTzoT8HPLKJgUQ3njNQ1EJIG7VTc7uA0dvoAKfZfL0C/Mt+rKloocVj
cttr6uc5K0UDHPC+V1JZbQS8EHF0u8M9r2Il5NCGiRo0Vh2tipFumGHcfohrKEq3OFSR+7C4sJ6I
FDDnz/cZgQ7N7Dek3Z94+KNO0hDezaevaEdzEUUTbMI0kCIJbP6L7CLR497nOCiYkCK8QT3Mey53
nhbiLeW12wxQbdEHJXPzGFdgVBslxW5AxopF7XJ+hHpuOlmCLcURVWIUgalWO4HNPmj5dkCTsSBn
UPSZcDoDANks5VlaTXxPoal5Bv1Jt7s2yzdaUmp+sBD3kHncDdzodGcFPMsag9x3yRmnqxbG0L/s
wwjeoonTqOBD/jdgR6aL7RWuBkn0BOyS5jCiZ4pR3Qj60wEcwO/NL3cPnAxXLppS4OIaNbHfPn0P
gUpaievYBYkTwEe/5HX6W191ZEKXIAHgEodAyPVZvQvRAjZkH+m4iUQABcnBNw3GY3kUcP1sz8zI
oNnRXVmjJlDIJtuvvQMoVmSjy7pqwqrCVqqpX7z8dsHcs9lMomjDn7usX9WsnBXgKh6l4fsGH/PO
/RgFs0/4SjTgaTNaMhQIx0P2eEqaijb07xYizBSPCl7obLJnvjvg8ya2t+GOcbUkI7lMj6xm6b2/
Mfx54brf9Ap+eTfp4ydgFAXhc6dvLPB4dum9DrP8XyZXwmfKDP45Nin13aOapHuocT/q+VQFQnOA
jBhXyFAUBODcpTsjIpPqAZ4WB1LQVlmaGSU+t1N8th9HqgvGs1rTnvSP5nYcxhZd9pmB9ImISN84
sn7ejHAOD5+w1Ei45bOQ1kCX2Kid3Xf0SstJuQS9EGAbFtwo2T+aGDxBtOC58b0HL26nz2FO3afm
faMrX6ev/WNmPB4IVdX+CkknXOmbW1w1yi2A8Sr9ZcdzK5enyOnmRBIcdgMCTL2q13l6BsZtbX/Y
Omt82lQLE1lL2XMr3HhWVAWKcF3OZMKG52wqDTNuWLsY0hm1WMO3PC54iQKNLEv/U+9hBDcs5mNQ
SpXRv9avtnTy2B/tM/LADEgpg8QGMYS6rJemRdJNiqDFyTWk82XKKj1Ue/viyKsI3cRuCrSEM5M1
PeRTeklKX9yyWH6FZNHdDHdfpOrM8Cz3RIEvPFLaK76KbBgWsmihmBiYCn2B0DcdtpthhiIZgYUg
uN8xh80LuvDvQeioGQLapAfySwyvNsr+0vixYdkRvsE6vPzYB2aAe3YtduOtspczoMZjh3xfhOPk
iJRkhIt0ZwZLRBrx4TrfIjW6HCX1iz2FNQSVlJ/yH5ROrjGV7jAGBbd6iTG2TKAt4VMKtO9ePMbA
n1BY9uVmSsZSBSXWu593DN9bTd8AJ5LQgKpY+GzplKD1UbeVKtV0c9gjNQEkYTXYmD0WI1F0aUS+
3V7DsLgmHrqJrwWoP1wlGtLka3KK28k3HrU/0jagX2IVsJ+l3zbgY0j3FxyRBHlj+M1QNPRmSWln
Qldrc1f2wFtyZnQ3TWOzPve0ERCk2FiMix+zX8vncjgeiWKOXDL+Gjo8brwHPvjqexNaHzIqsPN6
KFoh+kZiHDCwk/XlleTTqvKkghorfhBV1hVVUeXEwDhM+oP6aIaJArgw4Vu7yWntVb5NnIx2zvhP
9qxfIQgADMYw7ENTDjt2Magc6VvhPjKZUwBKqQ/EtBTLhIaHk8l8caNui2S4IXDPLuqhdodFGPzo
RsBTYmH1RVoSnndA3jGz0bY6ncw3GNGv+HGYp5QO3GlI2zgg1JQ7aS9h0rgTBUo9p7crdjGHWmTW
0TGnckq6lUxCgM9PyR7WQkvenL7g2VpV6UsBDdc5XEpqnjoLqX2RQl+P2EQEcP8bkBV0giS2i3lg
V4ZXixbRtlhW28+QyPqxZnqFhrQbHs/d4rZW1X+kfK510MyYYp5WV2QvO1t5ZPKlOQVc6/k7iSDe
1YjVpYieVz4Egt7nk4AfDkHIqhXxg3eP7qxqc098MYlaD845Q1u7AgC24Xn+3vwoB6CgsQoJXH3J
eVdts3Of6fihRKZCwlRuaJAmMuOLRWKaXWpMixZuAxaGAJ0XgAKdAKVmuYDKdYDW5ypzhnh5Hr1y
1oeT/z6/ik2XucsNMBNlvaXh9PFrQujV21peIZONn9R4F/TSIV8oyfknUEX5F/npRmVHO2b0+2+Q
rXJt/ZqGab8a0foThhG4D4vzLenbJbztDZ86+btKkNCgVvAjeAuqCc1YjU2HIvUQpnB4cgj8h5PY
hvgcyhYZK9MDPC4HSNQ/QNcnqheDvtpQLrrKg82GvCGV+YPSYnLYFMITuuS5tPmlm4JNbix7Iw2t
aydngmpj5q2AWls/+eNmJT8QMLJENpen4cBug5slwpbCwIzgH4vjTzrT5MpIr6oyU/tdMyNHoJCw
vbmAB+H37ELjIhrmOvQGAsAwSGdavPZSclrP2IKNJU3eTcmaLGZsY8JKBIXJE5VyFS7HBRVO+E2Z
nAsIQ0TchorjW2yHHqayR325jDnF51Asc5+vJ0zJGIZR0+C7fNjgw9RFpLwfjCan4/OVfVqCMpO4
7HzVzVUp5gE4H4TfBPbPrA2ZhxtF5XPk0sOK7WA4bZoFdALuvMdJlOKwauNF2n1EWD6lN6CM+GIh
vy8aqHfd0DnPEy+/LYKMCW6kKVekRiMnUGKqW+pxVZ8yDIZd9ECKecZpOzsiFcfrCRj52PL26OEl
yjz0kFjENUEKOj0QJoNeRxRwMK6v/vMCAhmHzY6hU19NWNnK/WkhY5dWnLom/WAGM0EgUArXDh/P
+ECqkffXkD8jW7azsiipHkZsG9yRntSwzbPPUBxIGavSUyCE2mt0hYT8s7tGEra69/2s6EKeVld5
r7AT4w6daI2enhoAfweOGj7BjsulaNXyHMy+zVivaSRF1qtBGHxZTsWgYkJFlwxemLmWALike0nZ
zmz9dUNkGyy+FqeZsgr/pb++K795WhbfFRg5lwewdW54OE6h6v08Zgp+eZMys2OndqoLZs65erCg
kmsQ/w6uuBKuRbtijHPRV3QvQRCiwIUoRu2UXeuyVlUPOWL3vJzVqCUZlk0MFIXkB5pfr1DZ5was
JbGx2g4iF/+p+s3sHv+FoUqB1Xq/iZGp3qFOWiuhEACpPd9iaT8Pzy0uwB87ti0CgWEgOEzaLgfR
+B3ZlNlTholOob9YbrURQwLpcygy6IU23P1EmKW4kjuJreuZuC8CNKzMO3XlFn4rbGfup+JBPz+f
mc7I6AzmPhfKUfxU6NHyRVtocp5rLCgj+Nge3rVbQChblbStD7uHylUd3kABQD0Ww6CTktwnFZ9N
7MujRUDjw/erndI042Tla8dE2X9GpbgUBXnNILepouQbHvgqnHYAA7UrWX6KqLnBxN5FIn87YxIY
0R6TSAlokjfeNdmHZEUKOo/oG6AzOY97lKboQSf0//P5AcXi5ZDR+wf6cP3TMVhg+NuEJumggjDh
miDagaCLyFtwjjYLT+oJJUZvjWUTC+vMq6dOPmONxHLG0CWj3K7RqfXMPedHigTKoZ51CogB166X
L3GiKbC8e+d5jxc2FiePpWeakhUWOjKHclM3ZCGAKl0j8vw5x6iq09Auujc+t+aMNN6Rf4o86+zA
9s+tNyeCYMPodSKk2krfKtFnPkNup4gvto5P6TFaAvrw8aMUF2hThWJa7uACUayvKMf6slqRt/aW
XGwpK36F3afExRtA8abv26QFoDcKhuiKb40nDBmnD+n0vWHxxcN4TKF1/T++oP8a0JEXMt89Braj
nPdqzVF/85hmPXlZJ2muLZD5bW0jZKre2GQ1A4YAoqKclLjJl50J7AFZAAZZd8XDZPPBAPRwh6cA
RWG9AIco3YFxhJ36pb41cD4hVfhSBk/HJ5iAk64jxksjg9RW927YnrfAUegdjjhZjRxgzJ0OOoVk
eDN1dR0jQeznvImQa4hFYBbYpGPynubKtQlkmD/pMyyM6ourQ1x/jPYd/NGp9/Cd49Wlx4CVoH2y
SWTuKZeYBO9+GkiWaUZtq+l6SPAKmZ/KvjbssOdpaId6YHLCk6kQhfWV8bW6vggdFv3AlgcuKjzE
fd3hmKcTKk+ysHoH1S0A8N4pwKoKnd+mblwxgejBpxeSqYDCsd3zv7+LAVw4sNh4U+PR1cxqBGaN
mgQprPAOKvkDYIxLYwL2Gn/t6ofjeak3j4qPMy5K8z0FfdUVpVoErzzIDC8kYEAaeLJNhRaKxGZe
+MoJGUP4EpiKU7fQC753WD27ygPB0lgQxXEODl1qHHRWFO5i5uA6DuxinDj43nae8vpXB1Hk/4Do
JKN2KvWhYh9Uum+pghGDAqX7lzOozk0mhcKJqnRXmefiGMBeFxTAIn1M5IzY6jg99YR9Mzq87+oy
LmCV+1p8aKOpa75C9hvevosl4Y0v3s8ztm8czm1UgUFGYUkc5RQelHERmD3XlF2u2z3hsrxdxz37
ooAubPO3TBAK7WBkHgefUbDEBQoS1z3hF4irG4kDnqfT5Cus0LpXUk8KHoj0PWK7m65kuG209JYh
MphS7Xv4JAvGVh9YpULkPtTkvP9ZwdhXwyfAsRUKnf51kt3HsH0wme/CEjMSFBOCQL9lV/crMsxi
4/RYoKFXfUkHuIwi7hwMyhsgiA9IVRVvL/nCLe59OcJtkPRNdTD6u7PKgyyvCw1slcbVsw827QFg
nVrUkimduseYiPAfXRPFPqu1BaFXWN0PA5hkMiOoPDHpNB1YUhIJ4dOkiW06sHDMg2KENqm4FGVQ
EkS7+KavUntbqAPMGNENcmnGGIx3cTyFQ2tGTPWOezWm/GipE8KZavgSwzgwvZtt3EEaeK+54HDT
Mrj/vlLgPI8BbHiavrFfoxhMm/kGGVZzM8X8F3zAWh0rSwvfLTjO9LeQir3lDUoyempB6mMGprw1
LZIRXTv/Ke0Cu5rKb3gAD3GeSFbzMGht2U+dW/3xdRwFWWIT5awhVXkwqGFi/Lf7bk8uEXRY6Hpu
L/X2GWwEUXgyJEy+G9VZ53adVGZam2gjT6/zMjZTvhOvQyuYLrJO1i5JhSADtHTNJV0vXi92Ma2A
xdsTLsZC3xtdwBQ3B5mT2IMXqlb0TL1iakZbx/cSjxbdiXgf8zuIIpfi0ubiSmYwgGaGV9x4PyHa
e1cNBrp58pyNnbaHG+tH/+K+fbMYrwi30eKeQBIe0Tr9bfzYcXJwZMG+yWA/iM+6MfAvBH7KLxP/
MO+jC9aus/j0Q+HpsuK/uok4VRIDd0x69C7t2ZsjJyh+xzVgMR9iCysy9dhHRpvIUcEeY3VNys7S
w4V8nhyiN3pzfVcuWlYsuubwDnA13rDup/j9RNO/yGYxhWVQRl0pA987oUnlwXKbrevH1c4b/GAr
z4UZy0Ut77lPhvMvdxgRzQ2frNWq67YLHLv+AT8HJgy1kMDWeD6Z7v7M1p24oGNX23SJKXYflgA4
aFSu/5n9AOFtsd2r2wkYHyTO0QO+TXMWFlYzJTGPzG9B7vB6bPDEO1lY7nbi5X0ATUT61c+VcNNI
co6qfEgwqHND96YoxMzOpxqMEJlovNWfDGq3j7l3oqpSWnzP52koMoIuQSRVPbjRPBTQJssLxluj
rLqH+EJfP5GEY+anhCZBZEM1SIepiqmerJ2/eu87DL7yqsPjV92FFw5Ain+CfWcLaHaGWkJzTFnU
GOHpmJLVVfgs/zxFbR7LRfNKMBSs0pzP5sUADKjdVQd78KHcktisNbH7FpHsYer+BAhASVtJnjuF
bLHfLFNf8DLdFPlfMlYKaBNMIIN7CUlnQ6lRKh1YOIeAgWm006dO05PSOpMYcjsYo2pKTddAEm+J
PaURGjI8uXok3WxHXbeWlIiZAjpa9vizLjc/idyHWl3RPLnKmugtMdqQ7K7hU2A8AvMvqxXA4qo0
r345L81+WRmHxskOzamiIE0psYecXMT2aBE0YGV6G5FmMpfK32R0PumRtzlGvAWfNMDopvpcOmqi
mEYt+IdzeFAoJwtQYjFuEqD+IXUKvEpp6u1Wr4F1g8vzti9PML4SSNqPFbJQeUz1gawEqRmB2XUW
hvm6lfw8gF9ym9yIPrbxjRLN7COnLSkddVhQKqojvtq2en4PkCjVe3wa/x8cD7r+oENAhLwWhMum
z8cWuctxUsyp1dqOLnLqp2xApUMaW4X/X9+nLlqgpfvpNY35f00jdhu2jYgz2gDIJJk5oyjyw2Wu
26p/DaCGGGxxGakrMnWTqeZtwJsQRfQmTGeLcu1hjKn6on2fx/6avHT99JLJ3Icen7ajPfl34So2
sy4gDodWMW+2MuStocNs5JgZWV4R1f8NP8HSCHb9U8nFRsNOEUhuRRIERlUeia1DWHE+J5nFv8+7
pSKN9MCigt4aFLpTD/G0oVKv3IMaBBugNqjRIvzXYeQKFspOmKKX3/ZGZWWy9VwD1g5cGELkDf4i
IkZasldM5Oa0a31M3zXh1tPfQ1vY6k4kAmXcUypLvoaAcDIaIx63LCcJVex/CfoBP8/Dr5jN/YO6
iNj9MmdBb5IQ5oGivIfOLOBLtTDleoRKMaWmR7QbDxczDwPgm4N2eRzqcc/k3dYeh+1BFZ0dad3m
Ptq3KiH5dKKqyhkbCU46N72+s0bMnBuXKWZpUJZjUxypdCWwpW+Ieg0hd0rVLxLJ+hSg/HrO194L
BtgcqBvQYZ9GIrfz+kqlsjMuo3MIoPd625K9zAez5g/kIMKPRLkD7gP4OXSemGNCtsn05B8910Ny
BPTj9NDNFjuKDXpBOuKeh+0Bi8EIoQwwzeLAHhKQUBwmfuwPJZmUmRTUh+6/ilf42hbkDnqzvSxn
2ibugzGZXRgtxS6WG/d4xjxkT/eEkG1fAWFRakU8W6LdDZNZfqktY/llpSS464LwPOKrwmaq9Hly
8UtBa/6ri+WbCy29SJe+f0N2cfWNMz3jKNOFLuraTuLaUSVisIEbO4EEiPbC9qPnlBFipP0lBONh
svM50+DQZe1iQSJtTi6eGPvht01KmeDrHyEl9HOZHhDMihMRIwLfBO6/CTp9mfWFa1B1VkVFfttK
5XmRuT1S6pRuox8WTx9NViDcjJPYizDjhpIJ2cR3Jiwq7oeQY0p2B+LIAzc7RWVxMk5MeLr+t3hm
aSNSw7Mc00zt2CQUnlYfJ53k5b0fUOltizGvz7jqThR0ZLY4hI/Ksv22keEGmFuj3p7GHCvwjyTr
oTQ2D8L3hCzSFF4CeIs3evIYmba1flgASlDVxdJj+gId7+nJzXF3rJJCtPgaj8VD+Y8jT2ljFV6s
v5x++R7ckYh3048LewLvGlaZCNcAIGhADe7Zc/a6snbl3HcCVhk/SAMR2KB9QocPUEitXd4Czsel
fq0vcw7KRzXqcw3/9hinPzJ0gZDOvZYZUOfurJpgtDBIhZGBPFsHthJKqJO6DCao12xDRwhny+nX
onCq0dJTVack5e1WnjIkZXK0LAHdy5dagGw6s7IR/b0bVJ2ftQpzAOXivLy3bRkgQ7+5lZd57JkL
StaKokSkBvpYQnAfH7ZyX+kUgdHigxogeXO9UYO/eeXtnuExsHwp7oElDjfcdxRhFQLZuR9OViMe
wyYivsqfOMiG0kjvU+M614ijPmN5l+DGyzoQ8SWTp54+dHLJCEbSF8zhML+NFplxbVbYhNFMkJGj
J3cdBaw6L4uXobac8Bu689H3pG0W7gQ4GKmv0gTxRl6GKaQYCVG3T4r+jX5lY9vc4rR+iW+QZ/l5
K8VzV0zWnkJz3tbh8MJHz/1iMAOB3ZDag4tUlcMNeFc1AcWm+TP/sWwB03+yO2Oe0IFDrQ1xft1K
z8jMJDUmCWE3FOujOUUPFpJhukWFrdhSJERhUmDuThnexUNB/lMtNNzg5d0vo3DMCrIQRZqBXkN4
uVkpHfSh8Iy020MFyq767ZgxZMhgmqWJ5MzbrSgrZtLcAclxrgnLHeUwfQ1gqQff+EU08X7skX+8
/BYJuGVcIqyn9P395G3lU+p05IkZtRq+g5AUxvJnu+4u4XCZuja6oHDmJmwWcKdX6345MpDCaWr8
rdtZR0MB7nmSM2KTcl0oA+MsT9j1EXzIUYoMYYu4FyBiaZChNfbv/SQdhCI9gbwAvmJX3H9SKCBe
lrTCNNCc/KJvKE1nqEyruthPoP9k3BdsKANE/+97bZTYgQFd5iP6Gfnm8XiQn3oN2ktbOirJG9Vg
vh2jL9TVvO3EvS43s6msZ1GsBdpG2dkKcLCi44pgWaWUNL+QG48Lh6WG4azPdpkA2NoJ0pK556uD
ZUzGlxK1OLuqnQ5IVTMyZbFNI04wT9D4hnyqEUbUAZYSGAhaT4Cgc9pXKEIJmHlgK3pqPuzYOfy/
isPgACeCKPep4obKbP+EnfyjIONN0d+T11zs4PhWMCEc3ofPtDsoY5PGUQiuyAoy0zyKwBVeJYjP
XvRjqoiY42dOJ7er8GZLFpjJtIwc0coNb1KpuZYrI3XrOi7IaUInfPe0kHHvoE156AHNuwq9gNgr
VLE+fKso4l/dTT+xb95ikqtGbjOr80YL7jKWIGyEezGx4Pjn1YV6mSZ2IpizZbAvxKa+Fyo3w/ka
97jhu4oQG0uFB1lz4yzH0rF4ByXXughMZIeejm0ltSdej88izHJKNVIopOBKDO8hcPQrui1V98aP
DXHIuqwxd6ZjRD+I+dG/oGup9LTaoViPdCWP+0O/oWobKoszItWD5Xv9LgCpmUHFBKG8JzQ7fRxf
zZZ4lLYppnppIMjyLhX/4UqfRx/TvMHmfIZloploTKfN2rIDIKsmBE2lImLIK+O+HK2uZX5z0yVK
oI72sGEWnhKIQHtR/JbVNWQIic7wII0TTc2zD8bI/zvv/wen8BPuzrZKVfRbO8e9acGSj9+kCcye
3wpPVCVdAIeihHTeHvLTR4eeRF8ZG8e7i4XH1ggcEiLctwB4C2IFOqZCP7kNkrdgOpUKz0VGXhQc
btM0lr6nfzdNxD5gSncsiAmX8olFxPK59PIwVfXxS7C74DqxIhNmrV7HsOrIJam6d9sQIISMOdgL
u8++aPBywLp/NoQO+Q6crsb8LUkTlf+1L6Udgcpoqz7eSyuQULdgTNeyAda49zNnTbSWintHDqTg
m8djhRgOcBsIRnuhfaeFOcR9RjCxhwL5wGU+cJ5jRGz2J3uRRBL+ZcOCLsV8dfOsSXvnPzg+4Ip6
Ey2i6+nENVLda8ydwBp7pr9FBssbB1L6ljkyuKgtVaMuITRDbaSyORHQYBlVYRTfWgtJFGojENKd
u0Nvu/aIMd6zkIFL+dVmC0eG/az2e1q5dT2/76HZxQpRo03gtIZURqU/ClQ9jLJz3foKxTC2G5x9
wFPNkS5XLFDBMHh3u5QQAl5WPLW07PlnuWO01bdkHyaUIw0vfAh5l8f+Ak2k6xidyGVr55Raolc9
LcL+AogzlMgWV1ith3Fr39TgUEZ/e+ulYgXehr2+Pz/6fIKLynD4D9i6WVM2NtXGBDHA7Pau/yUh
M8Q4zrbCOSxJOCGE7EmXy/QMYbEdt2rKid0ZqM3SSSVDjRB2Gh94w/4/XHdTrQYFp1VYTmTfGsZK
omNhKbjY+RvM/ZAaiKPSh0o6I7ECserpJmlYVqsAzWToJoE2mIlusOmXy95a9xNRZaJ9UcNh5sKu
LGTujZ58ENVk7/gjMhjcQbt7QIqVHs9nY0uGdNSndaEoXwpi+JLNibdYXtw0x/R8HygwolIIfa5Y
Q/EB6CtWUTUlM/dwJJ9V8T8ibi5ZkNL4j8aAu8oquKK7knpt6aCo/MyJKZlczPS9U5dVc3xSNWpl
BB34x0a1jhZj/DmaRhBXW3CrLxLso7jBFs1ix2QCoZHqaas48PBf2aHx6u5p6EjHt8RIo9nxNY9g
S02xMjpTXS8mh6Vvqv3Ym/76OAQFbND91FDjVyb3D7S+L9rzfPCVcgxQDjxmHcNDawKWjB4xKYF+
/jOE/CWFzk4jKnUUlpcsdoWeqNtNxaHZNoq8K3GN4buAz7XuBHtry7qvAgp44drzMLdXObVdfS2N
5x5KvMS02O6SPDEz6b0x4L2OzMH98JQ/mblOce6nzMbN+JpLwyJRbYruYJMIesjzoH00kvbQgOs5
Rf3siQTf7uOvG5xVGJ1OfCTRKlGL0uiUGlccG52JuhuLvzDHFSWCP+vzqke7aamMrVCmcUiwD189
JObVmm0lEjfeG7ZCv00yKjurZCfhqXu+ULUAw3BPe43M4SlMHtUqKgBqi2iPBIZmWwqESbH4afmR
3SF7TSsQzW7Y2sUd7IR1U8y47401WaYSgOu0INrhJuTEObMS3NgyzndNoK39mB5x03nTKvlNDj1E
ASVvbdTYPzgApC3QVmYJp1HBoh98pXlqtHFmqr02ZXeI6SzIyMOY1P/TGzAnXpjztLX12MRDhTKo
OozHZ/yYNCfblvj7ZaPqgyUReFHD/y7AG0ATubMzs+qS9Y25qse2+BVO+smmCkgtmSqbHFglA+X2
IOhK2q7IQG33YWZZ1k48HggovErtjWA4YkwgAevWytcEG2hawZyWbfr+9OPH9NQughW/4Ax7DB3H
qQ1D8b2OjumMAM2ZeoDROAO0jfvUtO7RsqZZGDdSTFHKOMZ6P6VtpCIeppgYzCUW1nv9Kasy3A9L
2qE09xdySvv3d36pLxpRGSa2SFEKsGkE3BhfVMN65N4kGrdV8NkyuePCeHXiXob7Fl5t+uK0FsZE
OV7XQ6NS2ashSwF3qguJfjHxggxDvcH6RaYnkPvduLsyMdb3d0OFa8j3juBjpqeRkN+R89U3yGeC
ZxLxljMSVDU+YqzMdvEjPv5UiCIiSuU2gvvqAt+M4vGq7fRYwKRtWhmhmnhwjXsK2EFs4dlzWeAl
OoS57f2NwavYv8wLEip/dzHxieDcqe0KMY7O0ghw4OusJpz/aU6DrqoIbGtEoLFrvgsU/UNuz1Pd
JDb+rTvpuEpr8wRfTcr6KJkkx6qymLajb7tUi93XoTfbJNvBeYy/F+BQxiR4/pP7zpHD+B/hK9dE
8ukePt8Mi4kcLAh8qLIOVibbODDaBllmsmo1Fbs5kqYElw3csT+SbwM2gXcmZAN7VcDCY90BLZLM
YIQwM04oJ98QQ8Qx/lmcZH/R6xgpnsr93p0utMtrcGqaLDbadj5FiaPrRGF+aUXg0/pf1FagGVVN
yYcxEXTQlw/mU4TX/bYby1Mne5BzQIOyfJwR9oBuFGJVupcI+8xJzXJjKrCYNPPtCJ16fy4NG+aM
Vwsm6Rj1HqvAxLbyipeoKGgjJfd0GlZv2x/NXtNZM/HbeUjF0FJSbafxVIJFDpnMy9wAsZljinFd
NfBHtwCYum5CoHf/PYMsEdLNGM6yfhoHFlBFsi/AhzrYyyR2BB5yzFSfi9dqqM4OeUmRpMTU64pB
J1XUdlq/cPg1FVsO92s7dF+ydYv46uN+wFtKud+ULUWolTxSQDJwAD+52gEDL8PwgugJuJH2peVd
LcaNYo8ijfdimksvDjWmnCCJi1fXVqiYSoqvp6NkuLPyNluP/QmQxsMH6+i+lt8Bt2ekV56g0n+p
cSHaxfLqpX7M4gpDBILBAwKIA/zbHEffFlGY9pK0XIkfIvsoAPBiwLX3N/YQZZ9Z19vatre35vok
SGOJlkgswNxsK3aZqG8VoxaEe3l/LoJEIoqtcxAKn1AH2n4r1iH+kyJ0W0vS/GYbq7LK/jHfgdtE
SzKRf0kzU30roaewV4miXg9u1C7C164cKwDZQnUiUQ6GgmrMErEvlpgtHGZOkMRPOIu32p3rglLY
RHbhx5UgZIUrhBSDwcdO4JmP0o1fggZyxyVetos0B3oAWUQH1+gFWV/+nRFZVpe3AIbug9sthqnC
oCfg1/UhJbW/Qu2mOuJb1fsRnY8x1lWeOy1J+chlZsLFt5wMwTRsCjy2kTQ5wfSQTh7/NuoU72kh
E7jd274uO50glfGHVPU2/VY2cg45ZAcJnHiOf/mHcb3e8Xdu7tLw6HDuLUm16RWVl4w6D6fj3Dx6
zz205fmJWwh3Opoxs/tsvDnj5r9q8zdFLWGjX5+GdH8iAGSO0S7/4j6WMpuqsEzIZ9ZWz2CN5XNG
tQirxKt1kp7n3YhYQWo9qvg6IpTTPrQNvd2v7/AXlWSuWvwpJ1SDLQU3Ed9mTqOvpz5uW+tKaQvs
fkw+1Dticd+HiJFdXQVdQFzMfXQBlYWHdrFjg/KDxhuq4WjVEoqWDiZ6M6A22AIjuJCpMWeImjRb
5Jok2JGr41Bm1KQTw6hGOeu6GRYWhvKh4kT2cDmM6sYIEpdEAnLCB5Exz3lFyjJ1Xe4NdmbB41Eh
aA4EErh8xnEosFwXIXGKaUC7FxEcJYkwcLCQ1a/j/OVZE17t1X3RezwyLILOjekogpxPq4JAIGCY
32kvxEID+4RostXwpawXy/3nwY+41MFQ7NmtuglLcJlrt5WiqhFZJt+jccRnKuD915WT99prBH//
LJaJnS8urGPPdZeWXKJgZdSAu8fzX8S+I/JBSHilKWUtXCMpHzUjz8s2b46/YqBRMc0CNcG0ceQj
C5SMcvbt7QCGd79vZt4LxEsfuXPPOrbLiPmy0VF7eA+QfWkjDUwmzuRdl3EdSu1i+POL/QM306eL
HXzKvgvdusw06lzINv3PjvYWDZLzbVQS33xR3PJ1njF0tIh40bjkxcfFOm1z8h5t9POFBiqIQqCR
UoocZLU0oo5BaicHNGhLe6efhgE36r+siZJELx8GJ3AgGatfi4OGH2L/UaMh5pnNo1cTRvp9ihmv
mhja1ZzqTYAzgpIXIBg9FXYXG5b3DzTWwtdM7v2//JcK47RGfrOXGfsqr0awHyfSqm7y4XZeCSzA
3+wC1OZVQunG0QnFp+ATajCx9esahuWMFjUnc2MEF5m3Ztv2N1eb8MI/o3AnICIlC3QWbqp2IfIm
FzMrJusTn5QdUgluLeF1CKYdJO8idtTTSU+Y7zFuRFdf+q0V1w8EDz9NCxO3+FUkyFSYnnJaCzuR
5YPnG3FeKX508tjAUQt6PdFQwWqoPP5DDew/ZxfsS9P9YdZz0Ep4ZEzKA7LgnwqL/V96TIjbxmRg
iCtqoaZYmmPbM4YGo7nMvRSellHJ9xat6Id1+SHrH+/7nubctZEFDGct9i+aOPC4bmYHuM+LRwg+
Nmmlx9ZCLyG+BapbjJ+VEY/Dj5pw+nyMLhYLIX5T2VS8gBmOwW7X4OPWh9q4RQ/Aq6zNAkAs3IXd
XKgtZeDxpfWNtP+4eD1Vi/Ihdm6TnRR9VvkxOCTqZJR976OSJfVv6EQu7pJCqmJYpp7GrRl2tyYB
4ekoWxJWYm38tBX8t6EFAjY1GVX8CqQ2fpLZy4Bzd10TjKtBl+6mwcQ+dxDT5N1B25NC4TLlgzxw
xttsIQvDa26ceo04wxdkzcsLWgEnPb7xhKuDiVYbEx1II+RiYl8rxRnjE6Awq4avKVy4sLNUWO4h
fnfKRGJInThuKeaD2qfruWqfcVSmRgYAfjLAc0S+oMod7HjO2aaKwLsE+Cbl5K8o2eynBt07TBtM
KGGxEOQ4yxbVe4L4ptQjXQf0r4BXbwvaALmnL1Q4lvvRasjlBKqqIc9fzHUbgU81kCujke++GoI7
RfTZutZ7a+Hwzk/tnW+pdgdVwxR8sSvyDzzsiwvBMFmlJoFTO713GEFqkRjm44tlSo+czXqpfU9t
qErEJZMuASzExHfZELMEBa51Wkz6k0+TrZG1raBRWq4gKwRx7cGUUu4luiCbkqpETzDo2efUXGKZ
y3YQzUdE0A+gfkIV8YJ8kts3Pfy2TWGM662g6JGbZZzqJTjA4v4uDuVW+0BqAcDpurzKkTww77zL
udFn7oTuosIVbUsr4MfI1lIn/teKeNMh1e+Cz9CtrNuezauVdyhs/p3xS0s0gmgG+Q0aonI/WJO9
76PwyQwz7XYns84y/9wQyrIGa8ZOrxDv13V3EDd5rqpX+jloT5GUH8CCCti3TCNx4zI1G5t25rTo
8Soy74yZAvSskN9TJij3OpfPeadSBNmRZDshTVjRiXccTAfOxpxDrJ5y7GJ/iN2RupTIcaohANoj
VXYyTGMob63JrJ6SMsKc22BgXezAQqjIfk+3OClgGI+89pCRIkpA25V+TEl5Qo0xG6xV729vWxIi
t9qMOM8bDBJUnQRLDQp0ulXKMrZImx8Q1My9CXK42kdVSjs17KzSjm126kAbFYMymB+2E1vIuK5Z
wYCni7K28m2eMohwTThkHkn28MDdT9q292wojcgG4QALW/b1+hRDKEDfvBR11IOxEKXTJhYFzwPp
qRAPGAHTob8BgHSibj6uTfUhhdHmex3Ubja0BCXADPupWpb1JJ5tLZEawMa3T2W+S4YmuEVORXIp
VpCu2lhGJlqJuutXE3/qMRZ61Y23hM08tGdBhuo7HDx+fTf+9Kmlqu1xGDi5BlaYGGR4FFT6iAPe
VjbRUHqxVxNLdMLR+H6Sk3aLvfx+g5ZG5sArYfyf2lYv1S+BxEHp1Gj+DeaxSQYNi9eoXBOMNJck
8JrgBvNXYLyFMGDhoVfh0Jb+aBtIW1WZc4iwg9euz3G9CLwWb++geWOx+M4yEgLH4NI00V0eL02o
X03Q7tnkkZpTgqhBxVoXE4+h8DurtMJTcnMXAFJQVDPA9gzQdoZq465JQMNMFcCZH51IdclxvnFm
cYoOncKmFwkJb+mmeYJ5F/rZSqA2e6+ej2N5g3sYFQbKQVRLaZuWEMsr6AtETSm5D9BikCufo0C6
OfExgL7ss36TiLiIukOZFMoqLpi7wwxE2PIQ9hEDVOQXBMmpPj8F+sUpYRZOaGkQdWYgnuhBIa+I
K4R3VjHSHfzLVPapEWX56/vg/3BQo88woQzz2iA4G7VQho8C1FJPD6I+ce7OfPBVfccsH/+34k4r
zAa1uHyuzuTmrATkoyf0KTYYwg5ihyHsmFWV0k1oOM7QiwP/g5Nv/uK8J3vmQCQxHuFGkskqDHq5
bB1W4SSJ9WoeA0OzyEtJljHA8pnAo3e2TYQamPxQW/8cJRoj56duAiMBa3xIMc6fVJgt5VuNJdmO
ID+fEqbGZB2P0nUVs87ksBSQKlEjyeStjGfxTtGBLzmS+i9DB/aC2hwm0OT13fzyMZX7ipcKYTpb
c2nwIQ8mZzzznxmqec284cRqhCbegPCYzHawThA4l+PTdJCXQqxzvtdb2ZMayRiVaa76r5bC9RgM
R/FFPQ+cl2nvatnj6vn6qacC2fbm7I3ABZnGvMEYgsBrRGDSDN+a45fIs9jHokbOZjyVt/yb2P/X
qYjsrPwqHRPUhGdhXGX1vjllwb0CZuz1r4MfewmfdkMCToSXJm8HbFLdJiAuKCsrgOwuXtYLte8N
eR59IAhy+8tOh948VrzgjXacC3rnj90lSYZhq6eIvfyM/yYiWZVTJc3CbNJLmONtRnWrYqG1z59q
jK9fq/8A9wwCBt4ll0H4QcYaIlsndVKTPCyFw+QFhq48VzSR3vST2piK/Tju4nZ3yBOPunvz6s3t
f1PWjlx31W7dwSB3Wg7GjAyYAFYWS15cWcTNEC8Wm2usZlcYVaZTaI4cY1dvVA6iWt/isd3aSoV+
n6RpqTlBPJ4b8HQERBLt1cS1bjQKV5b/mk0FY+zggGnT9K2G552toyY+jjm4K3JvyAqMs6t0fcLk
K3CDFyJX5L5dZvWXb+nmcHjAFomHgIGX63AMSrLPuS503kXnYYoR5bb7liaCqt+s31uyirhW4Fkk
bA62TRXizTuDJHHgLond9MzVUtya9OAXy/BSEEQ+qf8KDQDB489647+stDSGTDpsSV8ixybPpZyT
/JZaFHhIwdfbRV+5eULxSouUrNjk9nd2jTcidgnZccrkOJBvJSM3yC5GTL1ZNF6BuPok8+liNmfF
kSuwESlBq5rnelXC/VPBXYKKRvxh61DAdXQahl+9xMOxOYU1q5N6HOat5VlnWj4CLRXS2ddnR1l/
ke5zbmq/TArRZ+oJheRFUpPgFTTEfYpKMBjN0S0GBEMj9rJ6vLZGxGi67SViclnu0tjivbXYlKTW
ONyPEJpyAY7YA/Dup53GpzNqs/0YZ5RZFVOTI96PVkgs4mAPAyTreHyZ5A/7uCvpU7I7Qn4M9Qyk
CZZgOxbf3KQakcf1P5GGjNWYmNQfW5mlGt2lUvlzWCoHy7+med/THK9u12n0jnufQkArI4yk+BSS
b4MggfZVDW8rh4HISa/5pMG1czwJFiCRqSxx9YL0v3OXxt72k+Bi8mqzeYZxQ9uYVViOfEstCglj
Pb+TiPjGRwDUjcFyhh+BSw+J2CMU+LPFgD5m6dMKHc0qy04woqjfnX4HxQIDFTspTHos+R3O+FYs
NvFqgofUO+N9/W3mzwDFxKkwZtq/tm3pbJ8Sps5NYsj3dQJHCNboOXzo3e51bXdJ2bCtW5Aa5/K9
GHnkQGkDYBV4iC4B/M9bVaDZG29fb+GhofuNymCmIqxUhvVsKjTjV25VBIKeUrFZt8waGu1Wsfx8
cLCJ7/d5IL8XuOaQBo6tkNlGxOATJO/jXGE0HosjU7n/7NW4cyrmdv0jilNTrgDKz0VaSRn1Z480
E754QEGM5e37Zzvj6pCH3HILU6aKTAuk+5MTHqWJe1SHrhfQAS3ufyf7QqQKcWFR+v2DN+rkYKO+
ejo2aZIG+ok767YxoZ8kJA7fLD0PHv/oNBgqSOMiXCmMlSrNSd12Fw4NrZ9WWPTngeNT+OfTfbM4
tDUZ4P99endYCLVAB5V3WUBTGWXmvNMpBu8ihcalm5Df/nuteOQHbp9uv4IZvcwEsQpKCueJPOWh
zbUvrWfGqmtD66yMDz/AMs17h+FbFg1e5n0o/ry5BP37iiL+hIWU3YwHbEGViUd+4knpKG96Ve9g
MV6Y2mt2MgwDePnt8/bf8qsSaS922hlpk6hX9AnmyhXPPi0vHN95Mv5mpP3QHh05NTozVp2K+Ltr
BBrcSFpHduzQ6kAScyd4KnltiQ5puYIv0HVG9sifOORygp35ZxyLV95dTCgjX85S6uyxO6y4BEvh
xGpsiHygDCWUltkH4CHc0FsJVGGG6cXpdQtMXOEZfEKW5sy5U6h6IRkKksLvgCGp3QVtL0Pi8Gq7
QdqtQ5ckKVH/+QfmAYt1sNywKV66ecrQXKODmjNKiSHk590enTzhBU5EoshxIMF2Y6bzSd/s0dz4
pN4zMxbJ0BgWp5f+Ysx7n3zjZRPR8SlBwffzaGIEY7Btc2QnB1uttkZsHjkMbV58EoFNwh0/q7kj
B79YIyf8/O7WI0T6Q9vERwqq9iX0Ej/ASBe2VArwQIG5j85OCclQkeIbmaEHrQ2IBVRh9mPd479p
q7VQnuG5gLNnMiGvXXrW8VOj9KdT1kCEO+vNIkUnz/iMuX4jI8CgiROevGlRXxct3lr7pHOfWNJv
1JAIIs4h5pjY6Mzc8nKwtx7bR2ww/H5MaHFFMd5+XrgLXaKsshKjdQwAxE9y7KiSQk2derOz9o6z
aGu4Llyowal3/Flh11q0J+iS9rYJ3jglXwcAt5iEZQ/nto4uznqmRquWFlmdxUQExl8z3/pYT10G
wSU1eoEQ7mfsp9UDVQ/1NManreemu+Hy7AT/vWt1TyIOpqZOrijg+snHE6w16uJN6h9UMsMOmQPp
1dpwwE81GosspIYaevda5Sk7kvk1HLv5EgPcZ1+2oZVWc+WHOqTeQdTK+1LqRRsv7GQgx0zIYtfI
64WZaWher+h5wdfc9QZjgLntY9oZpkgUfSgSe0AXxNs8aZG7ChRHiuqX3svKK8WX+x9+azxjwYuq
/gTbHoe77MvnmhWBv4+0hdabehBP/ydHVJ9TSdJYy5LUjNDC5RxsowrdtzzBkXbIZJQWqvaJ1ivr
RkHjpThAdRBXM02mrPe+0tDq7Dhm87qCxWT3oFCW9TwgGrjLfnWgkoqJAuVZBnK/MgFMk1mTwjoE
B3Wr91/1XxCQWhhiDKGlSFuUGdqxmYuJXAn+AxxA9fXWwvVYqY97uNf5koFy7XBNu0zha6J8JNl7
CZlHY1C4GwswhcfOQvJp6skgchl89bb1Ec96dJUJcae2XsGqC+UNq3H8697/Lob2VjK1UHVi5Iip
jtRSuRvrva+T58XccJExmLwkvRoyE9D5vBQhHtrcGfs5MweG/xa5CxCuYE5WVyDTj5X9K45LCb7e
ErnQUiAFBodulY3kIj5HCMKnzxjP5nQ4YXuiEdc0Y81pprfO2pkQw6WD5avQgTFc++5IcK7AiCS3
1Ppal8XxI9hOXUNrKaPaqkfdCEe1qzPw9vD4OpOCP66LB1CXES2uw41HlTd0pD5N2jDan6XfZzz3
gjb2lNm3zMLYuwWaTB75P1841nBc0ZqO6qKftfqQvWLSafyOPBLBLekEtU3xvC2VjW37u7iU+OW2
AHc+iIt6EU7D10OBsVe7O6p/Jsl4lkTd+sPWlkGpKIDnjjnDZ2EFL3k7slCmuFAQ+zUZL+dYSeUL
PddKEsc4n9BiCASyPzQeSOxnWsuuep4j71EnK76gbkVtbJaWdjpYy7fyGv3D7G4HLqgiL5+S43oj
3MmYhfoo5wWzc+yr8KcVgYpPjxnGvNZEii5lDp9sN8L8O89kp48szthwOqoZ3dxnqjoMZ26Qr5N6
s6vxfMQVvQcNgcUuw9mi87D/XzlsZBOK4fV1FqJY5u3N2M83UJ2wPym6wPR7N2vrIEQeGQfy8fi9
TL42GQWoP7B8QFJ/VE+XISAlfODGo5/fnDDnf/xIjUhzj/QqD4rt3bHtrVvx81jtN+rIutMm4apr
pVPulKgABFJsdObHBp0eSZ47XI5VJIfQ2N0j/fvPa3de7SDFUTEp2KNmmQJ20XgRtIYfgflq7DLk
QDc+dKWGlXOH1iGkommt/3n+bAE2Quc29CbqiOznCGF+8JyGOOQLYXzi3sX81MFunG6f7LPLl7uK
XIe3liCyBXrUAUsPBdCFnLaG8BDQgJ/UjC8D0JfXbCzUPdTykrcUlQyFoFKBHkeca+cRrmR5KYE5
lMFUM0IG9wlobKXl9C1cWPw5RNJ5Y8KfBnGm/dSWrpaa9PH0epxWLWpgzdFTdkWBuXcxJkwqxfA6
Ow5NR7R3R2vOGAHf2WRT50TV8+sUSgFd/Vb9i2sORKpdWfWsF4crew+L3fYfWhmGpdpbUE8H6Uhd
jJiJlFzk9o76IyxEdA64VH+MW6G4BMYhmRctSpSLYTtO2IZxzoPjYMTyqG3SHx4MMwnLTjNrqA3b
2QI8HUrzar27hyJi7111ZuRJygZ4kbol4hYaxCHehXmV9Hk5WftkDvNToOt4m6EzFfL/mRVrWxNK
0qpz2Gr+qjC72BmghoyAfHxG58uSefXgLMY8Wn8pWpCbsOrqqbQ3iJPTc9fSCFZfIw9r8/UoHrss
zIFEmPf98bzMIfBoDKNnzbIX5FBuAHQmJq4we0ffkeE8E3ldN/e9w3rxhlvkONnR/7h/8LcNeEmM
a8qzdCczUOVP+EnsrKHsBZvJYHw7BVIlpRzUgVD1ADqFVt+lglqnIEZmQROfzIqv8FMAdujAoci3
wXmNz4qtfOw/GoPTiOUFStTZmtRUiJFF8WtErSe+6DZsJDeHC6Q8PqCTS+eB69wPvQGtwW5f1A5s
v2eABwQG0zTSEagxYcETPJFgFOprYOC5CMNgF2bbYzqG0TlYAuC2LfihfbYdEacw1jIAJcRiBqxl
gvffxTT08RvQZuozbX+Tr5QfkOddOboLjyORAC7ifJdN/gSPD54lK9C/cG/deW03ly3+00Umomxq
wma2SFjeJSKgQtMiryFf+kiQutqMDAznqFp6UabwL17Q9DoyxvjW/85jPHSIsybpjW5ii7wa+x+a
KPBfubfwxHiD93beyhFz5Z2FuawRpTdNNPHVXKmWPWWB79BOGlLz6RnCLJ9G71eW+qv/FRIj9K7B
c/jveUbp5jQJugrxQ6sljq7lZ+S2/IzxIaQSoRPynDJ9zuC90bwenl8hdqNly47mCDPpXDJPIbnP
+ouAoTPnsuKUXTMhbso52Gs/KltPXzOnUH6st5fDFgRGKWd2lecRm9rk2CZwfnxePRDnw6cSnAdE
eoijE4Hc7FrHcu+qdu1Qt0iYcs17ijG6g72fxXz83EQQF5nHhisQgXpBEkiD6wdlT2NTGn52qoqM
z0ANWp4ujfCKjy1uSfqf6ssEfIpzG/UMVU4rEugMy+c0qfETlaQvcZ2eoK1UCTBf4+/sD0plJA9k
FTTHTDMwNa7p1cW3MALI7j0Hy/F/tYjTVt+4fGOMRceR7GvHbm8WWwQ8goT3ZMt3tAZr6kDANks/
Ojx8HsJO1BvXRBIaQvO7nbDDRHF9UTuoUGOt9Kyj2nPyWKuKuRZ9OwXg6WouZXpBc0v1Y0Q6hg2E
CxSXTRA52ZpwBUy8+i7hkWYgyLIkulvn/Ysen1juq9sAc41pcZKroxx0uiBFasMLC9mEXqKQDHnR
RqyvkjJLkaSndX/apNRacR/BBY+/yf+jcilzJCPeggi8m2PPFWZJMtPtMiJ5P6gERyggPyEtwWyF
6SNULtyobNo8l8WXZP58wyqRkWMRGIx74kmn9jIl8K9YcDZ0apig1AWwt2Y5jUPb6KJPnwBOGBot
1kn5wxEuUaqQMPpOKAOVRBrKQJZ0Zo5lalmvidXtUyaNmxLG0rE2h+U+1jnktZmkwF3Hi1GQzEBT
U9S8Kcg4pwMgSRJu3xNG89yL3hg2VjjjDP+sda23KHLfZm5/XZjKKJBgipFXKyYL6UAxmh0gBw7l
nhiMoYXTB8NznFvQO9rtkiQfbp4H6Y++N8wC4DCQaxXHDCmvNgYpt+4/DfqU0gyR9qqIlshR2igZ
GCrP53uRz6WCoudYoAF07G332mKgpRhI44V00TRt/3hjFP0WIjHq+5v25+AMbTkoEnmLgzy+yrMw
2PAS8JAOXlvYf+h9UVNtyl10QebKhV68/uYVOGqem0BdqkgDlMe+y1tNFdLcUmr3+66o6IixOM/z
H4a0BwpS5mGgUjhQ3fxtUswAcRveRQUk7wMOaeO+ivjBzHUKcx8VuHWgM6Vxk5QrJBwOOt3Ojnxz
wawzUNN+iFs9P2NriUHgJawiiv5MqAXE3tADvqn8gW2g6p3onDyDGsID/9HgGm8AA6sg2uzeqOGQ
2CHerTHxAosWwAs8ssEpqmBUq8FQfXMOb2G4BCD6cTOCSyW2PtVgTiOmOC2NRA4UT/eQT5+Og/fe
IHJlWZy95ULth1uCghBD/igsDlDTQeOxkrALSi48LxbQGiyN1Zh+z5yPZbqJyFxC4Xqsgok/IN6Y
zi+vvgbxtp/RV8N25h3DUa6OPfbpmMVixARPQeEoPSiQXZBuYZcbDuKYhCaRUJ4CN7s7d3vQKCx7
NnfRiHEf7+qTSvCUuozm4v6YYamGC7DoGY87Rr99Ztfz10rhudOf3SHwYDKv1kexHgFhhF+PJpr3
CQ2WpCjvlJorogWvSI4IN0OEs6NMYdkOLEpPPP09w/Lx0/y+s+UaBIt3kyKwvqZIPehuD7BmXt4s
9+6Mst/nxJcijB4rXXmf7ZHQW3xfblv6c4mpS0YkPGLbsIBBECs4p2kxpOAmGwjFbPEgtRqH81MS
8Fy6tl+dIdJvnlCf+c81zUeVQhT1hCPVgXSpHnlTdSa7eFOdEV9n45iv9ZX5d816r+QiHgBdbTnT
vKA9aTqESSoHLUcAuAW5D7w1QrU0SK2U4urIz3Vm+ke3dzS1dhQzmNTk+kaP3EsRLNwAEZF+eZfa
3uOncryo2d42KwOu25BgsjJSoZkdzufU29Jx2UEFvAzwQbz+8yTSod9PJbns/5KINLsAxbsKx1RQ
f1poBD4Q84rY952lvnU0CzyIMUUSt+wsRIOV+8jjCCm/mxD60ai7+xIDG0FcZXydYY2KcneK1raE
N6KrMjI2yjAjI1K+YieYbXK/6mbUBigovGjSyt3JzDbisNAgca20TicbzzApd3nlBmcxGX1lwMPI
kvvT4cUHCetosytg21fV9aUqjBrmZ2qPbYzh+O2yQFaBJcYnMJ7JlU8xWOBvu6DuiJ43V1cYaVQl
phhsIUn374+izjNKs2vsom/nUSWPqSp5kdbXPZL/NAZn7US6t7f6l1K5lVi3U3/Iu4ebymyyoefo
8IEzEpwtcm4K5btwelkDc9I42AKPEGf5Vtx2emv6Vptm0AIw6pxMqeewSsrIx++brGJNyJ+yrFg5
CSqrBzJhwh/PdgvVB1KsfcHTa1NHLJsgRfjwq3Dm1NmQYaZbqapm987BAeTvBxP+MtytEqlozjZO
/ma70irb2kWwHMnc/cjmfmpedUVWRx+BSptFqXbsbkIxzBRJ4HwtokrvgmSVkL0ockZw90ywTu99
WGQyNoveKGfBjBHt9ZGw8mg+imjBJWVIBbOqIkp2CZ+hwiZNeijD4rZY0BjJMQCnXcufQxJ3nFt8
NAUmT+WWTGsdsmud2YENWq1VslrToZG01KeUI1iW7uhpyFl2mbcHcE/yh/UyalzMcBCZb/cuiH77
sKLUzSZjEW6tLLH8o0+FOmZGAOGn13th9vFdRNEoHXOQV89jK/cpTgx6w5I4IhQp5k1HnN5VixEZ
BmMB3DEJbjBaCWsHxxW1iwbj/7lyq9A4S4vSwrK0+UcnjdVDcGcmZ+JZH+CM3gbuFDqfXGV9ZQBj
9Pe6VhkI0Zvz882tOYtpPCuUBQ/UZoOhRB/Ll3oQB8J11mRiXZHRLxgGuoxnyZDYF4y1H3/ni5Lq
t0eMD2gA/9lbjCVHF7/EBGZtw6lHuY+WqVkWWl5TChWu4U4g3u4yBjZMMTtTyX//VMkfULXpoytD
64/kSM1R8ymhDbFOjGGoH5jriPbsUC1CpS5CEGVQR4YuOF4TXTsASQH7YTFZKL4ZkGXSgvH+BNr1
XooHw0jXQ+iwWkECrDbfgzCKWkg0wQK/5/Zs/p81JbNl7W1qNAwGpW9gStEljIyjcCBeeed4+3B4
0QHYSXyLGqiApKiVAsElThPAKjUF3ttnY9e1jzuHLlOIyLA7P6W+8JPVkO6DIvV0/OmpXuMtm666
uUUg8876QU5yAkpw3wAO/52XXp743ZWZmITkzof6uG2wEMN9soLyJbPX44dw77fC3jNdOnIpdVW+
Pm969BkmNuYrPUnDh7pXQoqbqJypS0//N8L2AnyoWz1DQq8YVdcf+uIImLSo9bZbwBA2T6tW3JsL
dP/+oa+iXHdA6OTjimzzzVVt5Dn8ynz9IuLlUi6/AMdfNgx6NSEYuQJwF5I1ZO7dqwRro1FHDs7W
VMEcngPEAPZxUq4qyvducLFe8fElTh3byd/1BqgtXcrRgT6PkJ/15NAaECtwxGmt3xRU8HufmwfI
yf4mBFQKjKou+rFyjswONTpdYpGtyYU7/yjets0wQtshrW+hoWP6kvyMfUCqPNyoz67kttbAPC3w
uGsBxED9wms+IWO75hPkg+gMMHnRS7t9d1DQquC8W2S4Jvl3fGOhHS9ve6VVQrAmzp3C4veDNZO9
cczSs0GpYkScpHPnveOeCna+I2vtw7PF0xxnOFoQJW/NjkepwhajFVg9mloQpk3hmO9ishzP07dv
71GSGI2JS0FhKf5N0zuwpKibwGhG6DqYi1hgxJJiI/nS+ijGuyjJWFvIxnLriG3ha74oNo/XpPtn
lh+cu3if/yWtiiUp/b3Oy/xWYTHUN11ggbESuMnOV00EmLFfyoZAw4LXe2PtWr1jx1UVacxUKcLK
4ki9uftYDXOoWqU1OAYhu6O/wwNeuo3nHDfYnerFxGDAdIFj0CVpVEhdreHpVNiCigIW1Fontxbf
Z1YmWGiu3Wm70/ARj31Bzp2yHk2Wtf+vCAIksvno45itC4PvK1TbuzILnXdv4DI+QZdWYhb4jgUV
3/yyLo180v/KVqtT932TU9XBlteFILOtu+bG2XS+qNkSmj6zlDYvOixccAyXEji3N5DmMMXaNsrO
OZR9yyGLV0Q1gVcArEt+hjCYhbVdgCAbkBCi9b0C0qsiMcfJoBtCuBFh39z0fYqfG9CjI8dWLZtI
Sed2VqEVoHkcpBvhRRLZUIzOaRy9lzw0KTUSc8dCJjPvKDJU5YSPJRUHy+7aFV5/+dbSa8Hpeqcf
SU3RjbFuOqgRYVUbmUqGj0pbFvHL3CpGkAdgvjiMhocm68uvW4vBj0NTCgtl5l86sh5WUXH+dYDL
5seZDkLlu2369dX4uXcVBRvgbn4qWBZvvn0B03OL+aZAccZvmklLXm0ReqnTbVpom1My8Ev5zw+o
nf0hRlaUjyTXF/3aUka5PPHCvy6G+6R5s1lw+GrOfTVCGBlKWmk5TgFXnCnR019F0PPPFQ1BH21v
yTOHq0uDCE2Vr9sOuv5UgTUTND+BLeddfH2nMN+1yx5InHofnagA0Z+2+wq/y7l4I1RqHn6sANUM
XJtB5+pwpwk4zgnRIyeIFT49d2VzbTcnIztOkxDYsUMnYL7/zUI7XMypsYwj3sD2vcN4U4zcoavt
fuA77WFMIpziA9F6ADzJaXU9Nu/zRooeLsRwJW6y9dg0N6tj0KhvG6b0UfS8s3gNZSNY8x4qCuk7
jrHqlxJFR7OoTYd2/EpzOJ/2kAEc7/h2cySjrLCwaPevsaCFWASnPatzM8jKISjbMKWX1GfyvI1u
YXIinTjlvYp1I8r7oOfDu9EojloUy2UpFMpMjznffVwWkrTp3YyfeYJzV/Xej8LQDXDNVQYyeV6V
iVtwTFuNH2O6zvhasEZE4J/irFq0gab3CmHNe1HCZYgKvFfciR36ed1KYqn0LNr1KpoRf9PBEK5T
P+DQlAs/0FKPWzeq19lj8oNIOP3q5OmiAR02n8e+eRcrNGHP/4RXnVn1DCc2Triso779y6vr7O89
UZjJ7cA+UJhpVMeZdZQL7MnQ2S/Qo3etMbrsjx1c9+bYIqBTGaJRMT4tskqCy1rVMjjpe6gP3VnM
Mc42byCbKqkkzFDsdFtBd9doTB8n52ZNhIMLkcpDGcnKV+4z0Z4UtxYvQr46DGLQ4oPBviIQTFeY
UixnfNYZxmdkgpDj89cORrY+7KzR5ubbZy4Yx9i+cQ++PevXZ9CJRM5g1q72ugnF+Tkz9FnKJaep
5WQn5crQFKxwR5fwNXODFRdGS90oIV+uUhkwkMT2anYdFo+RYt5oGarvOjfRz+IgZlk5OYQkMtnE
tH9HQrzzzqh2rWJr11NdBNUS2vcU/CWQ6OSrGifGenQzLBJOlBlvB+dul5JXxW9RI3MXoiD1tuqn
NeIjoQ4FrShIdKAt07QG7V60iEBFCecVbmmPe5Ghv0lb/M38AkCWqUv7EYfAv97uRGys1OGCKPUf
rk5/vXKt7msa3ghyQGkGn8OCFi1MoQMReApJH53XK9EGWxI93E0SM5jgJnWB1qfORX1YDuR8WDdV
97ongKZvoeDmzwQXgpNB81FCzjpfUQcZ5J5xN7+wfK7PzyKHzmlBkNJemBQCzaJzGqdMuyAU99pg
5MoD98q7+5sqSs9m9ULxcdimJetFsl+SQ734uc4nI7NjuS/wfQn2gvBHO7Zcf99uVCg2iBwV9H1s
0IhrCpdxhW0Y5LiWVP1Y7KZf+yNWp91pE+7j0k16RuR24gioLw88lwxxWS8N4N1JDpBS3QBWqKkX
a1pEe6rKv6G7/hP4GhxUTDTBJ6/1hF9ATfnjtEf3fV1kja6fsOifmGeQMP2mXG2JQKPYzKZ650aB
1zPsjIUymzVuknw0JhLbLlFoht3qjxWCuFyOIWC968KEp3AHzbiLn4T6YshXdTg6DF5X76Gz2ozV
1yMauSbCkihpOr0BZiIyrQFDDj3TIP0NKKlMgKbfotKxX+024nVr0UQdO9S9/Hi4EnWtfgi0iECs
1OgVc/HMGXHZaPP65G8E3kjx0wmwR3zfbXxMx5CdbUvU1mESWT71WP1BQWFHBe0Z0Y72uAz2cU8a
sfMmRtYOOjdlOTT9xtLacTVdXjN+ib8KQyLFSM2v7KSL2cA3hxNGc1353snLEsQo9A2rGD2c1oxM
s/XLzbPZoEKxEV2XxNcwBlFL1SXabjfD4JeVHZWdrt93BDoJtuRMComs9uV36hca1tR5JdSmJxK+
jiteD3I/Z4+L136hgW4lDYu2osTMPZ4X3ze0nm91KDdG1b4qDJ7sMpO0162hOeXwdjJTUi5SfdN1
bF6ay3HfStO8Xk85CKH1nYKenSZ76CBfa4LNru8oNzm88GmTgJSX1RnUwDhSc8+c+xu/SU4RNzqG
dZiCcJeuB6QZDJxyc351Ysh5H/k7R2NozklUUu5VUbb8S/WHVjYjbZ6u64zDRl8bDGrIDzNYenqE
edGZKYYRFcydNTxTzv3B9w57HaPABoNeLpl4fghq1nmv73VaZSvwBDi2DlhkTa4+5hRr1MwgEmOw
WAuaIYgzIgnEZAEKtXzpGwIHSd6P5W1SYl8p4ZEHB35PmqyIQUzpOXZh+yVlWMERCtjC0N0jG5jp
sgU9q+UL2o5rkrSdEV7XXf4Yu+R9ZggaqA5qICs5L0y2u0+LcqQ4wbEnfrEMDMducZkK0vkHm/cY
Xz82lj+CMwGraiKwoqK629W60myWdcLkzi4TeVy17RC4aELK+HyzyvpTF/qei8UDGXfVM3IvmZcN
awyJOOsw3x2sJ0y+R/jQrgua1sd46K5Xlah9G7YRdxeoOSYfpdvF192wJqxt4a4s39HjsDf+5trT
bcHNiqA1elGtuXcxq/9FKxyJ82EJXvblWxjgrHCNmZ+Dmmc1Grv07E2WjT3Ab1+Iyvc9aoIBNUXC
i9UXPH9fLfCpyK0wU/Bsq4JewhVtUZTFdtzEMZLi04RfcfCHmKMxIuUfEMAZ9iGu3qtacPgY81L0
73vJCtqgy6+GHwRSwceoCMLeZw2EMayo109ULgQt4liEMPbHzyRS2IRBSFBfusKWdrCzf25Nqq4a
3fSldr5sFE4hsi8L/0AWdzuLtCNHiIeQEbgUn2JjptJ3IuWOqMtAE47nliGDdTXPwWEoHlpK3hI6
DtZYbnBT2cBvK6B6VlCOvR5XFS0+1sWSjBrQPAQ6v7dGRIPWbN0Ol0CFYk4vlJXa+qSl5HCXlm4f
jZmVtooB4MBrAT+zZaziypPphOpMVaCVEc1YNc7lQTZ6wH/0AMgwssWm1PytMFYr/54QQygN+ZO0
1Cn1scBuZf4mQeHUM2m1ga+l1MqPznoONIdSH2xsL2Ig5Ugt9OxaT4HNlObIrnzuEMalxX1hb2GR
Mdb0YQD6ef4tbGVtvMuXRLg2CH7UWzkdMCRVr9fPBhLLAxeQhi6Y4MW+3PAApSoijgUlH+aQdI0y
qUZ6bFWiJ4RBUyMGI+IlQyS3tAEyd2HLU1py38wxDSGdniVDyrhSrr1ytmrxOb+pJoY0Y6RwFpFZ
5lNykjtZJhjKfwwoRRSecRGV2NR6WZOEivp75yeSouNFGqKParEpsKBi9Aa4hogOw3J50Fow5vdT
Q8NkM9Pccd527Hghwtmt0OYI51HqKUIh/UXmImLbcvQ0mpvZrAbPEVUCVIBLARtLpWIEkizE2xfo
+JQyXa8xS36jkEDh2YNs4/MFWwm7D8lw5fOhx/Jemgra5pU0DZfoBvK7byjX3kvRJcRw8GOh4Lyq
9wB9m2ndHEKkKIEpoaKDwqXCKavp7TpX1OWh8EWTnYWV/p8yHyMPc3wE43waoSXJwSbcUcEyycP3
H0tKBDCj4/Did06fSICwRQVa2ocJBv3gbHPZCph+J58Rdp95dQ==
`protect end_protected

