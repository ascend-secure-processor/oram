

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DElyVbHQlTD5myh21Z3j0wNJjFws5VTNrbLUSiUWSZ/24AuNXPddyVhrNaf7MK7EugGGDtralqL+
I2keUnk4ow==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BiF4dEhTrLHF2+c7GyyiYcOTeB9gPtdqzD5DxutghpwsSOJkHRjfqEI53B/sawH51BQCtdB++BYH
szhuLEY5WzncVr7+Wkr25EXgjmxmpd5jKke2fVDnRZuByZ3JAEPUL3fJ2h98qf51Puk56aF/NZqT
CZJA4SJY2QA8W8IGFM4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RoTyYQ5v+NXtIH2b2hxjDMrVxrSHy9UWw5oV4DkV97OWXAYXp3meNfg3aQPcXl9bijTfVtLjnnE+
NMxxW5qG9Kz46RNp0VB1GePzw0EEd40gs1/jtUnzbboxuO9T+RsDaCf2ARHrBi/vfNl9rQz/p0ja
5fTq+kb9sJoUSMj2eYwwPZlaxh9r+VMiPKMvkV6hHfVfv90nBdOuCxMFrv5APpk/GJizzcZYJb8v
6fXcMmx5GRJlQYMS+qfNqSlAU9bqhSQQ41dsm5QjK98AvAMg8pQZejFnk8jqIVtczNTZjaX9jveb
CAJs1ryT7uzIuApzavFdq4OLCz8oJZMWJSpVfA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NzeRMU24aT1OhFv95ixQFsHHDn/w//Ibpm31c39gZU5dYWGBi9hxwkZQW2aT7XjmgSLpg/bBa3wj
unJLGUk69tp3IKk8mm3Pvn3if1FXI0FHvkse4UHuy99XJaqGfEfjEi5HCtocf2yfkVbww8Bj+hcu
sQosFSCVqJ/FLrJqd4w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y/EvVqMDh29OZYmRAeNF8+hvNMppRl6sjVlutqRXsE7X2XR/NYAfEvOeMd/QNBQSVZHteBi9VdiK
+Qy2ga9gGb1ju/PvnRYVajMbeYbUo805VslSTHul/cKVHa2GmXgpy13DM+SYdCpD3IDPmap3CWZ9
Ji+89z3C4f91uiqdql1LgwIxssLzFj6/8f/bAlK/d2rDT0hkMICQvHPb/mqjxgGKxpGYL60XHAFW
oMFVCmCa4I526vOnCcCRYF8J1q3jFvyU+jabTHwkm7eBTeeG+tqmF2fKKlPG0HYcDzz+outrSDlR
mO3uApFJWrNEK88FHiXcvOl243F2FN693XqW/w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25312)
`protect data_block
4c0m3fsjfJ3f3wUTcb4uXgD9XtslsyQCqpyk2V1ObHgsVAOgt7U/md6iev/M7sRb3xDNroktoR74
luLkZOS4iS/327ScrvVP98rhcnTKou7r4/0B28dOfLykkodEFJHz3YmeoSOhRkotyb4fQk3skRbp
6YIC1TmJSdjCKbyTar0iGflnXxYOrQvb8QJH4O9O4swXkVrp8xjcP72oVsqTISRaimCwqZV2i/Hb
RhuU5InpljVW8Puiy2Ge1Q9bZWSP3n14qjjIENetaY3r+5Hu66NndwakoOad9vs093J5QoTXUJlQ
71popXZ9vlfl3u/eLZRPgqRj+pzxZtcEAq/emSkjI1SXVjyf92xFi6zrTaY6BXBB2kdv88I9ZTeN
CbwqNPMZK9L3V7L/wIRv83tocSODpicYlpxqQp/3jcLiC1xmGki511gpfPcIGJ9XcpvIpHo9FHcZ
LPwZ55FlgMON8mu4cYqZ7BLGIPLu3oh5LPhCdtqup4ZNQGtI2si3j2wBdw+WTRxJRbqMEhGvupDO
bcs+zc0F6Y9FUO/Jcfr/XdonzUSqJ9gh5y3d1sOP+B2NYq1k84u0hiZxN7OnlpN4EVvbgzjPbivV
RPP79u8IozwyBMe+tWGjuCUMWDpzJEKHRBrd7+xhr2tfFh3z2vk/2M4viRr4gBMh39EVXXukF52v
8XxEmGvVd+qRFPQD9gEtJGXKVlwFr3fdXUyDsm/4zjoxRRrPbGTiT9hZzRfnC143s4fF0fGZwlYP
7WEhPD4Y+uJSqxoILjCDw691KLVK4zxveryrYLVnGOTIlfw55CzGYhnBaxXoCPmMF5+M3bNno9F6
H8njHakyr2iZ+idaNNoPQd16C2De9Iik/wq811/JsyJB+bdRg5jvShGJ0brXaAw/ENb8I5BGzmEk
968DXygaKoOFtt0wcBJL9DZNPiDwDby+fNBJXbukq3gixXeFP7sGSnmW6TOirU+wXDZn/S8JdiYP
M26Dg3uf1i9NWYnWR77bu7+Kgnigvau6evtckFua2RZLPzMuASaQJjZyb1qedTmG7d4d1mHhzDsT
AKmj7IJGHN7Vtu51WkSblR2ZdgUIGP9g8vNmxALnjwco0d3MWkcIcTAv1XNsBZXWVjjfxWxYHZYj
S6Y91qjmvDQNWT3KyCPxKKnWqIm5hSkX2PMTKfBgZg4jumEcxZXg1Tebi5kuHpTwRlOKy7isip1j
SCR+XHASmGh9NUoqD8/4PgX+4yz5giRjBJplhbKT1Yu87aN4mOxS/VeCDEUDOpOYQI+Q1SoOgKKu
zbdSiRLrDpHj+YQsd7HZlwg7zk35L5kHGfSGHvu+Si5V2iTU+xLA3zPR23Xn/VqYvJODoVcJi6dj
U/KaX3kowEzUYbY33JZkehdnwQk7QzSTPQWcTom50iqDT5tsoiMdVY4CPNObMMzrktpTa8LTj0Em
nbv1l9l3576BOIdnf8/ZpIxu4rviI8K/gBr2i49JdhHciilVYPnTGyFwqtSTVzGAg0uy3a/+ZOZf
rYjBl162GpvMI5Ho0pgVLR6+iMPPEOnzKSE3R3tJN/eygYK9DauHXr7+jCVcMp4vnHff0Ai1Mt6r
nR1oZJBBZbhKr1GZL3fWaJtwgGPMzjW8jFruvqQVSYuA+J9GZAVY8z7rAyJ12Md5wiwhaHexZiLN
hYscIrztQKc8GfOOkgDppFw0xebAjwMqSn5gCdJI86tb0r3xSeNlV0/QNNsNSFAXwVvdVj2gyUJv
3IlncYPUE6H5oGRfgzab65D1aeqMdod2ggngRZQsLungJ8m1NNK+q/ik5lM3oHFhjaasyAmhj1Ij
8iv7g9Ja2WE3i1B/EgW2LpNLVX2tbbJDe7FG+bNbmPNopzozvT0ZuLmiSdtGCEuxsUieU3ag1Bmj
KFOHU734iemu1cvxPlYmzSXAARmCf3t1kuOMzAMcFeymPnPHc5zqIR73prEXEMyUIWrEO57dDTni
aMJ47LfWBREg5nadipIwN9fQgFGYSJR5f+peM/PRHLJMq0eP7NUmLUP7NQBOvqP6/g7+j6PjHn0p
kQQER72PPfrzhE/eMOrzQms5WOgERaM1rcRQIAd72mLj4DBmd8S65vYIHzlRltt4lkG/7coaSeYY
qZbWiJieKZz3c0ztEXJht5otLp/Immg8ORrdOC7hWDRZPY+SQSwczj1PQ8kIA5zy69imtWVzXEnD
ykibrM7i2NSU9i8jxG70K32xMPPN0Ym6dGIJHzRIEYXWFxOIDsCux614ldr2e3HpUJqE74mCwh98
EhmUpSltR9+7gGe0Vdy+JFcj0FhIK3n8P5jMXP0UuE29IzlmTPsMY2krYanfWNR+aEqideQiC34l
+OHyxtvHuIXzfEAsBOUkzFOXE0YIMQ5QHguGvM+sWLlfB3+2k6JuCBnA81hNwb+1ZGH4kc7CIYNu
H/nDB/WHAp+VmgCnmkYG1Sn6vrp+VZp90lPzXS48vZQsdVCUFFbRcpK3hpmfBwUXYX1cJogFKeHj
1ZCKQDbNfUnfoBTQtehbviI+w0Qlogtl8pcrfR8KcnW1zJg2xpJUsBGeEzPE3dGeEww3AZyuxqH2
40GlNbNuaArxCkNAb6nm3TTLvgcaBp6RpfRVgnHnvzTVb+pzHLX28QqxSX+K9wYY8xMnbGBSQsrA
4n6/TlJEKy95bBsr3RoaXQ3SQySVCc/hywcvIfpDuTsiiJqZt/LLABbNvlgvCmAzo1najL95B92W
/5Hm8YWmMYap8KTX++TPGRqAVwyRUsTR0PeobcDN6R4cwxw7HdVNSpeJDvLGr9UC3qGEds7bQOEB
dvUbte/SDoIppvjX0pFbjghVQTBLXSejhXL3G81TD2qLoy9MwQj2FeT18CFzgvNmMjFikXWIsG17
9hKo0WDqQ58uN6Dc9EmdyUiP4vXKgHecpiV932UPvxTF1rFoOFwkfVFC/+LYPhWQ9Mu5I2UEIzRF
FHk+G/SCkWnQ/Wkbsr5c6lo4RpWy07FXZ1Jqr6n/WwFTYtCq3gmUDtxZsRoBOV6V85UfuBZDot9+
qq2Bb9GqNNIxxOCRhtoO4psa6JbD3yQRCygRrFdi20Lr84pmx/4vy/bx0lOWFl3pWw5iId8wllj1
RxYxq3RoEbimVgG49fUjygprhVlgcVP9s2rQCQSzifZ13Snei/9qe1TeLqTYgKpGSI9ID0fs6Q9V
BgzluxM2uSOYhxr3WTHgg1FF6if2xOe1a9HbeFIAQbjCFEDaHgSFN8X7yYGLQN1hMdRbVfrG1NJ4
xK9gn7RCy7eEVzLpcxbtY2wlpvDGzEy2fm2LaIl9KWkh2VbuMfA39iGPvw0jpzB5KKKdc48ThDwN
X54TWK2ihJKJsLznnpmwJX3JHWGMnvYyJlt3o8MH9bftxuX+GLaeT+zEjLZcAkrauDIhH5YIRMTh
kNofkd8Eg0FrZIKY5NSd3TtNlP0PH8bdJgApworALQedZJfwYLtW2j9KmamhTxrsc7Vi/7/ZhIGe
MoMwRZ5Ekgv9MYj8GdI/BUMYpMguPVfjeOi+av/6SdJs2Dfm9pQulvcuZj566UebD39eYZYPLIRX
69/kp2h9PKnq7e6/8a9iqnfoAhSIpOLnCT6b3IFHmSV45oD97RWcmAZLDxEs452nbpLpVEIpmP9o
prNQ3rNwMhFkAYJt2B8wmSrPnY+TILcxbN5/M2PRpxd1LPmeDQjhmXUbVbudz+Se56+mswWZIjz/
TqvdrilWdp6Ls4dDul2hdKRLlc4a+9bKNBwfKgXcMJjnMfudHe2FIP8ti1xM2bDVkaY1bSEIbH8x
Fp8LxRiofNQny8WeJe1ipKq2FRaUqvpOcH5Q3yi/dFnabmKfUn/fR+B12+KxLvR4m5GlG764oXzI
iiswACeN+T6WcJVyGIpVN14f6rwv6V9RAFeMoOBdOHtAX89ayPxK3DUKZsj8qAPHJ+swkuWxNzrT
vECxGHibYZDkran3A0+olgzt0aryt1/76q8YhDmF5lTMkAO41quh5W12hhiDB9St/6t/fNkz01SH
57Uwvr1Ty7Hk+ANkT6LVf6XEoUdD7YgU6t0v+8QTy+D8yI6cfi1ImOVbryDTpJFVKRDwWGYSfHA0
2a1N457CYKb29bkfJVzCU5SEgI80GHQ2kiryL1pdyNFWS0ZtAqWTxztsQA9EqWW48hx1xnJhr6LH
kxY/ClZRAXWNxfwVq/bqcv68HE5PVc4xceYnGwJzPTL/S/goxZx9UdfDHj3qc16qy7ok6b7wibLS
5Y7nCAfnSLpsgDvR8MvpK27Y5bIHsUSuj3EgLute7JOo8c7Xz0nTjGuyaDH+gAaIFavI7DfMpTpp
cSrQXy3NVtJoaFeA/4m08t692sCdDr5fCtpkfEeLzAIzMKe+UrXwVkj1SwZTL8NONMYpE5YQkqev
UdJxgvq8lEqmNRK5PbHtuBNzPlqS1g7rp/WmilkNpw8Y+vykp3VdTayujsS+Zaz0Clq3E2Mcoqxe
C7vZlX4p4yed/1Fo4Ly4jM1J2Y9W4vMYEZgf8/LbyTS5QfPouuDjR25BuuGcdRlq3yTnIXFr7kv0
iQBahdHRFq2RV3ObnXqXydg3UwJKS/ksMmHAkDLG7z4VQ0LVoLtOVM1uY37DXtVRg70ARY6CP/1R
quvEmh8SkXif/whbhrCAqZ2w2y2nZY88MV9vEEijUbCZIQGo27CCIXyDIzIFfNamJAomo+QuDd90
IniqWhVNLP71PTT8d6EofsESEepb1coVVlwC0nvjLBlO4M55D8ZCGZj2ybPqWAC24iS5CiQA2nmp
FFrwJnKaeiBeI+QJ84Ml2HDqG/MVsyUD/tZsiiYWxK9khOgzWRh7p1b9gJ5E8c1+QAdXy3Y82mVN
Cdih0rgXpE/CkPELCvje3q2gXkyRha9UYG+XrWb3AfZza51wHp2bDE54rzStjnGHd2DT+sBE4bP8
Yo9i0eZzCuMftZ/T+umr6JeyABWt76JIV0RjnAowq5rKWJHxG1o/rfoLelP1gwg9EZVFbUVTCm4n
XB+uO+oCXYsesSruEpvFqNntTJLV8PXuvEzXKtcjfomzk7J7NahiyMRuVnFI13mnRKxa5tb6RQW5
5Mt7Hi1nq3hovZD7WDYveGDEUV5piVKBR4A81Dg8VxcnXc/jnyT2FIf2aNJ2tSFFGT1j50npvC0D
9HkkF+ABfyxJ7o0ATmHut9H8avVOQia/xmk8OKAFDHBR7EO1uECDVkSPnImfz0e2iO7y6f6d5yU0
j5J695m6W5mL/elYuSjX603aOE9aqPYnRKuUZtcdtfiN7kdnnhE6Ny/SlxELe85P9EPQYQQg8evf
F+EiqXSPimTY2HS07HaR3gTvoXElxPblKS2jMgxcVDm153o/rg0nR+c5Xk4fD0VUKFf3QiEjUoxH
gwb3xqYNtxLQ8eOHx0lrPsNndwCQB7UoyIO5s4kGf8UrEpfacSx0WxnYNyh2z8/d3xACtmu9zeYk
iiCRzjVOVrLxM3YvQXvDFT2kRfeuJBej3extD26Bx1rGeoOlVcLZnpzBqpm5KYaKjVifL6E2SHOP
Z/CFTJKMknhCZ2F+CV7XJnj8yex8MWmNlJx2zEuSftkAWPFqHSGg606Y9ricaLEcdUjlbhm/PC6G
KOYgNzkIHkE4wZbBxYHLq058xr5ypK94vPRAeviQ/dxMuy3/19iYLdGEDLE5+FRh9ShA64QU8MD+
TDSJz0rXSI0LyvkEYJbJU1DO5ac3IppIwO8fS5xQagLc4FbBsjGrdiBG43HYCl9WGFvxCLb03tvP
6rrgDTKzeRQVhL2X4xmqd9YLtKGIQ4cXhUHS2P8GzPBES77E6xc213+q5mpOA8D0Rjxlf0gJM3ES
o8C3h9Cr33ZPsFcBY3JQ+mCymhO3Sp7Naun8ROtL94rt4pk8dPmfsjqGqYKN81fS61zyk1OtO0rd
BD4MdCp2Ym03maVCRanwfIFS4OCsJDAPc/RSEozzWzYCmwvV8ofjDHZnNAiZIJSVcwnJvKubJWSk
I8kaxUBqB9CvWkF/HWlIifcmw2kwv3XxcmAHmHizB1GWCPh7BPduRuemKRMy9gKeGiIPtEHlOBwR
fvT5o+5XAE/1WCop9geGNEXgt3BOXmtofg4bAZiNktzD4ZAyXLthGtFONvAo2dnXP2GNQCjmUV0N
XVh8bnWRZjjjxKrosmGFNaaVjXsV2aE6k8VkOKWRXNFFiioQnJyUO1Rdnf0t3fSCRVnmMjZYi/Q3
1OpAVVRIzmmf0lBz1hmdp2fAHHgRae8K2dTBLkyn3/zbl2O5AyZBS6wNkhgxQnGOAJHxLnYivgy4
MeBfSY+YfumPXRZa+r+zFThFrO7UhTj0W3/Lv4aQSA2Ud5uAqOHaXht4foVJdYz4J6elWyDNzjtM
vEH5CzReOpvz+svYDduWRQZ3BmdZS1WPNDUsHchXic2MENSxebDKaG9K5Q7mQokYvP+2SfouMnjS
VI2LDaAPws2VrvPsqR1mzlTATk6JEquD6NlHeLYPAMUJ0JZ3qpAvmRwYcOXjEr2JKDadr7QhU0rs
fcPCHD10nmzNZh4PYTc/T2AEkXT2uvJQdO6Jv2qTnpOFCJsvrMcNWegWUggUQEOxhvuZpxpDjnDt
NvvVebMpBexTVeX9Yzh2z3+kGxDUPVZYCsdQMgGoczxS5DehX9HaJwpIIQJR5VFfxu/SGvM4RRKD
4r7B5OjY6bxtT3y4K8Y2Y6C/LI2UOILmA8SptcpX1YH2FcKel7SKZjaVZjjhrUwoExi9uYLfaAXs
DF/ApykQoR2TjCyj4pcl0okQ/r211Ufsyc4XTrKTBiE5vb2KZdHtSxdwe9iH1vWxvlzNiSSjMOq3
d6izdp8fBoGSEKNO3tJTv0SMTklYHctVUhWdBaC2F0A0Z+9+b+KBlC0168WEhukNt90Uq/Cc/jao
znUinEy4kOoIIOfgT0WuaAICmdgBvx1GmywXbCwTDk7ZsbadIslTNfqgELNlMBrUCGSXLwVKoRBQ
JiT/eswHJsccUksGJFBP5yo9/8f9iTz/4uxq7vnDv+dunbHrcGTTSqzjwXN52Ecik5v1iMfpGGtc
kwg8RyfKJZqn1lyTJReroHGb9DYDbujMiGq/zUtpDWn1szwFj0kWruo3D/wcsz0mTpDKI7j0ZToW
q4mjnJNvi8ZwUVnn8IyxOs4oOHW3k9kQjS3g1ZfqB/eHEr6ZrUDY7dW9CZ3DaIA8VEPT9K0DfI04
I2nj0+l8bqb83Roqzw/TfPhbgQfloUx9Dzwokmjp0rLCc0RakWngkuoOu+wmLcPWuqyEiwjfwln0
PvNOlRZhFLNh3kNXLkvp4wjCAxqubs/TJowHdBTRAwxP69n73lZigan2HO23UBiorj3VK19mmhkP
3R/PEQd4isqBbuVVFWPhcixtb0bdopBhs5HUkCWqTS7x5UHA7wMBlepuQoZ9UMUmmL4QSfgAv9jj
4p0WugiCmMa8MU8VZB/vl5YjFvnUSnSfJZMVk2Vs6YibcqUxjQZy7pjYfWA6/UL0wnMQt8iJPr4r
pnI0Iwe4feSKWf2nrvAfW2qp24+NotbNuX2M2bnPhJYUwGWbgasaJc3G+iW1NgwOQre+m4t5crRv
qgZI4ocETYwL++mywfjZ2p4dxr/Co5uIHUN/8dxoQVyQlrGGX4ODHtLdQu/QlcC1R/uHPptHI8BH
BhZr91lbvkHvjX4qP2LXYBdgDVUteCqF3yTjEBmlvFksatQN3I8hHsQJjSGEoZXQE6qjVyMouffa
MGbeemdHDMG46w4phnoHgxkXCwlrazkEmJewHGkPh9/4z2LtcU9KroqFCpebRmsqx+gLGPWfZIbJ
UD/H+4ebkZvSZoQiDx9rxJGI5GNnMzCfalL0lLahBIFKFOOw5vJ/awjtbbtTHAcbnJNIIfqdm6Ed
8q2Iku6UHefzULUyGoZpVj29jdQGNDATAhOXY4xLh7bNjUFCMB/66YbUn1oeIg5eF0p/QyyqhDlK
udR81oohdfOpnChcBFliYXPDpipkpIRtfdVBrLEQ8v4AWR1WhDYF/3I1H1DVhi+k2YB6cI6T8uW7
6zb8KFG4zkIycfOF079uqVddbjeNjYPXzpBr+a/AxJ0snzvHGon2KV2zR0+G+Uhhlj4SzD1fMlUh
p2/ZuYmm62iwa2/mkD0CIlNerBU1tYRuBd5M263Hd7NONIxMdDExpftr8lbJf1Fpjcazhw2ZljT0
A2d6zc2A9Phyl1JVwDTO6h5UG+blbgYn/s+2DYgmb9Q9a8LNGl2fC1pHqxly9T8U1uv21JhY3gyF
BO1siJ3kTY0S2lmEUZHm5B4LqkhIJrm0NBBHmi3eFAaiyc2EYaQd10pnvQndcffk9+TpVsF07uuB
oKuRQHlAUaOGJbxtKAUcrY9kd78W/7AjwJ/shwdjWMpnt+FY3qFM8D8wupgLtoOiaDzRvBS4x6tj
W6Utio6A0HZkz8A4qjB7MmS2o2xVf+VFq3bX1/Z6qrlWv02EYQTTY6mXPd0ZDuo9qlWkaVBypgnG
B9Mr8jalDaeO00m1BkJ13+DII72zehlJZs7Q3QEFvnEtvzbQg5DiIVh/IztIn90jSP62dIi8SOW2
lTk+G+rfBndwSgJ25DY8UDZgEtBYuWdfb+2rXx7iXNrks8PEsyRiwh3OdXsbHY2KJ6LL8yxa+YTV
5rJQnw9kFeyrWhOK53FTgcGZHqjuBoVles+xmTaHWS3H2RNwV/ArzcybNkuZR6xSH++mU+d+5cEu
L0XVQM54L44gQfOA2Zp1j87UI31lbEiebGtzeH0mnL4zOL60+LxC75XIDSEP9tdJTfHGkmPMvhw1
upKucxeXsU8cN3oSLvgcSMNcigrWzon4FYfX05cdAQ4RqwmxL+CPo4z8b4feo+WdiUbXvoxWQYKe
AhORcTPLsvyusWDM1ZUH0OX5men6zpHo11UzN6aD6Dd90q0K1DV5r5xJfZ2hRPUZXAkOgfZaBUsq
K0FDwcx1lsvOS/pInv13eO75rfwlk1f4CFnEeSu1TXCuPxqQssIAP/JTdAw6OmVkMGYRbC3CNIli
elWN2VjwA4KA4EYLr+iSO2D7wlLNMyXPxpBxB3d896sJ3kFN3eNVK5eu7re0d0PbEV4mhrNp2mT7
6Ng0TfmkE9axqBK8F5aYGT9qTNrbtLxAJXXNKUikAO2tpo7JhYsWlZvVRyOk9NS2oflSjEcxYep3
93xRHh85Q/5pCHaq0Q7mli2cSiitH77818b1FdFBRY3hoKIjyu91EK7Rdyc7X4GLWXUx5F2rApqk
9W8V41XkIk0/G6aubiA7y0T1UEA42Wi6Gx4ZEfhk27Os8UZFetsDi49sW9CJ+vDcQLSUvHuCVwDx
SQwH3+m13IpO209Ng/WvTRRvM8vM6ouM+EwIJ/5J+3075VYNjpBVXxZZlS3GnHvQ516p2aH9F3Xa
1cXoV4/54i2VW+I6G/Z9IhhPj+ZZpWSXAGV3f+OLEHk26MdFF/6XNqSdGf6+ZuFMGKNxrQdowUnZ
i/X98HjdXRUyH759BAQ487Yj0gBio+4NaICEs+GzUpZFSRoA0JPdXgEDvgKCTyIbyQKiQ5lEqnO+
SRHFbByWnYpsVq9dkU+zqsh+Nx+TpCJFZ5WvuWPy/aDHVLntdnVZJfTHwW7LiAxIQfLzh1woXiyi
VwsjT9kuZAYvbH3CudX62fHEVCMyb6yMJ7SLgIs8cgVa1rs5A9w1UPSsdl2VumxfmhA0pvUJnfhU
qKeokg34A40wAmVv0BO/qggyT02Kn/9s4tCpZRxNQS8k8IIs/JUrmzbSdMKkAUjO7gNyjoZiPVTE
0KHhLecJuI5YPry1tU6CRxBaJAvCInza3cJOELagGqVqEVhhespOYrUQXfT9T4p9eQfPvH0FmxYR
4PS+M+MYbBUazQptVrkCQ5azu19o7bz+4V4wKhHFfgnGrNUYAz4jGapzt1C8lHQj/5x3sSYkIve1
cnAOf8+0oWwHHQCN9unFv7bQ3pFghih0H5EfuNdZzXl4qn2hS/HqesirG7yY2ysRgeaTcZb6u2lD
N5ND/TDZVyMEsN+LH5jnpI0yHrBGuHbCnBx1qUy7dAab5H+PwuTaK6Y1ZzIuW8HwPKU2ZDnyKyvc
4A2muDBnyB4hzZQKD+0q9csrI/O2hj8d70egpGCKITAgguYmCDyYT7rSKAoV/sQFT2kRgWHpkVtk
vLHc4AvLsWUN4QPKtu7NAjBSw3Foy8clw84vPQdiC+UyY9ajQERNuLagm1dzZKVLNcMQWLlNLWxQ
s2DYMJjSiYjNrVlnISoeKEjS98uT1HVnjlq+W5g6IMH8jFr2EaxTtR8ZIwXNnUnQKmfkCJRZWK8M
dOX5jC4O19IkUyMM82DVxQXL7mvA4cOmE7Rnpzr6SIivauyqVcxk1y9Ato5dciZeZykn+c5WYXep
X5az7sIjEWEyAE1kN+ADUOApivOJgDmFDbSdK5T1426W+slrfrQ5A+O82GKg5akvOuTsQ3RzkpPQ
D2PX6aVR0YzKtS0M0hj5ZHEBWUheUIWnkNUoW49kejNX8CtAbQAGQjL4xp0wyVi4qte+uDjzjaw5
qCAno3ydh6+UsETw7Mm/fcYraS1cXSQwKYYPZeQlXat8/cII8CXvA8nZ+iBlpKLY/zt9G3zhZdq5
ByGOUl2eOP/4t2/duM+4KE74hK3TS1guGdZB2gN5l8kgpdTPvs3cEyblxfSWl4PpkFB3+LIVYRht
JI9NRQO8uzHsnUxr+ZjgCv1oRM+2wEJUECAZWpObm6+T27p6/p5F/JLAUQmVxXgyyC5xrOQdGnYA
G+jkl9kSekXqVV8DQkyNX/d1HdvM+/A9GSzBjqFbdwHfnAh9R1u5Ihax/L9uV1NFjXfL0/6KEbQD
i8g55Cs8VzJ79OsvSyjjwW6Nbh/D8iEygRAW6qOWyoG91Hxlzom7rAMVpdUENefs9eEAoP7+FPIp
b8Fw3cPmSYiCHobqhrrAVQgHPn9AcvE563/lgi6E1a3TNPY1X9eBOE9omlYCM0u/Znfri4bLZ3YU
ag9KSHzbYCKHKp3S31GKsHDoHIF2Cxx+h5REVENluScHWOS5Nl3db8lZEWTAm23xzV1rSN0ijuxi
DbIhaawAFGtYg7F/f1Khn6T409VoPMiDMI+nmTiQEcPcJyeeCIdjplFYiIaF+kSq1aXYF8CwHZOD
5HMiPVvtfkLgyZN78iNVnRwKaxHiJNJdU12pRDmuo0LmQmvt0EvNo6vECiIxNYWoobqE7lNS4Rcn
kMeGBw7GjthxlDEbsetGOnRkY1dLnEWW3LFNiIFL4KbRZXFd8kgTdwyCLHAh0eDYfmiBiTzeWJfG
vnGOJpNMsA93/OcYr766sOFM+v9XMBViiWOGxfH6bgpbloRzK1UwCtW7yf+tQthafOdr1h1bvc5d
QGrIqd23FJqUBk6mxkwd7VrOLXirPWLkZ2fYuSo+VlVo87VVIvmT64vRKI64rPkS7/Opqz+ZrtXk
5uwl340+i2RyO0fmpC7aW2ASWpk2f5hXhcBJnzwfYYi2ilUhu9kUZQpAXbS5Q54iBkkoZ98bM6A9
Dg0mPyDbHOfJgc0yEfZjiaoVMtZMUjfcFeXQZnZx2O+6BDNRhoANpN0gJyHEjzL98sMXWrzCopg9
gT/ywOVOYtDK/cVBmkUOREPzyA0wCFG4dZvFEGIRG9KBwMwvPA4o+7uMqj+4G35jtKeUXkwmPHBL
v1fAf2+4kNU4PyKClLSTmBttebzpAvHjL2f6mvD6s0Bq9v1q7igTadxKtBURJyphNzIj1OmX4mtE
00GvByjswNtC/sRiciKddWO6iNIdb3UEVS+DlHrIrrG4dBQE85fHX7He5VG0dVUNNwnb0HyzGVzF
19vEN8qv1pD7YThrdK966wXbtb1ZPTK68FQ3xL2UdfeUqTlXwiSojG0My+q8ZVCdrBd0sMHg37UV
RVCpQGx+YKuotmIVXS5+cgzJoGhTvaoLHkOGZ575zFlJZ2GAX4Sb2xfGGR/ZV4NAs6wl18IFobH2
j7Q++dKOAXJ96LOQpo2EJ1f3IE887cTsTb0Z3TU9fwr1UAkXH1UFJX8U80ecKdL15YNZ0ykozBdE
IpLKnSRrHBzbmgzAO30Hf5iEQ5Mc7KT45CxwYnnkSeU7lUPuYRKPnohE/4tLL9Bf7qN/YmhB6bZ7
+nxk7JP9EG3c9jiVzUgZf6yEEpRMVRtX+21+cd0ISp2LXFUck4vbZLm23i/ukcM99PYkDsLVzW+C
IuOHEA8qBPCJMOHwPCoHY158bQV9nn5w/jkrdtl6TOQLA/9klA0GshsBZDub+EeU0ivrwA+nrHyZ
XLXPz/opGSIyzekeBn8MIhEM79DdO3/nsJY6lNgPhI5hkwwICITV1sZzdD0jgw4K+fQ4mlCZpJ34
f++1yBWBczQnOntfNSzSEl4De+XABNtF6uaiDCvclo9p3aEJLhb/5N3NGAUA8WTKJ+ebU/KC/h0j
EZK7HIjeEkVW041Si7qkWJ/rFz5h9v3MQE9rmE4c3N0OIjZ35ogjNkVE8X66jgOnsVOQvHk3LV1Z
oOW7jZ50ba6HslBMU8dSlwehVmHOpu7qhI6usYdjPpMVZTAYqpQIY8U+XIyBOgeyGEHZXnKlkjW0
T5LckkP6OMZLOxfdm5np6YyZHDObA5rqJHSB+NoKLrMK8Ha6e6bpvkYIR/PrOfDjdJVPORn5sj3j
O+TW4xXKTSOUFQFx+Q49lNQXgOdylMzX4EzsuRgRMbzUJm/+ehml9A4UFxwGO4U+/dmohL9CQg0N
bZBxrcCg4ksBZ6Mf5uvERfyyDo0fPpUZjCKF6XdZrDpSHI2/yGGo+VyzaU4U6xk3CtlefR/bC/Jc
Z9lLPqSJR21Kb9oQBVGKgCuVtD3bEwtzZgkitxN9tFtcEb0T3npZCRhZQAj9D9FLdODYeMlZWoVt
9vDvBxXyGRa0D/elgfxNkU9hqvFRv6p1y7zJ3NznrzwcQuPzNRzYeYCkHtOvRpIB29nQPBzNO/Hr
7XjTNhzMZey+KqxxsbllQ99vUvVPmImLSwzcePz56EcDIWWrZTThKwU0Tb2dHV4DwyH+Rfy/kACd
U5nPuLc07QPech+Jd31mGZJhV7tENZfxN/OJoJ1Es4ftH6NmH3iHhhmxZtvxQHA0u+BCtf6STb9q
94EfDiaFIHMwqcZOhC8FH83dDzxogUe/JlB18U96mYuQXcumaZmlcTDuv38VLprfcooLIiiN7QJe
TupJLYEFLsorcX/niTJ7DHBlzCnXm7PaKpX89553yJfuWIkbNs1PT8Q+FumoIxYt0R1TZ/PhS3da
PcrvtRPCvl6ySfvqPo0gVtXdbpHZvs9Z31WqZkBL7daTwT2tj5HnG8xBWnyths2yVYyK5BsPJMxP
2xrWXKgP2Rfz83IMdmHUnScXKYJM40zhphIArmqThprzTa9arIhfLiK3tUVcDg/GK+JG6fggr087
hjY5c+lV6hUJpswxIDcZ0byIW0nT/5IWjXjUxoJmsCULEhWJfNdeNLwBkc0iCGu4rJb92jkA90l/
z+IapOWopQdjJR97ArXWURndZ6UwlFZ62cDwt1zUUZpQ4Bm+KoceTlYC/9Iw7QjAojWemEhc22tx
tet/rv9qgDFb8b5uQ0fysOTYyQXv3KqzzhakKe7xTgZKIYpT8xEwEL2xqFeh4dR8znpVKC04XJgz
ELx+WRu0wLYHMsG2AM+UlC8isVgNQUREwi0GjPrqNuY1KZ95sDff0v0jAVkCSA1mVNub4n4KwboD
mIMbUhdPvcNE+DfhJ19Md0Y2phALMr8b1uI0KLZ9Se4s8hsG8FHDeyWJ4hbKdySQ+yxmFKJxm86N
U8xVon5oWj6nFibgD835zjGI5e9n1C8ZaeQAMkZnxwEdtUymhK+dQLFTD6LH0+ntG6BEFAFIjLkL
FeU4cwcXQvXica5RAunX67qq42i067DIZaF+c2LUKXYzy46ZfFcfbhs3fHTY+9dpesmNS1LDkRdU
cDaaz/7Q7M6pmk6yspps+l+z5trY1xHMcWeS4L00+7kfmNMvVV4vYai/uquS47rfXVCtKG++gic0
W9C7P11ezhnUrdyIGy5G1WU22ZV7IZG8Qq7jYfHMq9XeIDt82AvSPCTM6yJar38Y8qPP+yZMZ82v
cc/VxtHxdsvd3X9h0ro3lYgZ5AqXG1SIYZDTrFkY3nppuC/Giq6Jd0TEb2KbzNwG4ZqwagFL8M3W
m9nzrxlwBbjfvZgz1tEC7If3p2KOgl/5HAWUuyXwnwm/VGj7u2vbKmaJV4kDHlmENZCrMoJyNumX
ChjOUremL6nuaEAVAfkLb2/5HdbdaE3GrEbngHcQuUFQ7HchPT4m3tMSpY54ECgdSpvgwDu8GuYS
ljZSjFIoLrkT52Ug+ObOzO3wkZzjMcrN6vU137mqL2P2SjQPa/zJfCf1zt6XNp0j4m8n9VFJFXvQ
tGEfL8BiQxyNGmHyf0aGk94/1bqPPHHDpTW9x1R3/xrEj4p6J/apjzaRQErxIOAZiqWRVBvVkEg7
bo+MBKZTP0+qvgM+Gn7iv5gSb+M1ctFMD5+OVn7rhMTkQ3ynqweEbbQNLlHjxj1xaNhjkPk7dcuJ
1VWK8QI+ihZhYncXZbVO6C1tMuUBIS75j6EoHD1hRpWfB1gQj//ZFjx8mf+sGT1qA+2+CgBXn1mQ
T9SJZVaO9y7aBNMral6diXkg8Mj/HG4+wEvwtFT68oFwc9r27HHTsBQz87bJwCpQ/xQNxM9JHfpm
v68OXKTMZrnTPMgyxJq49zO6JHtKWofnPTUjBhBdEOfE6mWa4VWZpmzWCNyr0kZoIK1RZcRgv8Z0
gHdtbb1zHnka8zfDEJbtMVt4kXt+9i6Mez6hkBeVh+iQf5S//LHJxR+fdG59E+148+LbIZ19nz5h
M9TWkYbCqY2O0R8ZXDRhIkWDTRLwyLM0ZOmdGNHOKCh2owlpJtkTkO+mQh8CSouA24ZARo4Zw2ag
7+bn76DDkqoikuF34+boaEmK/ZGec797EbS9GnzKDKJlP+tR1mrCKcPwhARiKg5lUUxYsTHC2vv+
V/E1WJS1ru1Ur89hzLCh6Avl1CUJgLOCQGYDtqg4fsmKMCw4nkz/Ah4xJvbc/FGcj8uF6ocw02gD
zKddsUUhW3vuc7iW6lgg/KGJI+JAjS5CCIfaqpF2yRBplQEdoU0eMWHC/iMhZ6iCCOfDq4+F+dRc
CYxH+aX5m/ZKDD5Y8bIpsizAttEQ2rH6UyO8o99anAC/zbf6D1wUDGyxIVvAa5w5hTmunou9Btkq
olTPlXMXCSpfN8mGgXvFpvxzbFD4LQkHxOrhChXBXwA+39+vRa0/h5SRRqx9OvoGR2m5BPimhjkd
EqNtW9kizU+36y0RioCsdqZOGP2y83X5KSeibtx8yhQMPsMpZlKkDZrgccMfAJufQEKF7iSgCr88
DSZ/+NwHrmcpQIPOdLHmZ8YHt7LcGbZqXBLNAJ4n5+KMUHlI3bX3NnBkBKw4XcvdrWFHhRUxptUc
TaELLl8c6ydHdGnNZWsUiWbY5RNm6+ni6B3dXhXQGyE1nEWmF76P27B0SvxauKqaLJsO9rr445mW
0bTxeVfjJ6+Qs6aoADPdVrxMAWkfDWc57+4jQETBzHMiz9lcm+V6Ybi+WXoQ932iMGsR9JxMsUO+
jMjrOyQ+wVxQgNC8dwa4hZK23OXfxyLhEsVOHfw/jn2951IuUih0OJkAJeTQxmsM+vbJZLPi1XTr
RvxOlrBY06Ek/NEpvRnoI7vhQazlxZhj/TQpMSG7QTQ/7l4RtGOKEofK9m9wfrBe3QCCkQSN/h43
WLLufa/AUPsPUZXDsVI3MBUsSrgNQlGadBxMx/kTJ/KWNcKEirYE5xcqcEr63sDrYiW3WnjKZ9KC
AuBKz6UEX/BmZjmV4gi2JzSL9YpJFXLj0nVTfUITRP17F086J/GXGaHkLG2vRMzLsVFdwV7zErV/
ZVguIhcMnmRDZxya4qr3/1AfzaKlNe9YNRMak0CpHBfI8wiAls+OxpE3ajuOhJPbfO9OxSeFfAYI
j3/LpfhPYukW0EvJsBn/JOEojsAxsML7dGz3ZV0iOtfwmrP7Wn5ZN5VzCptRSXPqHb4IIQTVFMDA
RPSoYZco5Le/HGF4tmvYeVYdpNGbaJ4EBu0d7IqrcQBPJBSSFCMJO8gMyra0U5QLcI8CPrr/VIzd
Hjg7gx7NylmR0aFlwhWGcq03f/aTkvjXxs5JO002VOP/fNPt+JN04PmjbrsnycWf5WDGdp3F4gb5
LQHYt/SberaF++I6Hv/So940tE4a2sw1UoJ0esaPI4l3Pvj7QHp5PdityQA6sB+0qVWyqg/snXQi
VEfkwzU6khczsEUtQIrZCUwfogA4TMciS42C2rTZz8QMQ1mDQ6NMkKRBLicMusumQ3j41iKyqj/6
/Hod3xK9yidOM7qaSEd+bbTR+3XSSc3APK3RbqtUtvp/X3ZFkkK7ZwFQWh3oHIjm37/cbFltGbML
4wcNuMcmuiYCbEH0a9e7HgkbGRAr/AigAXyk7SzHBlpRuultgNy2u+jI0R4n9OJdK+ye0ka4Bt4g
Q56TFSGBr2XAgPOkCkvwGPaI1h4IPhqWhrkYR9uDs7nasKdrZ2CtvuCJ1DgwpjewiLh/xvc7M3rp
NwJ3hBPD752D3KcD9TxVfAWtQYFoVNlK2giGYY/gXHwF46lQqzqerGF9WlypEwJBYy3bYRLS9rfe
jcsyanONR+JHUdjosVe45CH8TsO4qFzFBHBrYb15HAoeclV6DHn02F2+bRp2io0M9bz39kSClqdl
MMDkCLu7eMR16Rlwu+LQSKZKSvMidPbjx/LQXpl8fo/AmPf+UN7Scfpf0GHaRLEFXB6zZdtUaBXe
9j9hERs/D5pAw5HoToOup1uAByNuGoud65QP160MWpfVtqtCD5K+9mipi2eRNjcikjrZHmUpzXct
x7EFtqRI5opsf84p/uB7L99i2pVArSmrK7NiljFsunOjxVm+CfED7rXzR/FxHx/5uAuabw2dik24
CnmjsE+qUA8M/80srnyGCGMsaJNaAuyLuuaKGQy1GPcLONBp6bxrS65o3qnDQjCu7lhrQo0+ilPX
rPFjw31CbGyF+d7T7E2KAevNtHm5Saz6OEkGu0qGcUk23kWcNs+YjZJ2iClQHPosXb0Zs5U48A1s
enRf1UAyL+xT4hLSSnYqxKQsVob/ObrB69iXMP0eOJ5mrutzDqQAO++ZwaZyJ7VDjLa2F7GXwnxs
f6J0FNdHZIQ5XoVzwoOIez0wbcizLE2Ge7VjsN06YGSDwZ2ziNovpKMLy4ZbG9aJg3N6Bu10U3JA
rVATNTtXdiKSaXcKWx2XyWBAVaTQx1vr5QPFk/yYIpNxeTo1FXLt+IyiXWgPl4FDlfxA3YgRCIJc
tgSlUJXt6FxeJ47HuC/ENNyUYrbXzCVVS8m9BNXqlq4gXG9LEXaTgNb9f0Zf8+BEMNJvZTmDEk6A
GXkkVrO7f4nwq08yBme9OegaFahtCcgz04DW3+Mb7XB07VC32VyL4FNO6pJW2HGdXRRp4/hxV3/J
WNQpcCX1MVKugVcasECGBdkB8x1dmBvIu+/l3hHDP1rBCvUTqzW8QxHzNGOP+fHfDb2+hEwCObyJ
DrfOLeemxbl5TWZA4nFNSahaSpgnN1V8IolSqm70ofm62woF77RtWdA+h+Uui8Kl4hcC1dY61c9Q
4v/f/i/C6JrtL7pUxFH7wQlaeZO+desoHexFiH7CY0+lBc9eDIjhvYYqp/oxhNOAMP51s99ugQrA
RD3Ev9aV6dKliTaeM0eAtxA0KwPXtsv7BDWb3SpK+fMfFVSPZe4DRAghIk0r7TLo1EEbclYiLGq0
D0F6xLRkZk23bHCf5MncyZ7MduWAey1Yla3jw4j5c61S3MxldQG0giNSjSIXSTTHtt1OzWpIZ+V6
LOMs2cRuUg292fNyUg+3sW5tQtV2pqw+r/EA0mxq9d+VIdPYMy2ITmWLaueMF5HU7KH+nl7B155b
Ai7ASdPNypZAGMAVBlrO3PFnEC4/1eneP42v7Ki7UHgnhbMBKRJhKo2WfH6lItI3HuJMLiNKgV2l
v7fbpp3dTBeiNs9K0ps2/ZONq9Jb0oi9Ayz6ZNt/0pmJpCi+lii0wTcEITT+aunIrFeOcAgXVtmI
jM8A+RLI52EmNv1Q+suxOQEdmZCpVs9EiXu89PMcnz2iQAKpECh0z6DESznktiE4qguAg80C7f8Q
NBE0REezVhZIRLI/ieC5i38N4pyMNi1aaiiGQwD5neBVuiZFQ8ChTM1olezZscxEjVbk0ApkJ1uE
N8+3++cacZ/s2kR5UHu9ZZp7SCe9XmLAUYBP2HtDO0yDMeUQ/bRycVdbipvSWHWZFNoWTB6+Ng/x
xmFOETXVIWrgZcMoxuUeGmz+VTgLjbKtmz6ravLCLk1VNFD4biMWJiD4m2V4mqafnCSDFrFNPq1J
jOAlPpIR+nh+0tezkWNLffzaXE9NY95zCoKn9Bu47qwoD/5w+LBqrGA97DBCFBygOEaI2+oEKHhD
4p+0VX23bhzhjkAlNVMAsNOI9bQTnwb76LPP+QOU7McJc4DsrMqEQzQNWkEUqIQTThUvdfIyBAjd
VKuz9YcDdM08iZNasK7jjP4UDRtdI7fhIUe0n+PLh0mj0FCq4Ez1gShmbzNEp3d+svI6qS4BxBtD
M9GqT0T5QMhK3T019eRYq935CHBRDEvnouqkcFV3lGgaWGPCxDgZ9Mx0UCXdVoZ73+ea5F1w69bX
CaInW9bh0WzhQTU1bOwDi+dQ0E0gFSdz6vxhVpChmygKbOCpnJ9tj77fH5wdXbh8MByuiuLNhAMO
bDotaI4TH9s/M3u8ehLi9Us77rxRLxaFMZP64JS2AJ2Q8CGmyMNU3fu8g8T8unl6J6YgLr1mpQrx
K8N9mQJjBBn8dRKJ4OqQqQwOvg5BvJjze3rj40KDryMlQh07jPZZRViA1o1QX9Bvxt73iqOoWU3b
O880NR1/V9z1c0L9RVxvxv9hLeZb1cP4Ny2PjjBswqGR9B9y9b0CIwGfVh1tbJf3X1Omq6IBr274
xuj1uUE4q1Lbu2umDc89yFs11zSqoBwgR3TNHtN0mvi1PtCZRrO0N/ZEhBgSRLS13tD/FQQBjW9M
2r4HRRaBOJ/fnMAHBECtpTrBxSVetfpL7CWvKU2T9urIdoAPJkeP3jDZfLm/6ZIOdVG8Z2/eB6qY
HQsP5V00JQzgUadye2AxCxXfiE8IzNiW5MuDS2srfEOw1bYteuHSjqiJZogQs2sMXFWOJZRuxy8W
H3jQxvsmSby1ch8BARv0F0COvkLNm6FtGfruxw1G69Ut5b43njYFtdYTo9J42VXJOpYqBKzmpo9E
CaTvMNaxIptCsr8qmkZKsBtcLyuCc6VMPWKpcJpiQsrrrmDgJKvrEh1cBfhT8urNpTYTExS3Funh
VLZNi2pw+Nz3ppJ/FGliE0NaGEqXt2WEWykOJL1WZ8Ehp9SSB65CdvxGSZq6gkVXrLICY4JUWFK9
+dQUx4m7FQ5ORrqAQRmajkdKjMMqBXaeN9dC4UEAkEKuwstNElNUK0bdedYVHkNkNZLsJJS/1S8r
+P38WhfAwhO07JUwJ2GJ0JeEFSqtcDZ+7x0da1zWSlNi4hGg7WExNzaWNAw7IJ4EJ0oly0NyfsMr
35SvNynK6I2K94XbP0BPuyTp1a806zXHCrU9YFPLddgEJ28BoO3CPMr/vWL/7apY6PTZLwy8gOV/
7QMYplol+4kIYp+zG7d6Vbi/9tJzMUXQ9QuJcCzBfHUJMz3LVaEV5JhJCoHo7fK4arr7kzHDTAvf
8GD02JeGp2xkqP6oHJCtC40kUHa9Bh1i7d9W3cO3Te6w8nnUTKQi90frWh9ZG7MEdGxiyLZgdfzO
FBK3Q7O4SxvyMUTXGLS7VzUQmYUDD5KcD0hu1EtuSbVLnHZ3jxI3EONdt0Gsq3uMFw+WsN8Qdrku
k81+AoK4BkRQk1jkZ3s3sYSJDLW3nbGfsB2+bacUnu7MumkpuD8CZ+luJc63uiAiOJXHhIogFSnc
jPf9svhNwVGQt3seOSL2v3jDav51d+H83VTY+lix2XqkI6RxKmW0SjBXGknSFwHbDBO/65jxp927
EgGL4IYrZG2gNyKqSj8z5/O3fM+I4Igq528Idjut6turl8D+jEX5oKxIyRqfVDP6As3zaMVOhd2r
eY+zTBI9rYSkWxoTHKXBXxYKgPe/AtbXYKJpA17i1Vgcg8kxPVjNDhlW/7gZLhno4Qxto3m8Cp1i
JsFbad7HWu6o9Bl++SFWNfE2KjitV/mA4JhBzJBYdee6WT9EHK76OHWSOI09vEdRzYO4UtzKmHzE
dqafbEey+Wj3vFnuw/UAtdhs+t32xz/6OsCV9m6JBEUZVgLNYq6qiyv7Uy9pYr7VF+Ibx3JnhoE2
nYDljfFvQMZDXaH+7jZmMmCGRdMWwO2mD9+F7uNvaLIB+H5T2rWwR3fX77hMAya8+IwLoNl+JbqS
lm05KUJ0IOsY5pjqvPNXjofClxXf2/WuhrVtUYPVjrdLd70TLjXkAAUWQZgjUWPRKcjsGHMshLkD
2RvlltTtVaLmSIGIEyc71RQGy1kQLrwTkemDP7aDGcu/Mc906XeOmUmmG0gQU9rl2SSv8rgaN/5v
5yYnSxCrF+hgx5Dl0sef8lVfyzNdLXAt5/Wi+2hWgVPR0fVDYI6nhvhQeZHEFOSFeWLoZ/Msv7/k
W5A+A4ZyCvCUhpkJIxlcRLYcXJAsUMtk1AGyKZHYwGBnxqwF5dgMXvp5pGXfw7NUi9HGXIPliyp7
PTtyaoP8kIQY5wszNXAM+NFR92gnIpAMH9y5/3NjO/+Ky3Gv69SeTtrNmULk9hBFiFmRbgBVPWSL
aLZ2CCH2QJH4ObHaS/EHzC8v7RXKK0DM4y/cAJZstX4F70SD/TLr2YLdCyf+QgaTsn8J5LeP6N9/
AqC/QGlW8WGNU2nY2XKfuX2ytJGz/VZmvOCkhqkMrQu4z5qWb7RCqWEbWpxt9oz3T4mmPoKpBPI0
PnW4/1RmB+6bI37prd8ku4Dzw1Rk7AhhIT53n6ZUYHIFCvfud42YhihwvBkAQE2L3nLRVQmPvsMf
cvZXzW7NjqmEg65COc2FEQOxrwpIFOc0Y+913eGfiWzaH77axNwCETJjOB09SlrKnE6CNBcHkzfo
TSCc6GTv0NYozdUNo0a3tSczPhywycPq7oEOKt8TS1qTI3HMhGLDgdphK4Txf240aVA4r6kWgUxP
oc5kEkYoBd5x0CE+eyfim7GIBnHFpoq7/2v1dTYSV45VCE7WVlGT1VcSJv+SOBapQz9pDkJCi6Uo
kJzI21Lg7Yf6R+hqxYayGV5NKOxR6tMnTywBEN3ZbuU1hCE8l7PyRkF26aaz7KmVlolhkX9Aswl1
+XDOxeIQpWLQc3yL1O1OghGnbEU4FPI/Y+GNd5H0wRxIiOgD2ISvOoA+7dhtplSCg3MGrl2lGgz1
3uZm54Sg+/+meYLTD/jpY0x3slwh9ivdfidWoj4nOLPFoBCiRDb9xzIreQOXT83r95W/FMOPRlWG
S+8HJmLmBDo2e3ejUbSVs7mOw1FbGpBZpas4bz6ntJthCJwl49PW/rqTECkmUqKFjDnUHLQV7qjV
nK4Uf7tmnIzXiYz/g1rIdmtsg2FUB5g29J+GkdMazZA9KVIrUoc/8GXTT87AFRM31tMdUGrkTelD
2UG1+RnhzyQZbJQKp8E1L8fnxuZy4mc8iGVnBtWmgbnh45FkCm3juIddu9pmN2j2mgV44qmfpZ9F
Jm4CxxIPu3j1SVKMFXbNtFcuFDPNJNYByMS+qn8W8ZWMlhY+7FQ1LAZUU5chsPtoWJ/558UjAhGj
gfW/X4s3pSS7QAcneokIdo079GyFFsmUHOgMq5K35SIGAhCvpIbd7mq0hRWdYfJopkhiWU8VsBBv
eFSoZ3Dzx5rvWXkr9AryxPpjiRBEEEqeBzjWlgizn4x8RYL8dxm3weWqGyU44qahG/MewIRaqC7o
v/7HiPipfZx50Ms08Pjze8654O/SqCH0P/s44BcUgAJK7DUDost0U1FguGPx3A149XdBQfe1dsnv
TEvQpiJBIeEJAzVRUcBIWvZRTmH7UU4+qrv8itOKAtlabq7vUppwATsQbux+yFgb2hMRvr33wpOP
ZGY9zGZOhDeuBfQMz/2rW8nvIUP9TfrrnAS7kL0/prryiACioyBeBQtebBOZrWrxaAWbLNKcnUB8
y1rYjBTRb6eszlgJWHLV65CuQZO6p4y/hAM7iaGu62H48AhNcS540/7Yhxfy+F2ZvH4SAm8/56bt
8usGbvfSbUMp2dcZRyQFBoLpV4/B7XafYxS/iT0f33m0DJoD6Gu7AzJKdI7kuJTwP6j2HJ/+zZEh
tO5Hox2AbDdceGvYJiPa1cMHGjH07n6EwADWx8fEI3HKUhmYEKIPd1H5SV9O+5xrGWPInZPd4J/V
XLm+xtS5dJp1pNDxJCUEdQl4kwZJJYDFAttlUDBno4m4RcZIcFbWRYIt47HjDCT/5GvmHUXXn0Qu
xR84BDJp7J/maVzsGdAxCe0MhpsDYQSHFUwE77VuciFO3VerWVm3k81lGHxpYuDuVWa0xmx0OvDH
Xhrrifv2SGtwHHjOdOrMzCzhEtVWs2V74chYzLOiqOn+1hinLGEy7wxDFXTKayJxgDLv0S6QQJob
a0vXk8ZZ6U6hy0JvOsgqqvYqgQyA0jSKVra8kAnk7C/3qf9uIHduqdnIajhi1TKiLikFm8Z4bhaw
NiRRNNwc1dEMlNUDL54+J0+rvHH8hDjU4TlgYfB0VZLIzMsqug37mne4L3U5Yeb2cqgdLUutpZHE
qwWrq8eisZeaCYJ97E5Oa6pbb9ZZ2FmTgCCfAS6Xov7TSNCOA164peovU1/iJM39kpwc2JAZcO92
PFwasYYkd85gmwHfdi55WhBRDQepikU2kEXfEDKrdBVcLEPwBjNEwb9fvcVhxB72Z1pv4GWQH0iZ
dqd4mtJ7GehgT+4ZtSgmF52QqnMvTbVmYKSIGA9KFWXgAVZF/6SB06S6iV6NFaKLmBtS0hr7yS+q
dBnJRKYJxWOFPpiRCYVP4tuzNAadecx9QZwQq26cTuhE1AbrYCrOjdmcigQoA2Uso9THdFZ136GU
QTkW/DszgkfU3BGYBV7Aezs1ybViIVvUBUEJ6e1J5kdHxKuc4CKjycZAQUWQE27hTPHfQ4U0wBRz
6pBrejg03+QeNj+XUgXWAQOQipVv+pn17ldVWFAta3priNUe71c66v/eLA0kP+Ei9TobfZjiz97S
vhec2p2jUHQowoJpywUHI+PjuLdrdyPCG/xTlldghcOCg8loh1PHxGpfV/oN5PDj89JcOKa9gGCq
JmAm53o5267TRl7mSfnpqxTiCWpYgBOOviGk2QNdiQEjtSW//mNFjRfccYDooi6UTpwZoPak6LnH
4/1ljBLiXyUEEXS3+luKgOMcg3Svo471ZZ3SsZgp3GpKOCr1oq7hcvIoJ8PCz5/ifDevf6IYhIR7
b72sERulXno6OokGo52pZ8pqLeCTAhN5J2CTKfItlBC/7s8HefnxH7VplT2QstiIVcE44XmgPhPG
sBwr0eqQ+OZSH9tk6T5QmRQQKo8n4YEL/aiayAjsUTLVQ2R9tzGaxIMNxP1lSy1N2WRFIV07uTD4
0finPELvnjDlPiHPCPbqUSi0AzU/7KXkEevdRQSLrCxeOuT1YbxOK2pWXWI77+hYLUy/MBfZgQ53
2znKOWKE7DiGAgV97+rIxVZJ3K2NNVO0uAbxYpHoObiQOMLlcOkCmUFJihmFBSYkaU7bm2t3mb0P
viA1Fr2NGuO/BDH+e0LSqOnx0KnH5aqH0QJGPdV1Ex6vPtMNwWw0KrY9VC9GpcvKKpVWUX2PT35Y
7a6jFJEqkB0vTysC4Nf/0nExLGG8ygFhCnWxLVGoDL3vDDuU1u9zhKJM2eIH4oDdDB6m3qJ2XjVM
VkPHp18HIhAfvMoq24GaWcvrN/1EF/DSOwV/sfKoOAvgFgkCCOLnrBAOYQfJweaW47kS3Djh1DRU
L++hni0BcKuJMErIU3iLgJVpFZnSf7McsWNGObagMBp8ID2V0GITw4YtVsY04RlyvEQn0TnzGlw3
KNi8yI8AD2wRY+aZ0VFXj3uDFwkXLRAuig+iJKdXcrCwOiaaFZmRQJT8DG8iPOPiipOgN84xrPxp
fwYr1myAST9Rv03d/CsUgCNkiGELF9DG5JPuly6pGhXXptoeHktQlS6LXXj0A4jRfB2qTg8i7NIG
UyyKpPEcVsdkq4R6sTD5DgYaCkbq94MwV9HFuGVotkuXX4aeDMDXGjERLPsuA78VzL4f53mhV4Ub
ov5K1JT1GqKHIK+GQ+CBk8IHLErY/sOhtkocXNbM2xBBbIEQuSl/nESHCeBdm5VcQ+BUTC3dq02p
H5INHrQO4gmY+R7RO8VX924BuQngjeRiSMGHLBlhC7zZckSysyXqi6gBJNMcTidKS78/eL1o7O/l
XB7LMFSppmtV3n9tyQc0Q5muRLx2GA7kvbrUhgzAvYuClqydQm9LKCmiA/80dZv280fl4y0wkmMK
jiktXtJOl75/aUTt/5a/nY2NXmIIb+GPn3J4qBRIN1+1VMV7UIbD7R+TC7rw9Ki5zxqjkW5gTdv/
2QdyFZ0Qzhv9QFIpmYLSiUoq5QRDah0IBLuz2c558vkNQkNztZQKmiB6TNx5nJqI07pfP+zY1GZm
nXTEBIz9qUEH0uh06ZnjOUb3mR85zhU74WADK1UI35qBPRedSMkPwkqIfoai8nQk4+YL5n09i3HS
lrYgETZu3YDVj3kdqxMUi/bQsMzbrrQ2nGI0jlkg3X0p0QDhyNDzo4+r0lPqu8yDhTIb69QpOQ0a
fir24M/qmkGG36o1y8317tIe289Obgk8jaDrYYER9HBCRA7lgm7ViPfC9Z5etPNY2Z3HIvVPfe7v
tHilOxQocP9p7BDenMeXfpyY9RhlE9hFvkKNkXSshCqfzXdASyVRdGvyx5m0s5rWhyjjik6R9pt2
aYF1x0eoG9k3+/XWmh3BPzC4LPsu9VPdZZACT7rCB+MK1RSg2oK2eVRYpK5fa9Nlft08Uyoj+vsw
1DoMYI3vQkGVfX8M6OW8C2obheqhPawcwE4B+HBgeNk4ed7NtkBjnmFjOHchKVtSA3rdx/MUm0f6
cfYkmIdDoBLQrumXBGOZQ0s2MRSUIMUiPH8dHFLT7m3YquCdI5+GiLeYoa6VhMciWA0w9vC3KRLU
mQkbsg8TqBs6spspJK9wygnsdKie9BH4TBCJzjGlFDmdFdMJzjt42hmzuW1XuvFmrH/WpaWmxXb1
ia6N2EKE1jjBYRM7CTbSul54bM3lLH+Fhp0poEFNkvNlYBDTZYf5EImvqV7goM+0nGJ9rw0chXWT
RRWUClRiUzKx08Ai5IR1mxPbibshUCmpzcyIHdpEMEv2gmiI2G5KpHpjmdH83gk7osvmEmA6FgmJ
6SdxpVNrwS0kBPg2SLK1LHIFI28k7AyAvUojHlGchAuLLj4XWylytYp8qoUhk/MtiyHB53QWf/kB
+sVePJwf14nC6vz7WNaL0DEkWM11SeipTui/0NVsuBreRiNTu9GSR4dvIA1c2tI8TevPwr3u0O3J
pTaJ83JmiIBV6XTLYD1TDK7PsNx2qBrVpacf02wjSDleNzPzBd1i127xEXG+6p0eNtl9QfiM48JN
Vi25oZx+63GMeZhzOQtDWPu/A7l7VA4VJeauPKxNXoncrYUYngQD6ZP/X+Xkf20sx5yPkPxvslyC
GF1ERqaPHWuBeYEBbYOuVFan2rOsuZ7hR5JTClD0j/2zhJ7N4SPEJMPfyrvY9GQH+YaieFq6dNka
6TI7DtgNAModBgTWDSHuv+WGOST8VwKPikSuLFOmK+XfzRgTbA3IpJ5oPr5GWf64U0ZwYPcSLHws
0dMcSaGaefZ6zYJqKgH+N2AVxku+/2QC+xy8PnAhJow0XgJjMChszGMw78BCEYANiIdjfYIyzwzD
ms6OtmGCsYSfmI+PlC5xUEOlTznnZJL2MZ4VhqKpnZqtMk3arsOmaZbrhb6nCMLSv9FQ97//evkQ
r7wDMRK0HrFHKErJVHAyKAJWKV04MhODJyRzo2ccxuYzcR4/i3oiUX14NYoCVMLZItN9/RbXaR79
SoVwYB7fEyEazGiebtoGg8CjaAndFQAZubrwbd7S62p+VHsAl0B6JEDomm+mkq1gKl1f6QpK32rx
Sv6kKHa6T2dJQoM4oFH+Hg/2mETXy2CIU/TVfGUSXqzaX6fm6nLJ10bdlIPHSaiej1wtVAhasHVT
b28QKrCgJUt0hJB2nOlz9zXtbNdnubrjMDEe1PE3/0kMqmeybsTVgdBlhIvBd0cElbvEd9MrECCX
j0vu+dRLy6YuzSTITa8iOTgZHU0C/jZ61lqokMMClKnqWlpgniFeuYh2VB71CwsdWRF5bIxajsaU
ymy75oUqaHmWQaMSj/2Is0QyCEKlzKNGeISO/5rkx3ON79diCTfD2Oi9SqcElisGEL9WXCEuHJkY
epSnMAOIYJtitgR37P3TAcuOaNks02QPVyGr09V/FZOFKI4kVWWbmmN3kIYeHaRkuaD5aAdeXjBy
z+TZTwpwlbWDR0rsm0pb2CI0yK5d8Upa3K8y0tpxC6WXIX0a8AJdbqYsLt9Y23bhInDRPH3yGbuX
4OSIg8bcvsdyGkMnUunf9XGsWTezEDlXro7QetrEHsgTWQjpufg3i/lI2RMtAp+yac1DhlSJCfpl
m7S4R4Kex0hfCWLrvASVrlwG2QyWur0EBejvxjFqzEjd1/9lEV1CZMs9aJGwUwK2UwDClKQA75vE
JM01HxWPl3wb6JQR79/9B3meHvkKyxpuycZfmt6XrZZYXVv/nNmbDf0xZCgm+UnREvGZRgmZwQL4
9OCoWCplBvSeeCqRc9LQll4xEjNkh7A/MchPeQYtzjQW1hKv8YQF/hLO5phYLW/Uh3VDe1wA2o5f
olUXCEiGPu1yAZSGsy7pWthzNdqsqC7bmR4ExIRfujcmtm8a3Wc5E3DA/PRbr5qp26YflvI40UvT
zwV6t2B7kyyhRp9+rRJrzCbhMuKpJeeXKa8aSvwFzljUJ97DV2r9/P93TO4zFN6cSv5OeSmZ/Tej
ALE+JTjungejwoYkZCNP+4xWxLQSmQjcdYAGXbg00AsFMGD7xoIu9+tF8Gmsk92ooyAEspqr/MeF
1CBCUV4080rBtfcLwNYPUjTX7hYOPUoxsV0h2wxPRSQbA46kzTu7ttyAxbo5/GDLrL9Lu6B9TFt9
UJeBthVnfWWiqODG440k/b7nWkt7TWQHQR8t5qJD3mYzh6dR9nSMVZjI4aWkRclg6va1tfz34ceF
PvKy4V5T4V5bMFRCpJzpy6seXOdcS0i/SKN8/zA1T3CyH+TjmAJd5YaGMBFd0xlzfOWhAfawyjzS
W3Zwp+VeQuXtS21ZJ2LM76PbbtcL0z+Wx9bKfdtf2Gjutaihbcf1tw1jQN9DXiekLWZI2n5gamg3
YO1JN9mQqr7hOC5vuxynLG9v/aCH2aIMhuBYOx5sUTtEeBZVgVyHMQH2sLXbrfhNjfol+uQ+Y/JJ
zBXTNXoEpXGMhlvY1yUyBBnu6VaFZo9klGjZL5C6r+psiAi+rrWkDqaCg3X9s1TbVmMh3bgWJCLZ
SSAqqOV2YTfgkYUH2K8m2lR30WkahKzeu6jQ5TGvq0eG1u3EdGx65KNzFRBcgFEtCVXWyMqNQSWH
59onMMS34ecduZtpM0e8ARm1S+tH6ChGSObHMoEU/bbP8hvWyrXlv1BxEfqSVv5dLeh4tRgPBMX1
mqXSL4K7sxJZChNIvpmGaPclo3saPfYaXs993VdZd2OFpBSF7P7MNvNsQ1n1WITmvNn3S+B7gFTf
sQPlon7DwLxnrWgUmQ1+LyuTDUf3Y1PG0tHKNXDDoCCkQxvEttqVAWLvUl5axE23rJHSPMgCTzws
+bhC3LCzcCHufhWC24CbvyewoSx6W5b0B8doJ1zp/OSINOlCZuF5NiLYu+EaGeDcz3QEoqu1HpIN
SWqW+x9iK8mcbU86ixxOmOZLKS+3HnDh96vn1IUgPGk2dJqAZ7hnTRLgGSW3XWH9752cZTjmNqxl
s/NhC4vZNRDYko+GNSSypqdwymHJaUdXzXpooktAnKjpLgdMB3rtfitOZPPJ65WSg30YFF74KAuL
oyTO9Qu2lhPE7W8YHaG3+bmT0v+UZekTh9JaX90lr5kDru2V0+Hx91LQz3pf1YjyuaxF7Gb2OJGS
xsRvklOZfUULa70KSO7QikkAQjkqxxAxw/2auQBxr+n2WLRSjW5vrE8BsgVjs0IpAEe+G6V4/Pmh
2PwTkm5xX5Yt9ph5ab2Z5WX92P8+H3BrSBXhCcyqxQb10nc5ir1WUAlkoXfgERZeb/gyz0vzZMzr
iuEAzOGA08RXI4h1aWQBtIi/DbV60U4iHsZbIJ5kqsFeTG8bCE9swce1h2wGlgWAO67Bops8leAn
IGEnPojqFz1lN+YI/8V48Fr2vEyrMemIe9WJYDbeTbNJP/zEkNRF8YLMfjLIXjJ1DvYOL3LlUVI5
sGEqg68kr4PNWoQjqLv9/4d9oW168LicyVIgNXWz/2hFmJf6PYIfTme5BHGfd37CVeqQgdEbTM+D
KDGzD/ji7ACA5OvdfMR9V3ixHRMNFTJB6Zs7294f57BjpcEHAFsCkKyAsek8akLew8hkkxf5vR3F
e9iVQmpJ0JrVTk+JQVM8MNsmh02X0LhBKb//SJTAiN1QLwZAcx8bMsZUKOGy2IA9BjjpQrByB7kY
w6Ljnot89FRa5ZednR9Auk8TPW6Z0ezge8udrqoQsIBqI9XoN2U449q6FgFpFmjcY2YhjuNoa8A9
awV9Ru6U3mGsHspzTOzsJVdgJqW+3DTjwE19ojwSwsDcNb9gMk+jCRJFVSWIsVRiBvXT0QLOaAi7
/cri0oevW3jkda4WAvaKnxufrIbxHn++/F4uT3zzyHnQEGJjK30/iGyEbFh9hbvDhvHCsFOj4idS
5J3+UID4Ifa36FX45WGRXq2QiT6oAVb4AJsoxAGHGT3Kog9gLtE/8ZE/XnhcRfBPcqaOXCVvJFU0
FfEYb1kUTgmXorhytwCC2cx6HzQ0FGQTodvqFEhTZ4j7u9EdwFkZCa/SebG4G3kL3BX/Erf1PtFm
x538beTIw8qRh7ZTwOa4KdmAWgJbEiCHZW2fZBxgkckoXb+opLvnqJekrP0k6wh5VyEqaYcXtGKj
H2+ULLPm3JEPJwHv5VCF30k2buIvCoQrv6k+AihTmA2RulwCcGxBM9Rt+hEDbefjh5Ll6ONOwaAA
y2CKU9anvn1dFz87rc96USomyM6dwfJOG3BX+ULVdpuy0PDvcqzjuNZNpS+hFJ6jMy+qdujanCGq
luPKj3vtx+er6vQqz1GUoRyGrnzNjUfxx0TUvTJaEu8O1O/vOd7+7qWuSpKoe2aXrtJG9APlWKBG
4GyscqXfwLMzC1rM25k+HFNqU2xen3NPfH1mdpyjmB0ejI5VLUpf7Cf1kSAk9Zjf4YpGqEqKfE2x
g1C+4wrvCjf02dbJ3f9oAgslo2cKY9732niq+EgnHrN5Cdxc+by2btiK5wfQEWMxP2mD2L3UccRf
vx9Hh5ABOg87PalndOnvmko1wtwnYEK0urib3RDohNubOYIp+17XPLJkNPZcOSyK8y5ZJJwmE8rV
RNagD+rlTA2LsSAMLSwLIQzk+kIc3SjBnqDTmqylYBm8t4sRtUQDUAng+b9bztuu2uoHgCIdIxdr
cuj7ZlsLE1lQaU0KNQrc+Pwz+DBo+ZSDxIZdxv8Q4rg7xQTt4mxVkBbYwAkbvX/SDO+pVAoWmHp1
Bd+Mqu10whjulr4+lBC5XbWYe0nIlkeGRkoqeR0mcZUwD05pYOfnGFnuk4yE+VJhLXuQNCU+7IWX
nMXDqSQyswqHPIKB/T3Q7L+Ey3BeIAe0PcvnEMe0QP1efroGIb1W0BgRT+W+3/NS9rthRrFjK+Rs
vmJiP3Y4Gnsj758CFPpRYb+6ilgWty+VQVlIhhNtvjbTUJJ1Mkr7zxbW+1HHJniupteA2o9lETHD
7CG1k4Fx/B8k2ebUiBSFFTEMRz3NPPv0c/gldgamyJmGW4r4mbDh9wgUC0dQTjovEMSxO/yvtnIX
dk/OivkNmXd/PA3EBaGv53UiAv7Obz8WQw/3bOtZwtRjTxNXw8Nnv5Z/AetDySY0fcd6j8J1W/os
5EPwsfKLSQxizJQjbf56i+tADRryV/V1QDQik0WagHH+lm8R9PXYD8wudOQPPV3ro4oHGgpsZrgT
8nB9ooz+dBHwPKvOMUDRIrKFLB0fMirb+ZY+sJXkKFTUZUJVF5UExbhvj6iGalZLtwlh3+oz65Rz
5ELXXxzYlo/EFApFGxbGgnc2aQrkWZ6O/YebO0scvqcrJ5t9G4cvE4WbpoVjEiIpIsWqjsMEZBeM
u2EjgH99S4A9yyee3Eon0cnnTx/TBkHKHPCY11hhs7cls4FXSnc0Vu8ed7QksgU+hqTCfqq3HILV
lFQxi8NH/xawa5znIR3AgjJV4F1LqGC0Xtb9RXZGhXmbvoKXLuLDp/5MjlTif8fUO6aCY8SQ/K64
U0vNPHJi9Z2Iw4W73gHDEmhw/kfVxly/oJm1+xE81OGFZHTZOEPKXeYaKM9EDhczPYeRNxvJF/dy
eGaFfW4NgDDC7fOTSIgUieOVacFu3MST9vI7dNCORYDsEEGKLfBJFum1OT2K8I/U8Y7owXrNRxsH
9jDSZDJmbI4KF3H+Tdn+Ra+GWFww18fZVF7WEj9n17dPEID8Li5BlmFvr+R4G5PDojdRpxwyKB3+
KBUOjfTvcqm9DIEhmiVlJVapRXsgTV+n/gj9Q2nz8sP8xlJr75CnUXggW2jhvUrX4A+Pxb4bX2/K
5vemJ8QPkRd8Y9rjgbKTQ+lL4M9coFT1W5iXWt78QdjyB0k9tdEZv0pQeoWef/Xfop2Oz967iswU
0+dSJGB0hL6JyH/DlNxVFKrLMQ2qzM7L33H+wRLqs7GTjtM8cbwWFKuoEp4AuGhiqqTTJtr1iw3v
kxISXAl9SHTAcl4KHtAXIz9a16NrPF1JSOMr4Wamm+O7hoLbzWdzscK4Plyh0W54wPc1JJb5Ff6p
hdyZrrpdLUChzzs7U7guIK9ScHTNqp5cTSNvmSH9uB4EnnSKCQ7WSAkCsxRT+2v84gm5vgYvLbx7
TemFaoiibnhxzTc8trdgS2z4DGar/OTa1OGNh9Upp5NK6d3X3e5wn3W9rZ65invmbDNrU931Ltzd
I6CjCie930prjoUfITkUBnV9biameAR8qlu7jyVpeX4+4gcu/8GtOC989KJR9+1vM/lvdPrVs0mO
4aa+bA+V2MPdfu0RkD4M74wEOoSDRK+rqS8N5bSyIsRwxzy3TzjKeKydKXPimJHCGisH32zcS72/
QnqgfqaadXvaGbCbb1HUJ1vqLb0iafhW+9eZimsCszJrX8InrNBcZ/zgaUdCrhE9gQAJipxXVynr
Ns1fBUybaiBuKQlfFujzh/Ig2lJH3OUWTRholN9TQ/jfnReh9KETSZn2osHZdkzgE3NcwNa58KXm
G1iKn72IOi2i9X0FghADYJiM51+5mN5i9018DXlAjTOcEyQmPD+UXnQX9MKb/Z3WHarsgCluyLLu
Xq7H70X8NAv/MGOiNUz7jcc9bSYRxeR1ZCRQuanY9R7MdRy2fuQIBya2cnjQLMmNz4R60zMgJK8A
3e3B9glGXGoNMIcWxh+UajnOFkB9xRV3xazARr5AMuNoFqxh1LOfTZedf9S7/OEYAkwLVrbKAWp+
+8NCzG5tDUG8428S8gN2nd8Q1DZ2GcDTyHsY0ouU0cT5BTeOS1qNMnPeA0F0/yimQAxPE2T3yNlI
EAXfUJEQ5Xb104x4jNKioYRy+FaUglgMpF3kMrdAGR/7c5YJLpHH1FJ+oF8eJsYu+Msmg+R1UMTJ
8YUUfv48OxGBX+45lbcH5Mp64SZ/xbYi8IPYH6Ocvj1YEgpL3464rd6LYt7aKizl2nqMShgxaERH
oluqold0EJx1zE3PvWGaKCawriB6rGL0ACcwWRi8t7zQwKBZz7kqHra7lqxIGV9na2NLox0P/ikx
KspLxVDM9AV8RFRqO1OyC5Y22JCNN1DM606ZVHka5vhkBvzzHR6RePl6TTHJzQF0gAIRwdCM1yka
xzbo984XjhOxIu78YhcJdCMSUQ7uDfMZgvpeRRLE/VvsPuYLu5+okVfPP3P7FiHHl1cuP1SOJuKX
otdL43vNk0dNPQ3lcWAtOzLx+sFpnNJMPF5nseqNG4q48qwFzdt87u+GLwD/aUv10ERf7mt4rHi9
XFJYJVijQMt9EzQ2IA/bgGB64apbiOkDnUoWicSCwMS0Qf8q4GbuLxppEA1TTWKEh16VNWcVzmb9
OCIQ7Rh6YDPNUQoS9hLeCvtIk6A+SllHd9GEtJqTrcq9wlqlK7AQc+MWylLUzU9xjQZhxm7hA3iU
7pu4wkcQcIsHPL2BKy5fralC/P6mtfVo4/Wq6n+FhcOktuFpPQq0Om3WAWi1Gpa4zSQtAmKrgJuO
6YLOyUtCsaabWKbsuWp7aqCjgWiuO+KitHS6XfvFj28LpNPY5CMxS0Y8r751wQhAyNxMcjaAL6UX
bp14XEWCXpkwZsembWFA7NScbQmKQrXLz43249zU7uF927Zu2Ja66B80PuQEcKDWyWJ2NJYk6LHz
7tAv4GEbznMpodcZzAtt2Li+T7VUyQlC0vGDbDQh/c0Z5fhwGaZ0CGBN9A+6Vf0qXxP7dL09hruU
JjinlWj5kaOFPxDdG1faCpTUqdqahYBkKYuPx13UROx6WH0ZmYrJ4IWaCzDH+E1AxhxpYnN+vFSg
NweDUzUkCUuubxo32C7LcnqSnW66xruqvBPQZbYYNTSv4+WyLfPRhsDC2Dw+CElNq+N5pDz6dkmI
XJsHZGPYqlGgu0h6n8P58sjA7qU4A9u/I8aKNoXKxcd3pYFmRkeF084FMW77dUVxkqm3eUgaw/tT
8J1tcm988VUfXOO1U/ucrA44l+T3/TE/JhvqZ0vRe01sBENb4OvnVRsv35wsUdUd6fHU9aaZkJXi
Au4CxzHibHltO8uXq6Toi1aNhA6paOyqpXVyHKYTola3r7dCgJeiXRWyqTaD6S1d8YfSrANHvppM
C589HbR1o3xgUHXCtl7+VI2GLE5dml3k51Lb2HTKJlp0aalOWZ7BEY10wrCz7CKoLpj8vTUgtFVe
G7ERBQHfp+7o8SUFjqoWKMdf97supEMrW0+6f2xJW1djtAGbtEfVN6w27xW7Gk/o67gD0aKSW1ua
Z+MinhwCF0m6HbH4gNLGljThGqEcWW9KzyX+eMBzwFlQfYDsUwrl7PYe+DJDZ9kTUkAHpw7iYqZx
eay5PLwJ2QfCA00qQ1zQdV9QG61lEyRk6FWRKucM7Jz9l7N+RyOw1jQcOd2S9WRu0InMzHn4UnOo
J+2ADM8pAjYuPsIizSsJPTJ5UPfIo4ppzZ/RRzidQ0lH3zevyEvJdauyt/xC3fEXQCWHmVvTxS+0
vl3DnDHQcSmDt6qU8JuvAftYN1X1BEhT4CNhnVt9Uzfce1x/rKo96nTn5irNWMlvU/+87gZ1dTWf
AgoD6A==
`protect end_protected

