    parameter	EnablePLB = 1;
	parameter   PLBCapacity = 1024;     // in bits
                
