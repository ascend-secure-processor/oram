
	parameter					IVEntropyWidth =	64;