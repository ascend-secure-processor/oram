

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Q7hbl0RjbcwyKOfDj0Bh/cJ98heat/v/B6itvD2hDie3qw/7UKUwH8bHVmPvhUJFZGBrcoyG7KX4
k6IwWmCgAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MgsJCbHtEHfuaVY1CiyrOSdYIIK7rjq7OjYC3zCEllrgg9KSWHvHZNrKKwntDbmtceaj0l3vsA2x
omj8YSfqGqwkDVfUVIjLZfQW0DOQIJzJ2r5/U3O9vy9+l/bmMNZwe0Es7zzcEbu3M1rf1SGCbncb
WppuV2IsQG28xHpCZuA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YNWJAED4PZBIxsOb/SatK7nk54sYk1XP2cr+JLIZa5g7NzdhrG5gSvEPPVVw0PukD0xGyhU1csLX
pZht5dD+qCRbWWA4mJRLb+ur6T+YaBYDiZPWbLapIembFxEC0WOYryrjfb8xV3ELfgXp5I93hKdg
f3dIyRfLxYMUnVldHSzIcTM5bwnU44boF3lRqEsSSldWf87NT6/RTku1z7PdGbg5OoKywjgOxl0v
ZOF3mPLSSdXsd70b+JfZQWfe+sFV43Dy8TzdkkQ79nLOOirYX9z6IEyVZSVwuIfmaLxPouSvCn/I
pEqpWrYsghlXFygpKexT8J/ZGthVNW8QlgqR3A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RFRuJ4R7yNiEuDtT+8UKS2lgkpcE0RXuCl1d550+EWjh76QC64ioRSjvjvMvDWXvetLE6lqp8/I0
oR0BaoALTh7ZKHtPk9iFjOPMOJ7EjFyz6bH8l5+D8K3AowdlfprW+IuvY4zm12pgP8yLRdLg7FCv
nNdzvxJUuJbq+VjZya8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ci5XBgPzKUCYTv25+FhUtKoEfiRwOFKb4KCY+gYi6R2CmaBrBpJSautWvDNDWbAwCOUFXrx/H0Zj
nrJsceGmt4TGxbNZUpwimva89UR/qUTFIpm+tYVRo5i3Jc0378XWSL6i2sVzh75/BUU/4RAlCHtb
UzkCicCfWJlMjVc9mgouAVOVwrAt+8NeXpYy2Ti5VOCth7wF6xoERkXgLIneC7fhCHuJ1oJl/1Cg
hC4Wj5HmAuOsYWLpGtjb7DNyIZiqltbXkJ7AJGeNZJyp2LE4XfhrRf4Aa219Z3zh5EJ4XZrE6yEY
SJ6Wa2+NRzIRaMOX24Nv3pw7Fs1XqmhE8wwvPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6432)
`protect data_block
UNtxdcfkeuxkjuWRNE28Qf2UFhf5mWvEA8H189s4z8wTIyO8xg80A0X4s2UpbnkvFFrwFqFpD/h7
FBz0+6T/lvTI/Dze7xpLNxQjxEEHK5hYqTTwnZUvlzvE9IN+v51YEzn6IST5htnfrIqFVigArp6W
lNyF1mtECykd5KfPPzpX9V9ayobUV/KWnA5RGJjdNHzgMU20uQ0v51hIqZUjJRExCgIhO5HcU4wi
07ycr7OxMBonYGpwv98yJzCNm9WH4Y136C5F6kfDgXZ07BJMe5YZmNrWVBfi1OFphtoD1Me73KDk
hXYRLPW7/HhK1VqcacRT8wwBOXSnyMVn7bMDKS/dnNbWWEtDAVRt+njJWDVRZ4atY2zm6Jnsrsw8
jTY6zA3dn015Abj7zpiUPIBgEAKgfJz/U2dC+4/KeJgskjVPiSSmuWWOt+wEmk7gpdlb8RygjI3J
bWGamVxQUqz6ygE1Upa7Kndq5aJ9RPXo/G9GZfXR2a4XI3NU6DZgqBOEdgpVCX18HIvfyuvcr4gh
p2DOFogkRjGv/G70A0K0cgQuycVoxHGFNRewJGIf3YI4OdICc6U/GgAzo0rKCIcVlCo6KLnWViba
qWhIQsEWnA2WJf9fhbjxrqSUGdO8z5k8dkh0MTHt/yYqkKNeeeY/+ueyFTqiPqTbwwWR/ueD/GRW
t1PKpPMLH+A5eP3MRuUndY0sBpT7MOcQBmqLbQOvl/RGjt7Ip9lcVKuE36CGMoKNJUjBQVh+UB7V
tIEYK6uC/YsYCXSh/0yAPTSdYX7+mmiEvscwJeZAT5kQI5g92qobA+dOEHfWTx9OE3G1foepkqSA
Dgkk8r1AiMMrSrgElWndxa+Ypxjraq8UdUM+C/AMeaoiLuAkULOPBHUbMm4vcWDL+1jYStmODQDo
s+8ijIWX50HXhQL7pQYsiPgPA7ePgJi4OWmfpodmEFGGRSLN4PEtrjXVE5DflZzYdlZoUPGB634a
ocKlpqWDqBstqYjyWOwZLAWNm6SQEx/3jiTZqFqg5gj1AJPuPNscCMAuBRq5zjVPf+2UppE7NffS
LNc6rzJZcwT7tXEGR1C+g3bb7qL236QapzwvYen5E0TW6/SH0xhGhk3uzubLpbZKpdnzv6O8xH7A
awzsCm909Bv1WgM+2aGshOtHofUHySD86QUWGFpoOhfaECLTG3WaPXSYXXeKWO7AQfiNxihj2gii
D03x9A+3yqeLK5Ylx8zvEclglca4K+gjEQkAcZakEpKYAXtPpr3kIrb295dmunxODCQ0Q/5WW3/Q
Z2CHlhGpOk8xU4EZNefU6Kp3lk2fj8CgN9Bi+GiHg1qLZ9PBTmmOwlPNHqMq8tusKQ1s0tF1BVsL
f9mBIFkb+L3Ci65NmC902h2Cf5Q9QceK3fL5TLgRaWm3Gfdla76W8URkiHw99jAVxmZabsjZLrb4
f4oEaH2Dv4BAy8Zu8JTKAvTZwH6NbyvbUSvWR/q+EwsLjpe2sBcx4Smacgmd80Ow9Bh/8iKxRoch
Es+XnFNRhH+SChe8zse/XREuUJPh9lNL9o5AvZ0JsolAYkpEWjKXxv/6cr7YMuWZasUdRhShcWI0
y11g+UO6f5XO4nRnhVK3QdMZEdVKHsBpvrpp6klid4mXzPx5a0nKcswGZDnPDf+sA3MmBgNc2siV
ARJE52O6WrLq2ftgf8WS7Bd2gFGGKz+MNoWsIKOMnmqs7ruxZ2EyZD4/h8WsDuj3hxUieIcTuo27
KbY/3f0WYMRa35XSHRdIuJdg3KoAk3FAhQU4pN99hASRldutkNuhL/X5Tj3Ouy32Uck0oWJHJPAd
g2FnlMMmZR7P9klhcxY5Cbe2UL28ocF1KOiLKnca6V4Mn7/NzqpA/YDakb1R9ryZWBLggHKsibLy
B33ThNxvHwUwvJ3wAOEDbusHfk8lL+BrBorv9gyZyh0ICxCTds7DGiVWmswsgkGu33Ne3YdYfqUY
pVlD/M38L3gNbOONOmK4UQWiecSN4jubql30NEyXIED9nlCZeOKVHoxDWEleYWUSl/wUmk0+WG/P
aYMTp3raZKUVd0lq3sc7Dzrjwmh4lid6M2Oqd9JfXUXKS+1LmgQVQJwd3bLHXqMiouSLG6z+U1gI
QNFZSqJA/2KpqjeCxcAGPdVKpxIxuOgkqmpftoQN0Tb4dri+DXpmWArzKsOW7MopRmsWrxj88xpO
LScqHo7Ef5YcxQ57OHsUsIjc985ZoTppHG97VU9nmV7t0sSRaFLcvv95+t34dkHd5Xpo0CkbhEI4
qjkGULqie3zk6hPmckxDUTVq0TZC1+YRBl3eVIqzI6Ngoie2mCGKy4lEr7ReRMvT6d4NGDkT1c2E
AbFXjSy2g3etxisSf2ThMZyy3vdsxNKlfKzDzn5Nl+2/iZeDDc3m2+37O/oWhH7mu+bcxAQYtgM2
w2jl+vXWtEGseydz91xM2Y1PYQuKvg12Z6PVljvrPpo5ecndEGnXkcyr0/v4ycCYxTOGbz+WWv09
DoaXOSZ/OcLELdI34w8vDH9lBBdYyrSYd7fjYHGZH6w2MDEMUEf9gdepOikn3xhlrdrmB3riu8nN
r+bosd7mvjFTd9B6hNK2K0vvDAHBLhB7xGp5zxBl7qmeo97xjOI6SHC/ccN2ZrC3i6Di1OD3Tbit
tKrPwwnSxVVIlfsgFFPOv+kDmRnUQDMHawLPrcsGZciZqm109QgGpJe09BDUEmR+gMgofKfz0rw2
GAzWRVZtLWoRHmjM/5f+p4GDS2X+RmYkC5jUmi2uP8JxUqNoascevRwM7njFGCNxraFjntFAUSsI
pDnRenwMx4m4vbs94yiWSawCn9oyFxOGnKVGcHHGSuZTmvQnR3Qdn3CS8LkJRL8RnAtaboTpsmsN
O0Fuuu7mjxVi8rSEL5s3xqTDnKR7lf8ugXtxeJu3BnOFXiIMPdcucCP5iQmbF/sr0TYclPBvux91
50HICRb4tihoQs+gh4HA1SuwxB31btmvaiATGvHHVREhhKADPRvU3qg1qY7Fp50UI/9/XVBzvbGv
nNZzU2bopw4w664nZ4muqyl9AHa7UpCjy0QchS//+nkVhhG08mn63jwLfsse3mmqrTUGNi+8fGkA
7SQuc79BBsX3aOnIbowVxIkPuw2ZPdHoZB6ttvSdpzypUuSNzidl4cmbRZSpYRcS0QB/5FlZoIQ2
OP7S2xZC2KR16Q1BaDkCn91f6MI9LE5hH24Z9qFBONi8B0YhW6tsvIeoyh/vZNhHRxEl4pdTeYV/
sp3tdnpiUBjzfyLQL7TXF8vuhStIsl5YX8yk84w3yXfHVdlmUQJkd7MLE7w6aMEslLK0EatNeIFG
FzpHUpJMZLs1wOK2451oMANOksxuGbfP56fu+27pT0tGnySsSq13vgxfTarVDGLXT3XxXGn4Lth3
AmE0lmO0+HEUnvB5U7au24AKsRNg1GJvjMaVCjEDZP2X8s+XqDv7rEJ/eZuW+3h4LRiTezAljQu1
4diXHhAyXOPwGCA2wGmbRhGTlGkgwx1E/1TAIlwbK5rFFigedVcNOFfj/WQgphkO5AuVg2iMEfqz
yaQjjqCRexD9BPTY0N24KgtnWM6rH6RimIQ0QsjkFLoS2w5NhRSGqJ6zEwuAGkm4yA2eWdLrSKgE
97FrQmrwbQgi4Q89UP5JIN9vUv12N4khq6wnqZajXCCQwOGWCB61nMi4TSpBJ5xN745Eg73ne+uj
tGGPwnHvi+mfri6EBldX3pINVplRhxYLXFEpcZdcr8pICSRl2bMsEIxO+a6yrHDbgQYdyWBRqYXq
RrPaTrBf79kORMPCLrZL6As8a+KtUvW3rMNgXHwH3v8jNzB7INHRbtdCIavEHl64ah5WZ9HLm4yi
1ah87K0b195w5nkE2/pNl3e0O0usEp/t2x9IYZZbSS6xc3yRRPU3lxiqmAv8unUZh1oy9kVpZYNM
WrpKQzCXCSgj9BLC5rMOFMeuPse/5TriUQNg/bKwYX/NcKHteCVOyrVzJIdirFkFCDpRphS8Q+zf
h1Du+UHRMpGgRRjo5qxH4rhtt/gPssUIbmF9l0CCr/UjZ84gF0+GNBbxcyZ+2CeSvAN9TlNUXDRk
qPN0P+fJ2vGmkB/ueBhmY2hz7YflKS9cfQQbDqO0Rsrcc23h9wm8+nFn3+mDU/4dstf6+Aj0mL6W
zDNjc9KeKi0si/8z0LahNPENuNCwnu8xbGVJEgtDQbR8FujwZZIqDuf8zpkU85refr4afHN/JUzQ
c0EqUlj7OZxG+7nuSIbtnuEZrQaM3sw27l5mmfR1Tuqs9zfY7uu91JHVV157ZvWw2t8y3N48RNgj
SP8jQT1dIuwray1Qt86wJ1/tSBDOdX8ObQfOKP9xeIEWMOTccfMuqF/t3tkAn6MQ4mT80CflJzA0
xpsG/V4r56tHlSck4/GnKvaFgsXXvgKcaLJrpcn0QGGll4uaPpBpGmdzpR1UrcAQQRbKOBHSJkqj
y6oTWDYkr6IF/gHRk9v5Edq7Cb1ury14M6RvNMMwJn77wJgWgJyYvoMjxW1g576SMDJJ6QGAvJjQ
9Hg9abwxwlu6DXvlnt9eT4HfjBiuS7sghj2KpGbsLJ8lOhoD8xGF+2o0cEMTra/keRkU8AEuN4Ih
KxS/Zvd8OXDll7Q0/CfGUBqn9IWd09iqZZYGz5EKK+mIXSLrvW8Uoirm8D/Dodu1K/xkZ9NNa/eW
lIXrsqm8SHdPSrOJuezKxz5FzjoJsGICBMxkToH7M4BV6Jin48ER3vp4IRqdsf7rIGktIxTQqK77
NsvIDZXFJFD26rJVIMzhvZTLpkNTUulFh38pChXS5zK7Roa4IJp6YN7TMACjvJzKktO5+B4I7MUt
6hug4iHfBnM1eSUHx/OvL+/k8yIk/+Y6PFYs2YV3yzqTI+yR+gGP7oVIG6rg5dWtVwxutJfwfi/k
GsU+TllnIFQdDE/gSGxhZNXq6eM2tzFDr49iO6LIad0+hrxV1bSX1lVrYIec/FB9328r/UcbpZvB
/nblMLMolQ2huE8hlz9fwDQGe1OUb2Fk+aBMK95eD5nvSu9E2xQ8InAulQeP/oWVeqMyMDC47V5N
7MNJA4gRNSUAMl4xtXudiLadA0PCKc1wZG6hyQpjCOqRHm4q7HPwaYrzK8j9Pi0Df4YNYxTZ6q9x
5kJU1/ZU1as0UM4Y2uW5hKE9XVxTpbt9RvHPHG0euL8ogIVa4sRCm+l+gw0Wp3FwdC7aHA4xCDe1
ykyk4tG/1K6C8rjb4XAC8jm7ZvmBEpIcwtT3Vl94GP8eTLVW3opkAEvvkFvRNYH4wiFAZpCCyWIe
yQuiTTmpu4QdV6wUA3bmW5sa1BLq1iNyyxVZ7N172CqHR4iCl/2rjRVfJbtYgRbdJzHZoiB07X7W
j10kkh/cTtroz/AUBimmFP1h4RZwqrByZ0+/bC3DBUlR/PVUyjLxpG0PQastuutOBIwObxW+f/VE
GuU1YjNG5NtzpfpgU6OCJMWdfff43wQyub0Nxx7qt/8EX900ChGnnddDcajvXfFqVcC6TCT19RMe
BnnEkQwkvMfEsJGpaavQuOAx04iGZe1ahWlzg0/NmE1mJC8+G5IF7Xcl9MeKuXn92cQJvN8Oq345
phlIJDo3zUPYJkllPKwIZXDRB/CbNKzWC4kyybevumDVQuQAYZ3+iXzBHjGxucHU91ocNKpNPTW4
HM9nvbH/FrTd7yWq6Ye7RafKF5z1Ef7h3mUVXJRxduVdkzFznOvPWUQ5ECTwtSSUYEVylwIh3vwG
hluf6UqVWdBNG54a5yv1aedMrn9vNcUCHdXb5NbFnd+BgOh6ILDQDTS2+TgNiDi0wy3wlZLxLGwX
bbA+GKaTJVi+5UszmeqYClQNxci2tjhOWzsiO/JCgfOxBYH948qc6/OIU21aa2pynyYIhYnG4l+Z
vEB5+uUU/hSMUHfgl+BPFIDD6ty1ZqNajgB5Le9b3t5jdHMMicllcBPD0fXwyop8l5KpS1ti9vxP
Ki/LdV3nF0lEbQmCbRNGZPcm1nDiynTawmpr31kX30GZw8DZ073ic6BVntZKUiBoRXn7G+r/JuG/
8GUde2+x2Jg+EwdGGhfSCR+xT4HgC3vtZ3Z0OVK2QtADV3i3Audz0F9kAfgXn+klgIo7+R7zRv/6
zPYdiU3DW23i0HlsLEPfGngsFYmdi2jfGPwUq1Soi61jPda10u42OKY31H4ox+Cx37bFTXtlhNyx
wkmZouR6c74okQXHnpZ/OdK0K5WRD9m/EMbI+1gLVz8OGVFtgywnuy/N7sYmxETGPWSX80WjAt5v
zlUiebP3AEzXzn45UYhks9CoNW5WYbhUaClS5HXttRe0dWv38XdES9dUWOdMT/pH1Q330cfCtvMb
WM7RERqB/sUFSGa6fFyAFxxn0gJyUy9pPZbIEgoA303acrHzQuonquB7hLfnEXhQOOwVgHZ3dT7q
AUgvreRec5Ln4WIKaHs/8Hn9f1/QI4ZWHFLWRgHR4m2cMUN+GLuRZmqI0dJaVvHmgu8bo+FigKee
CeICgxZXeTqfAIFd/lDZjmHc8Lj4/8YWYqVOioqq6SFCcGLexnvK4fE3B+F/+YBFXBAmaBKtupDQ
+38XT2L2vTM3Pwa0f1o4SMsTiuXn+MKFWubs8R0p/WXjJXfesSQqbT0R8kdwlqlJIBaNxmpF0cMo
pGn5nw3G0wFrH3jsU63hAQRi5a1wovuml2folw70xHNLRckgUqMsnFqpgqzImpkkw3hkV9lXjGuu
1KFItWy0J0J42mtRPLWpthSmi3DuQSjqVnYAyAKZIcEdKRUINpb+2XA4Fzxp0eWqR9jyHpuwx/Sf
M69C3vYoOmeQD96bycUIJp7taz2s3esJgAk7dSj6gVn+aeyqJqhid5YIkULd1e2J4USGL0UMW5jV
M342gkN4zAJBmvmBjWV37LHhfn8ifm7eRhYr8SzZkJzSOA75kV4Gka0mqmwtRabcny8KKg2i0jJ4
W5k0yjo5jCuTKaf6Qj9IxyVNAso3ijw8argZ6XJ0hPcJuOWJ1qkmK2/lCiqpFosiz5qKH/uS3BpA
20b5+7jr67suHTX/gc+bzG21hUZNiVsuQGM8tCe5fe0jA3q7d3dIdszFqvf0rlEW1m633/nV+ya2
SyKGkx4WNFLqCqGCMyKPEiWC3e6MremaJnep+Nr5e0lzaamyDKxMAYesQYi5u/O1tbrMv7BMWcvU
n2qbSqCPJCne8QhIqaN8lkL/830xNXpxZDq997WfgOZt9gHstUtpFFvDGHkgpJnmHZZSfyP9HlBi
3Y3NAGzpCmeOXQ2wKzEmb2xbuqTyyTd46g5WHnv68s0qZQ0JwHm2k0a7so83h2zOqeGpY6aV15VR
ybPUPpeCXw/dtI+MesT2/OyhLfSSxUb7tT3lLzT0A+LxzWHAMNRVHHzproskCBT778ElPnT3n3Wl
qHhb6yP/AMauh3NSbxszhV0MbiDsGYxWr0R2wl4F05CkQlYaIQU6SgwOsvGaaOfiVenv9w4TnY60
LAqMo+1MGF4CvjNdhzRbz7R3skp9gDz9cmD1zAGqea6OGsu93vxiEqZzGiC6r7L13/4mntUUCJmH
+SZt7HK8KaMSt23GCqTA9inOM4IdThWKdzt/eUeSS2j1zx/zAxYWbfNw354Ju5sfk3zpo96ZLMv6
c8vyCbaYmzS4dBqqqJdiB7gJYkFDkZ/3mKPem89jPaPvKimM+Df6YGSx2TzNElHclCKjvT3lO1Sk
sjHlSW34KMAWW8NA7OtwZQLAVTOlrWKaHr3rKZ5JEBvfRcsWaihxYLO58a7RwRueZ5SH1QhnTCPd
iDgBcwXuyUxFVtXKDof5E2CsA4rQP479ZNPm0WF2+2eW+AUBDcDwbqYfG5wHEoBfi81Jv89pobsn
JqYZDMoSSLylmMNR1Hui5Un7Pa3HKTRqQc/9OYp8NanzqvU3lBhBX77GIKXG0B96541twwEdYqkf
mGWAisKs2fQ12rGCk3LVGlPqv0XZB7wfMN7CH2SrVRTGB2Qw0IF7zbCLnBjb2TduJV1wAYZtKmcM
O58TmhgEQa0ExrBVklAfWLFk82nPRy1jVqHdBmdi8Zjnfzoi3ip9EQNKBAUTCLDz9kqwV5D9lvqG
SvyugEgDtZOW2HP1300yW5we/L/4McwDbtkyd5x+s42uwImhx1+VYAHEjmR1459lIz2jY6zB1hzi
iBu32jLcHVBOy7VtFP4i89CMVz3ZjusU8aD1RHW7qy4DbkyuG2xVY1hFO5oG0gPln2TdZ8/ocsFA
r+l5BCV2+33i1CQsoVuLUk44qR+BbqssyWtZIhasZWrVs+dSMstxVt1f/IL8tJZVhspMohvQW9W/
+qznkzZfx6eCFIZB68PHzm01ND370oP5UCl2oNyLYprUnz/UuS/ErLgKw7w7f+TWU2TJ/H+rwtE9
IDE9cLFDCDkSB2YMy8o4+wRvu+oxpnSBXvCoc0mD0THh1iq9Z2AkLIgZvDgCWw5aIrsfJUIOA2nv
jf2MMynyms87YREs/EoVuTXtou6TmAyTgueAi3qNjbP0fj0tngGMRJ2U7ZLhEOO/
`protect end_protected

