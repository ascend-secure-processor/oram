

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F6k3P9aUcR+POD1v0vugqSgOHOxcTtH3i/73hzjm3G/Y7WtFeMPGlBw9mRYqkFMs7Byf5SinYMXs
f+qxOktcJw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gAXNQlJR8pfCN5KdBW++vcbpZhfcpgqUr0wiZZCUh6xICdJqGKC+nmcv3VhfGoI3NeMjttcKfKBc
5fUY9i29HuOA9z877uNFhF25esc2XKNsicJn1alndds2J7CXz7n0RyVz9/PYU+B6XwsHGjq4M7n/
8hXshGNN3NwZDtURyc4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
slk/0eyRMmi3RJM3I0xwfAYw3vuOWOx8pMhqatWvD5n+4nTkNmDs0ucxSi18aMep/r88gqh9DmmF
MSbKb9Joi4NZzW9MSviq4nB+r/cqOr/G+6kYphaXUhE40cXwhTQZKd7ljLhD/3pJd8ADjABy1+Yb
IdYzmA1OOhbl+X0dmHU+c+ENp7vUk2ssu4OEgiDHglsCB4E1C+mGX1bwFvEZ8T5PzfJnTIloA32Y
XUeWFkdrXpuzz5U4SDK5nKS3DG9Iun1L+hbs420cYgr5nX7aWz6Sy489Xh3XX/lYKLTNp6eCLsjK
mh7/jOmnSp5xR3exATW+mFof1qyKy1dSiwutkw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SqApNXbpr2t7CC7d8fZtb/xfvJmD05W1Z/f4uy/y5KP9KgyfkoacwJsu7Z96Kxnh28hTVbUr+XCw
DO4TkKolZH+V0q8mx4RozLHwDdxV51gziP5JyL95YBlj+cgGTtW8Pp1+IESS6yN8I9SYCcCM7+5s
3ZXm7KCHYFL8vQZS7AI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V+dXXGh8I0uauCzKNCpPJ8GCO+C5LCBRq6KgtN6MzYYF6bEUw/apajafXOWljGHKm7jCKmjn+5M+
NNKXVrVygNHMLjHpm8oKF1RbXBR8feDq89OnxkWRacklRkf2oM77jMJsLKx3zlx41FTEYDx6yQMR
95ZnhrFZ1TzkZx8Omgii6kpyCzK5uVq04RJnBWNpTy7LCQJWV/g20TeaWZusSbByV89fjKbZQcNn
FxDuOF5B99SmmbtLmcEW63PpZwd4ZehH7S5S+iSxshNAZppS7YcXwttXLfweRYVaQJXBHP3TI37O
w53geuCPoq+cQXG6qZ1Tl335vLK7ogAkSQuBfQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20960)
`protect data_block
FcVWi0vTfK0FCtktTreLFEotoKZRsQJ8TzzL+Ix6AUkIN7fQ8JpKeLWVYiGW/zV1/GEyEnox7r/x
7oeGmcMRmiWJCDQ76l6qzWA/0CoLR6L8AKEHk5H3anQKJypZ0ojenVcgUsCi6Z4Mj+JCddThYVSZ
moZeZQiD0NkMQHpL1/3dty//uISHqjeclzPZbcEwGQdVG7hQi9Te0ppSatyAHZRGLH+ufcCde6bl
EcrbX7HLpekmLcSF2Wz80tazJWIsqIIJXqkAVj5EI2mtb4oHCR1oDn4HKl47d32PhcCWypcqtuIa
oG7YXFtTTV9q6L2mexASp2qe44SRfDlksZxq3vWrocOYlziY4+081KRdtYGmKmya63MHWFwumWnt
e1DKvmjOC0NuFe9emdJeJTWx9zl7OnbIPAGj0tArIC4b0mfGWjyhVIspLOaRlm0M5t+telRj47y+
YCJAyd85yv4CtSm1EUu0pAFDHdCbaSXRX5OYdm5yvIojDCko0LILpFaI9sGkMMTs4+A287f7snkj
ZVTSE3nk/hvB90EzrRmPphVUwppDXWhskmVcMMGBZyDocPbdrgNJkpi1V13N4Si95SbAdT4LioYg
lRST/Y8XITHrM3oUgpaGieutTru3SVrRiMrY6LHPnb4bnYoKOGZrw3TZKjCOWtGteDAUNmJlR9GE
fGclo603mErglhBQoUMOlL8bUx+2/X0g/cnzi4Dd/YtYpztJBqbH3objkGs4EXOlOxtEhuKIToZE
+oN4J9ENizV2JAWEMpRQEIONYUnwmw+hxNCpx8A+BHI3fVKEuIseudBjJFTLpG/lNRbdI7EvX62b
4wh9L+qqcET0nkYOSDdB9TepSnR3rmQgbcd5IrbvlEttkSPlkdmtQOozMM0d/Pr6b1i4QRUm0mIc
xF0xFnddvTzQmggqLX18Lat2Dax3fJAgShw2ca9/xuhwwR+azImhRbwIZm5aeXPEpYwYmZ6ND5c1
fJwYGOyysohRISHiQE1iWeaRw2ACkub3SEJyywiJMd+1ufE1WjE/QGOm9W8GmzTZQTutTRGqQYmY
t+I/2QTdJQ++hyVXRC1QWiQYy4XCdrxa37Wizj/uYIWMhnlufZB4M6YO4N9C5hqrw4OBpyU2ElYS
dAoF4CaWnBj+/6eSYFZIIhjGjWdTtRGssw14hXpTJde6AAdFQqf387LUs7H6can7pFWFz75tclVH
jnTqk0IB+gm9+fOt2m5OKd+BSAykbCPiYU6yRk19IjbixMvm/Hx7//L094o1A0IHICCmGJ64KfvG
N5wloBRWt+LCGiUrpFbI+okw6XBUn3Sw1L9ben0b/HzehYIp2GTYTfqYLkQhQFYhOVcagsTcCQD/
ByRtYP1jARSYj4YHQcpD0VI8tmF3lMBHxA7hYfdgTznb2m3GtUmEwbtgkPvp/O8yfUaVxV+rNd+6
Wxuf423ibKtnrbSKDdPGqbbRpq+mto92z0APy6UoRtWZL835nMIX9MiqKJV83ekk2u0X/XT/3XbU
Kb+vJX0R0qOul06Ylfrr1HhMvGptTcvAdciybk1w2JJ2kxGSTYsnttWKqLM7Gar8COtFP+D0usXz
OyuG5F+j/EFendDVqkTGiaNER9rvrMorEh4g0jMKylSo3WzSJOeb8ADv/A34RCYbDyXruJhTigff
wWJi6Igy3UQ4xO1iRJlomfzaWn3b9cqMbyu8cwr2DWzXGF3iYHwau/JKOW2Dqw8hcaHpSj9jOs3F
YXR6dXljFRwj3klABUbR+yWLCYS4PDZW29eYe81gDwm8aWtOgAtyzIfSrDwnEJmeY9dZIreVuzIA
IpKz+rFqOF1ClPiD3Ha75Yi6lwHgUnoG2Xz9JAA0C0F92+1bz+GVZzuvrZc7mXkeSKv/lA2+ulcL
gUB28Ikzm2sTKUPCr9EpR4wCxJdZmk7Jzltet4I77u3dPxJaEs2tJIZ3OnszRulcIxB9QXC7mI7U
/1NrhrIiA9BzrVujgeFJLwh1T7pS2kK9hu13Ome8QUdAYcd33NMKOjMquzZsqL4iOfinIuqK9TzJ
50Iy0Ez1SJXirpeO8Vw529aeIqVbQViFvRwjW76fvdd1YKGO4uAp9JIQ+4PVxfdf/duYiwVBcNUO
gwra11KR8hElaT/EbFjdenFTnHQ3FcAvOxdphtjZMNICyal36cpl1df68CL+6KqbNN+meh1x3sMi
KLhwd/78ZWed58udbwPVz387Ls1P3uXz/Jm4gvOcaTZaUgBYndKx+AntCzvsn4lfrycf1qbY0r47
yYk2gcvLWxpAxj/D6prJRsdqka49Fd3ciR7O0VqspAOb6gANY1W0UYd2v71qJDTMeP+xYo3GJATO
J9H/L8xOipPiHL+Z+/XhvWhz6Tit5qt9uRX98M5prLqtjc668XcZVPbGqQ8GDbwYVUtulQlGAN12
wRvX5AYXe7Mb8wgmI8SVsM+Jo6Hv4hTTItJqOepeYkjoDFj+QSKUzUJ1SoLdgTl8HABQBBLVwvJM
tPSCx28Iq6b1xrP8CJ5iHXhD8SzuTPbG85md8V2xfRFHeFqPzlW+6BgX/b0UndgW6oz4BoMnB4d8
q9nMcSN5GeKw7pKZNGvriJ0bmLmpiZ5QqUJLeyk1AEH+VAbvssRBRcFMHlX0YfuWjzWLlmjbClMd
7JgqOrkdWuVpYnQEL2ZdIGHsPHRi3I+kjyqodAGvViKKwW859YDu/d5dbBvimi+HgWr42YZslLlH
5zRmyHK+qsjq7Nq32i+WA4cZSwMReU5AAtvzTqTIgh4cfKQ9xdoKd6kuW8Q0RRoSappi2Oq7bIBb
vZ7o+49iv9Y9w213pz16xdePH48cJv2XIXadoe287Q8trCkYxKHRtd+VAHLFvA9VY5z6HX1DUjJP
F6tfSYZSfvAaluFI6LWfB9Vi+oJbtxTxH+cvIIsSVaA9kw7DJnh1itEg20tOzfBClk1CcU9lPTzA
0g2m01QssDtK7H/3e97Er6anKZgDN9zGNgeGTYjrMSxw6CYosyM3cf3RI8XpNAtDPM3+/U4okth7
wU8FaTCIsQ71XI3Owf6uh6M+zY3n/h4TA19zOKJaxgDzdghoXLFyWU71iuU7Yo3npPKRL3g9euhC
QLFrsiNWP7r/qWXuXuI7a7QTQCoVRZpgTJJ+JZ/ZGnyPQeoalNZelDnDauJeTUHHTHx3snVVRTXZ
4pJ1/PpR4nAicek61qJd6bixcepw59s6fa0V5New/jiX2dqFRGMwnFR7Bvm7E6rbRVPrbZdAOWB4
qdW8yJqS7XLziRQNv4c8jPALN+M3xXXIihmeN5j9k+oP181gDdhb8HBtxymmbLKe0REWYB58i6Og
OKX0HBp4yhPTJ9xNtB1R/bXfz8HFnnAiekB9EWqVjb4XMRfu95S1BzecfI4KBL3MaURn22Yz58dA
HOE937HEyFV44UETAr7iOoZnZb06vSAW9H6m0HbQOMaFqxs40/RwWSa3WsxEKQe1OPehftTyqBcb
Cht4fyW/pnpkmCBcvPeOm7vvJjVLr+d8SogYi/NEz9APsKEgDhs3XhibSrGXkVE9aBVUFCg0dleD
DZs1BMv9YjVIISnpOeESE98B84yrDlDwHK1QLdttr+7MD/+nvxSL515Te4fBPHrO93Fdpu3WcvGx
jyXoWESqokXw4jD0WegFx4gKnc7ifhhWaepjR+JoDacsTbgVIxEziyex4Yanmm6P6bgLGs1C1rIO
reihraD4Kg0WPVZuP7cW3+ASWlJg537k1FwGGBfxq6MbuBGjEN8ZTFxFI6tzWFZtXipe/riqnuAT
2QmKalRC56vdmJoIDmy/77mz7SuVqA02RFLeI1Ao9BBOoiezIWQH3wfNgPAk8BpptVct3L3R4cgi
rKZtaJmrtqM7sPZn8HBHTH/UvF6XMUCu9ctV+MajQT4bKbyw+qi4FzyVjRXW0tXvb76RyN/Kj9M6
5g3/WQTVDFb4dCuMboqft0Hxv28ryEtXSf+DMuulmUwWKee74M+InsbQKu6i9Zz2sKi7FZNakYAM
ddliZyedNBOIfHesPx1J223HtndOybZ2MfOOjoOVCHGssDEUsJuHzTfDAhYwiAGQ0DZxf+DeUPrN
1kv+yGEenhmL4WuwFY7O5Esw4xGtNgP8igcke03PSXKf0Y23+mRi5LnTLYpI/Ujgk05KQUnDyyXo
afCZPyMZ63M6yyyOeXuimqHgkdgdvzYdZ0ye9RfuuIzwVry4gUoP9slRyz3fLLd+XdPYFrlSpn7e
MFONU2t/rQM7KSuM5fFhFdyCB9kZG3C0rl4GZspH8PPwgZSlCwygWlPi1l8+jco4p7KYgss4Q5QZ
BP1n0v6ps9oOA53Mf/PkGdpIvn892q7yD5DVJfCACTzDxaIXhPuh1GsORYmR/XUMgCgJcHLVp2xF
L0siNSsPuxfSx07ZGAscSM6I2CvqRUq2zVFqCmQHtkpvjBk1vyK7cU2iJBXSMbYvWsTLjtLJVV6m
VloL2nZsWeg7MGmLKbYMTzq2zepIsu895owR5dSOvgcVaH7KHjQX6d/MCBiY2wHL4oVsE0yOhnxo
3EUROmcd071P6enhrVlvlGw3BA1JTFMfZpLNUY/NOwkBNaMpzGhG8+wv3cI8nFBsLpO5o+Gjg8tK
IIc2em78aiPpMK7RyqXryQ7KZxRwOqs//WcS7T+B1Zir6/kkYMKy0UM1LRrumQcI2NkzQWllXnG7
v7cZfNpJ7TL1p6G3TR+uIX6YOzG4Cphc22srucwnCS3FIQ0+ofw9BMxu4stQd2duahJwe9ey0oYK
LKoxBwbry3B6yfhSLbA8D9Y3+CM5ZbGDlR2hOVHYWO0ODWZc8UKp2G0Z/6M7z8YmHX2FOc+7Cy5s
IXsQuzjvdkjpsRHxw7KXwYhVuxkZhDkcVvX4ka5CSLCZZet+f5tfm3YxxK4bSQZGtwvMC/FMjWSa
iONcH+U4uKeSjCOdrPyG2QSbPtJd52AxpSqN5kwykOiNBejknT+VwyeuU/lHdrGIWKl6Dd+pm6A0
P9zH7e8XDVu5zpUJUmrGajGtYBL260tLLaSyGmMk2yRGFIEBRyo2DNOBE1mKg9k0eq/MoS48M7AH
1GUKDuIOB7UxgkZjdOY8RpdrYhzzRv6nCqA0paWBdYgsbY8+fkB0D/i9tNzzryNgQpMYMX5nw/f6
ch9WDW9r7pXACa5xjNVcs+sRyGr8Q9EJHCVpp38J57c7X7QUETmrnGLPrKtvGD+0siViRaCt3cba
ZhrriIt7xpbpQ94BFJBvSA6S/h4Wu5lXLcW5owjf/OEa5EPE03Mjn1cO9MrHGh6aXT3NAY+hq3Dq
lpEzikjlze3BgIRhXOAHa8gFCA4SzY1USjEDQy55Vhx6+Bkf88bGXhwt5lnYN366snT+MjY0OcOM
P9Jq/IqtWH+uN6TqSzoN3235O2nUPbUdxN7oiDnABJM1hmIUy+NZkAnlJJcjFGjBV2krAFJA0DYx
W9dZb8vNvx/OKzekJopi0c62wV4JF940W3jGANIAA7+cuyMBYiGdln+ki808U4yZqX70JRD81c3m
vPsw+iFUqNz1s3HCT2tHDzb1Vg69iyI3b8aAS0w0PvwLPWymOWeHj2zXB9XTN56+x1s0Rk4volkN
UzQIDGKLbET3KuHw0ZtwDmKg0M4KAzS1GqDOi9E2DY82fVJG3pPzQE6ydJuaD7h4L1X+GDygaVjH
s6z06bMZUtclWsANFzGb5m3UYa6YKDuWSpuiNa1kHmQ+RXvHxASheSPg001URqXYRJAoLLZ8J/Lg
UyEmw0/vy5PCWXnJQEfICoR+xnZJn9KoZEOYwy6Pjq60bT35puBUeHj0tBTAJq02mnABQp1AIsM1
AXax1W3m2ZeEe8APeqokKdkIwPzmLjhtbwfWRdFClKgfe1I4KSmR7CkGlIQLNzXUQw+/aZBn27Gf
0Xp7pWv/4/KdAQUanYMp+qHrIIFVs9kHLOr+TVDCQTeewLfhPKtI++8JOiB1Cup+BhbgGLOL2eSB
6/OwQf6k+NW4aOoX4EUi69/97/0CsLwH1dVIqfgTSwDk7P9Q6TIubU8jlH4v0o9hsSTO8+jl8O/D
TvzKDRrUmFUKLqxBuR35263ruGLL8qtFueEE9+7VO+RZlwpAPS1w8laZI2pEXXn2h/SoWNgc1OLz
ZhX3Gp66DsCheZmleB0VIoP5++Qp/in2t/D9jCb/5ZIElksyTL7a/qqdLLNxJTlhpU2iIsLuNGMu
1JBSa5mp9XYcMw2q8g9TzgIc/HrwUAxUwe9zy5hkh54Xp1sZJM8cxKXc9wPZe0zJrZ5FwkLAcAvU
byxdjnMbpRsIhcDGgsDUVQ1ODpn7/jkVviF3ILDBSLhdlIv8SsQNds861zzvSTVebIiezZc32IyT
GRlsffV49AZqZ72yp5WpsppJSy0CgoASXYLwB9nRCBBkAQvMU5vDe5YqhKWPezy1xCW8a9A9o3Qc
xbsDU4c59baOJrMPPYfLYw8//QbQQZ7qFSF92vePUU6ilCKHf87Di0kmBAHjGaN7DzdZxyH0H5m1
fXn7W//VwMXZjASLz2XvPAWagk6LlWT6di4vtM5g1q8wRI6o2cS0bfngYpphDYeuuu3VbZfpid5I
eiq80aWxLVZ7libkWD4Py4AdUWxBIqr0n5ioN1xtYQgW1Z0RYbFs8ztZ66P3BnE7JHlOLpszWXOK
ZxPiZ2cUYZv4Qsix21Vl5cwiHZxWM6cXE+Z1sMMAU3372Kw3iojUl2zYo9TyZJI81bqQ0AB0bWXn
j7F6VrDzicyGZLUXmKTFK2+WHkE7SsYcO1vGY0uXeFN9qnzpeuW1cYhNpqxyK7vgacfEhlaIo3uN
koPX6NRbUfdU5Orujp+k0ePS1roVqkW+39a1mSmDSOJcRUjyeLr4/Ih6DxPrI5Iy9T1yHes7ImH3
UvAcexmMth0+UPb1V4Nts+KEc6rZu7jFA583JPFcm79r+A086d23shhn7lkJkgAJaxlHHHJrvRSt
BND+4+dxUsZRzApd6nrFn5ovgmvsVBPoHB123uqdDwHecAtRwGQxQK9xFAFhVgI16vOGzZBXCSQ7
w4rMeVijaumslhbWfAuydUYEyxPRdv0r6UJ7BeaRRUWuomBtcXqaOB9Er1ANnofYFRBSVVpAYchS
StNhIPG5y1VCphZhI9RLoiFTWLjTiXHrF39Yv7d3yt5D7iQNvRvKJffXTWQPJfkAjmW5XXviR6B/
hTgxKf4yypoVBs8KOpeXPoJXogD6lS8xDyE5VcNRuD5NffM3S3GqqJc5O8fcgFrWmJRh1ZBJWw6K
kfH9ZleV0j87UEz481iPdetyiT4Yn/PoZ88BW/qovA+Z9pC1ymwS5kE9l68jgVrHad2OhZ+RHLLR
M58UrKzznmRABtsjLwl9tVy15knVbRfKWtW9rsd4pb3xR/tcANWsYi6nWNP5lWwZbfNGpO9gI6hU
yZkAKong2q5BESz+RYJCyE2pnFwf1dmahgXIn05pFA7mgXhEBTcVKnFSEz6LJWvPKIWlPOGmzEje
zyRFjvkSUXLn3Xr+R0Sl6vMiMs6L6Qheaj3h4ofxh1usu+l6UIApti1gYuzSQ8bU2BNrsvASQqQQ
MKZiC5qP8eiFuQDMMdM21hWlkz7kZq8oTDOF8QAmtE13c87iBUq0pz0/1nWAv8vj2Gq73Hr4SqZh
phnwB340BebUmI3Exyt3b68dnwQw5d3o0UH19+V290RD22neVmsohZZ30AApMmYFoxK6pMuHYtTL
1nd8YuYh0rgGakvJLpbO4wI7nOsZob3wpPHb+WX86PjbMO6Os/3aHOWDEmMygfCRniLG5pTcpytf
87q1KdZBMV3KCcDbDCXpWskEVZnZjP19sIwgkRPcp7/QtqYKAwdLkb3oDw3kMRzkUTsdd8IPAOpc
QJuoFQwS90JpaC8EKfWczhLnstA4bsShaIqgWTF9V2CGiGvEuXPR8bFC7QiXT1gsn6qdzr4H2Ca9
n2edDjR6hr52imT2n+DKhsDhq6Q7X6qoAKCZWe3hNApvUDmkfx0QTsxWn0eg5rnr1hrXmMh07pNz
dcIGNQOtw226Za6f+AHgV8riEtIHxkK1RJ1eOvAKygSuFazSJf3ISL6GyPogl+914hoNG2wdJO0q
JiQ1uvRsRsnPPSooRQQyjBsuMGpNTo0HlfZCXL8DTWtvkfiwhTKtMXgk5meGrqLtk2b6BwSZP3pH
t5zWKGc327eoK3aV5DcG8NC+kmmvSGW+Cqa1xn7T5fFCGzCprshVCTm5FHkNFvSbKVponbXSJnxz
ZDRdNbHHa/wwpvCS3InITNXk7E2ZpjG/ANC8m7WR6Cgr/A4OXhU2NxdpgVskCR2hIogU7uv/ofh6
IUSrnvuyX0LrRpIGmdJxTRhf7nR+t9j14EvWU5IPeyP2bsvdPjLW5N/Uf2ZYArpsXO8Cr8fjPr+n
efWD3+74zi4nta+xxzLFSRlT6Ys2PiuytV/Y103+Tb0yXmRikLOf5cCtmSr22IOa+maXFVpLfeTx
L2EoZFsgwwdna2k8WDS/qyVneS3BSIjQtwz4BQ1msr8QP2Qzl2v2StIv91gXAhnUhKDtb2gkoccb
4yK9UGloq8JQaL+tRBgSGoJXEZL7HxJOnzu/M1SbHZu/kS5K0rxxeuvyL4inPfPc79RQbUZfRWne
Vdrk5pASLn+P9EM4iJy7u7HGK0kejI8ZkvwLTC3NHX2u7Y1CLfsjIhXArxejaUMkRxUHjHJHAW0G
4SYhUiXWKIumvAF68QCc2acCbL2niUFE30Q5i81nNQTwb1YPFZJ45f2MuC/ZdksGy6Sxqr+BdPGd
Re9d66TVsx2VKVKs41b1EmdSRCnz26lplzn8RqYiOlDVIJr7AlGieKwLDuscb9+CNx5unGKTDCLN
sl8cvv8BqufBzBn83pL3K2OMVf5bUfftVxnAVwGfvQtv6nxnsCMTMK9dNRFPJwOg3StHlNAXfDOf
+VQ5Sn6oPbC0SK9ea5CaaXTKiSlVBl1JAFMAReCTJv58nDFlisJg2yvUcCQcLtO77lxgbuH1jgcW
IEBczKGfDVh53nQ0OMPlF2Btl1jrLVenWMOKrURfjhYj2j54y3iLAmwDW8Jkrwj2WhOHyC5m+T9s
2D+7+pR6sP1bttghY3Cukal53Ord7yHYPP82wcI0AP7QcVY2EsmiT4jy/VW+A/vPwz2nofk2X1Lf
4u+wLyL/bIlh/t7JI6y2hBjhenVf9LiDZN4DfeUEYm4fuz5rcHm7H0QVquOKjH5aztHfnILTVIqw
iIbnexVkMAZV00+zCMVVB4wgNTDAXzzPJgj2iETnvK0VWMZXJuo8OuofemI7P8fVpjtcLKfIE0LS
8QAFzUo27u+OVrLh83qpyh7n/i59aBCMC8rQm33XCFcZkxVshCpnL+6VSCxsy/PZYIz5PyeYFeDJ
Go3lYWdTMdLdrMF3vxM0dOKSJlx3FkoH0EfB6n/OsO1X6PRlfncrqg5zYLuxdHKdX5k83kTqmb5q
Y4oOpCmSEh4fD4a7wOZ5AJHGGdTtaD4lVKI5mZV8366Bz1wmpOfuv841ozQWCd5qY2oImS+Fl5tt
eEVZVG3iH8+TN+TEYxN/pVoXPkaQt4vkeQOtbXGxWDETdXYow9Hg2zLROjvwnbTAUp2T+EFXqQNw
9oU6YgJ2ww+Wy2JbWuoLFzqg6xKZfJrsUJ23+oDsMjl+FofR5wR985OTiTC1aggxN5Q1CN0mgiAz
lh57E/AR6LJtzBIHi1mEffR3Y1Ce3l+HhRZVoWaWje3ziIr1rpUJYbezc+M5mwW4V/MKJSW6+mqo
SaVDfKyat+Nm+Zhy/Y7rH7zFUeAD3eFVCFKU8BKGPMysLwFJ6WSyy9gvhHY+JoLIwI3DIQgaP4Kh
5mbm50uvIFRgTt2AiXKbaODTKc120/A8WPbup4donH0SOcr4R4NZoI9f4STqtvy1qwUripaEdQwR
x0w2s+u7Se7F5NQ18R4IKumEv4+m+N6ZiN/vF+xYUBLPrJJl94iXAcpN1kri1PYt0WPROHwUL1J+
NzI3VMwcqstvkmZAsas/I+RharznN5eERWPfIhdSGjXivCG87m+YUh3ie6QruOVn0IIuzA9LWKUF
i778G6vo9oIgYr7ja25NYso4n4Qesbl+DJ4X1l1/T+ffdRwrqJFMqeq8nRIqpQmW9CFLHChagrNS
/eQxc2v0LarC+tNHav8RflEkAshgaJQ2KJSKmNVLvAsme+Q8Jk6w85WapCFLJG4YJjT7ySy19KFy
9MAkmeRqHyP+6ycVsstuIpyIm+HZSGsr4BRdeVn13XRVYiqwxC3We3vlEjc2WFWHfSO80I96c/bQ
J7ZefnnL74mgp2xClrNpt8PtRJHOOzVtO60bicOUCCbiMRxD8227rNXa0Jb4E4axPZZQqmNi9gJ5
AiJ200B/5TD7H1NKCDKvw1hXrpavPHzlTCrU6w2Js2zlXAeeXhN1D8CoC5togWPSSWTAvlKw2lR1
9RduYNoCNNZ15Kor1q+sZ/7e/EAWDOk0mjjjKEtYGlwnMtFAjUezLZTrSg7oXjdkVlb12FS8wEad
v2UrZcnB2UxyTIVNPfTGATZCMfPlQdT2Veru3HmTkzGSwJPVEPOIm78igKCFnzzj5iby92/aDWH2
jgQbHoNeVxgeFF4A5iGbbiSNfao4musACpL9Ozr64lAjPWmA4qX1KBGpEJqpmPv9cQsuzbxb9kYd
q7TUC4KGaMfPFmwC9O11ezw/BHxqGEBkC1Oq6kzw8Sv1b96fjrCVF07dN5q0g1qBBPhKBrYba8cg
P6qKoVLC29e70r3NwHpXljQQebLe8ulPSzPs6ILHMhtyRPwf/OUTxxlMTqHDDcPI2W5FIpsO1qSA
nbmeANb4KwDcCUdOMo9/KlTHQnSs3X9p8ifcsxCfHSwv1lbJ+sdta8MYHNm3928XFKItphCZN10E
NIabbkvOQzuF8A+6lsLrqKt0sEUfcGd85TLaDwzE1wElawMO/su/6Z6CqJVuDZcPkT1vJxfPACT3
8lN5DQY/GgJLqbgT8zsT91i2vrbzBL4899gzEwJrsg8UvH6SFFp0ttb/ZTdL7FY1MzFjAoR6i6Wj
Ukf1+AtH9TYZ8d1FDBdkkEfTrm70Dc8sveUruOl7OCTtmBrvayKCeyxiV73/I0Vr/dMtZslX06d8
4L00WN/YBTHi3EqupruDjAq05IBV4/o79ppL9prFyj3v25BcVdNAeV7N6Pg91ADqP06R9B948oRu
yJkOoaTLu4eGyJTI5JO6V+aezNiPDXH9wsO4FJrwhovFkkL0gj7xOQjxpVgeJDRh/LwNrJk66BwK
8oslynl5w8bMw5Dof1dpK4W9xbOVbaRjZbGlG4DDV87BaE1+o1Nd4Y1VaN+G5QyxIVx1Ja17i9pY
6tAq2fysxomkzl6crO3qzi5uYke5CnFnNTlNpaZyPJQi47fNAZ4zcmq87128Fscyo09EWvdFAMZ/
NLuGxvXQPCSPqgMQfe3ZB+S/WnBKAW4+qlvo18zTyYuz1olTO0HcQ1b9V8Zk1KKGzz887EKXP18i
ASekZZovCvmoNWZlkYsMjDcqq3a9CayNvNdtosMNlN8qhw8cDOkHAiWCOi0ypSbxZ0LJl04C81Kh
R1AQv6AwsvjvNVE7GIbUjfh/ug8/PhNtb5+GfQ+JwTQsO15iCmR7QYHfPLjrH89+hHc4i6Le9SCw
QvcwwpGmjiSpcqn/1kFGP84Raul+TJ0OMppU8crB9tLePAtPEuoSGcEb7hHVu8BxRnEvyD0ZQdrc
6O1FoH5ruTW/5gTSbxVj5LRKFAxiwk5KZLeSUQKRzEb35Rwtf8k16xLeuyrVMl2J6frk5MGwfuDE
Y3p7nR0vpAZpFfcCZDOu7XNfHSDFQCBL8N4FKgNr+i8Psp+8SIgCn1+Jx1sMbzklJrNwjT5hrWGY
SAtJUjT4aIU/IBmx9JXoMn/jB05gCyrrevmdIFsVBrS0BIP0DalH+GS1y7RcT3lsrpOrTYd3EWV6
4kOLbMYmLOF+b0NRzIoUpoKNn7UPWmKL7nrJPdPAbUW19oY7FlPiQ3zHhgYWo0UkvDLiEHENN2CG
0a48O+Fca5WjygvatrmWUyks9a2ZkFf2SwGGAHGcsXBEvgwAMEbojrfe9KbzY3xMfqPocWYRczo+
bxLkF9Z+mVm0V4/iOdsXWodT6N8Xjp7HyhCfhnIh8UPNsL0kmOeaIuz4e7p4BaqNEY1aQatnfXXE
obh8ygMmrzILfq3bbhZY3mdMYE7kIBpExk3Z0Rb23u7dV5Pv0sNHX9uXUTM9NoqrIfUD6k0Uf59n
PQvfeY1yhqIaPg7E1+vF86wZSH04feUmNHLlv6FGPRw4KklEmYeNlu+EOgKqW449mS6TZNQhtucK
uvI5nvfbMQzNbPFZ6pML4x/zgauuK0F6R8BKwjB5g5uDawPFiTLyehK1U3gzyKykRTnwnT290Sgo
gvsyxB1CiTu1lix8XoJ8gUAFR/DRU8il4R8+AEzHhr2Fanj0eDc9hywyxClScoR1gSOUdcOhlGsy
2zYypriOroXScqNhf8diFyZeXtr5ovPmYY+aAgufUbxgQveLemIo4Dz1zWxqljIHZrfgZbaG+8Kl
3dixt57492HedGZqfDmeH5/FzPVZCWn4Qdw0zU0clZh8xH/aYpFBEat97AFp5nc89K2XYUf3URN8
ak42Ox/tVShj72trIcg+BLgv6QodLf7HGURdZEEBMq0aIC5yLIJ5R50v2CWC+JB7f1Dr965GniM3
DxqybbWV3ZMdIeq+wGofF5i2hhe2OHpxbtRV7CVG4mrTUzmCKW6q09hjQWy40emJz/Re9GAjBk3d
fm5K5mvKAg0VZaw3brEKDjKR53cGDUoo4u40TeGMcYkpHo9xKYucv4soVbTpw4IShMfW7+Q8U32J
ggeYBa0uk3bU400tN1WD496l1sDopq8Udd6w9tMDjigJMpw5I97gXomuq96fURQs5RC/N/LM5B59
fAfUC9lanJvyfevA2/LQy5uiqmIIRqcy+hY9R9rjdxe/QmBfhQ6Ra9fLyP2SQcbt7H//uEcyoI9r
mwWrkZ5njrm+3KxrrVkMbJcckD8HkKIw9Q0NGLskkGxbfyb4u7glFbg9VDWK0F8dfyWMoZQ+GBe2
fckOrkXEnUaiLpI94OVJXCPSQncdzbuKkmVwVGcSU8/pegCA0pcJUT4+IUeEFAtVE+VjvpWdaCbp
9Bo5sk7LNzrmNIuHw5TvRudOkELe1SWDGA0HapjcsNVPx5Wwq3Vzo8CwTwz5kd9iSZ648Pt+ukAl
cyHvcXOn1EO5tuZE7qkwlzBymVgwsVgRqkasSUAFfcEz7ATREMikpWNu2DM3K4Vcp1eoQQYkEADs
y3RYgdcA1OUTZuITgROlqDomx61q6mG4U0EkPnLUsadTBNHW7uHAoquZfDfWA7Fe1QsMxf03GQCP
x1YpfnzSU2reyRXjFSat7MQB8jGrjz0m/3BlSLN7vZULH1CayLhZpeEo2EmPy/IwXNHhZ9+Po1Yu
rBTTlHe5KogVgAXMdecW67x6xtzWrmRZ2IiNuglsIerlKw6xTXjpqTWfMKqfPmWPmkwXqFH1wgh9
ziKz87ZZiv7bab0i9CdPzSO13EApPyCUAsasrCtTfz4T7Zw5QEh7C9r2t+1rbnXJC2bph8N6NgaX
4gyw4fa7oLTYp50fYj5CvNc87dd+wpKC4BEkRChtbDnbLXltQth4SuMjn+hdiW0rUG4GNVQGBHvS
SsNMBFQhwSzsx2FavqOXvQ5q/lansASdSLzxk3fvbdQC3MeSriqWddaRiKkGZrj2C8Eq3UpKloW0
u5F5SaPZb3ZEfbcXOOy2Ps51Tnaaf1+YA668fBc3fEZLzhNZ7kFwXazONP7ayFH0kpARrpGWSGmN
2StdaVNERFkMFHRhztvaXlZxpkzNWbZoCWMSPfas6VvobpgUEkyQh8vrSfDwEzv2AwdPhRodxACB
Cp+2ZGLlOkuEC5B9F2R4OLi/ucH7hVJwrorlEu+qJRrqqgDuDJ66S0E4rbhz83cIgG+D3Tfvfo6P
NHCfM2SvdElJTrnqfgf1SozweQcun9HLof+pPgvZyj6oWCFA9hccTYV2GOCiRdWfH3hwfiNckVMA
BENO9rS3tILh/j63jExs/h3XPZE/w9AMgvU8SEUPXWQYu9Bo4rHqH7f6CBaOZgXAzbl5Vx2OZYUi
9lQK/Z9K83zVos6uYF5CbPUwWjaA5GHuTrgO4uwmj0s6vRfeBZFFlM6tjm0lm6lePz1Xp5AfGA7E
TWdHinVCSKIHh7sYarltOSvaJRE9ocm8vqszj55wIskoVxseZ5ltlNtjaDIh+Ko922xyX6y4iUEI
jjue56H/jT+uymGDh7OcaGW0uxvCzxiGws6Axfz0NFiOjMFn1X5+WLtaQsVRhpTdlY6Qxcs45L3o
fLu/xhZjgNjvxNkhkuDFSIGrOM7o3y8LMmnI9CCPldbSi3s9BXzjsU33xKMminXD6BZi8QgpHdNz
UcYGFYtZuo9PPjhE0D9Rir32sD+Q9EIJavoxxF2E8SCTcqwPD8HVKIueRnEPeTVtEXrOG4IWqag7
aLMXM7FmsHkXmiL+X58u9XAAudELIIjCrUfIA88l2uTVTF1KIuIzzfmbYC8mCiNe8EST8QCJ897Y
rxyQp87XYUbQRT7hHTH6A50k6Dm6sDDP0cxRIifZaoAzC6qwCjVfd+KJK9v0EhuCyX/MZ1jbmC5N
w2uB6HPJvF/4m9DgN4mj0gWAh/MC+1MTCs6GgF+7KTvNEJ/QbkpusIrW5q9Q7PwvpSEr4ET9zPRz
0r6cy7GVXAx74ccEHGckWqYTslGlQHjwPyPqGbmiJjTPkoU1sESCGczIZbXs/7xhvQwxG0tUWsEV
mBdJLA8tcvc722KxwoVGA9EfzI9p86sPO4Z0VkCj3f4F0k4Y9y46H9szkxcwwHWpMg/uh8ZG6ZSt
/yhT74edM63AkXnXeya565A2tHwX+zz7cer1UDH5rAd9yXIt/XkqE/Eg25FWUinqZqrrLnz/9uoo
BEvrYxanCk4e4i/UgIvkiuL/fVAB99WHw80TRXIFpQBJPEGXoy83Lx/uW+jt8g6rANImU4cqrzEU
lgpiKRQqL/rxJ4uTKs2iZkg8PFqsDrO4ekDrpYnCWRA1X9s9SNHSOMFeLbyP1s19bb215f7yZ4we
ut327VDoZYkSe9ze3u385ryRhwc1lEsitqEDoUebpYTwS63zKYNnbHx77FeEyqsDkNyAqdgq9GYj
zHAAzR03Jovpzvkb8TdwkpBBfqUPZYETTlC9uV5iPauQ/lgDh5tSLD6eHYc71zglgbKSNBIzcAk+
I93Rpb1cA8bOBZ3NGfghaY92sFKPVQiFSMFsV0Qd1n7Pjt46xElPIS1iKI0jJocFtPhJkPVAUZhD
6bDvmS0k9K6koG+Sf+yY/UkwACaelDwZjVjRAu3G84WLVWebPhB4DgKmodJFLnOxhKND4odHLQGm
LTMBHgxN3eXmXvWkADQKfVg9xp9zsmpe75sVj9Pw3+CTE5WpzCMDfdVTBG7GByXMTTplM/xJiWP5
3GShkw9MqOhSr+FTDWFrRm5cRSFkOvsEKK+LJdyF2LFPSM5LEZnqaCXcihSYju36bndVOdz9MRuC
7gYKUDxSwH3wNqlZXDMyXlK6AEuf1wzmfFLL916OyAZe781gl/3Dt0MdRf6MtaFlhW5Qo00olst1
JXc85XyH1Qrq5r3eNTaPE6KJdZi70TFl/Dpsp390GsacLdZiGpLI2GQHE4zvFtCdIBctap4dKf99
y8R8qaZaDV4lI6mPdi3Ho9bpcFEJrbyrxIRJzjnQMhOn71HEPYCIl0mJS5qWjL4FSLebCB8UMZoX
gFlhc9d31kiBiFa+4YTgQSUuI9Qywc5jPsUQ2P8nj2hSSrd8xlwOqqwkVaxB2jtaZsyTzbQ0P2F0
2vzox/0ZTEWv5bONsEJtSAK1PgpYvD92gKDye64J4RhfJSVcqQrnoUFIj/HtLHfmIlqn61QpUfq1
KTf+WD+48hQrujffb6kyFwdgNkf2dPlDgRCr1JwIxJo9Tiqh5Wtp1fTo9B4CDdziSiSNX0RcoWIS
o0vlxxmzYg+8GVLRRVe6ZS+1Ni+9CmIjDuL7r/H0RYMttqdQnQHQcf+8kyeD7E0pbMWvwHN1b1Mv
k6a6fW8FLafHXzYgPXP7l+0rm9vc7YR6kvEBFqX5022Ajostr1lTM6ST6Rv8CMOAO7cOoqJjq8gV
TZV/yvh7stC626i8N2l41cQzO7aYQk+iLcXKRjhMM3vEYf53nJH99l4mDEDTWr3Qgn6wwnP/bDEp
8wGQ9iB0F1lOheFjYAj01bXsVF2TROJcCQSEGRXg0KxtSpbp2VAOFU8xsF598i/IzNLYcVKlssmf
8UJWTeMYqKLwfDrLFFsFzEYuD1HTOOMgjoKtuNC9g6J8WcvttFobLb2skT6E3A9M6733Du4HLYkr
dRtXCCjxNPGEckOW3tI3589jY1Gr+qRM3EwoSs1mcn7lQi6bwp2cvn0hYv1scNunkQ/KbUQ3TI/U
lmlFlqjvicRzU2pgCcuq7vi2HNc727ZgT9lMkvoWiCuB+xlWcG3KdrwAgHhbhpUGfQQ+MrXjJPU4
UCxuZdeYH4f/fClbH49gfIBg0c2UMDWObbayniDibFbKM6JOdFQvycPlQBncNmjJ6aft3aIzqotd
XANwhP7S6An65oL3OzdNhi/i8D+yZHmKlH3ziAFW0Sg4ddlBLiPXPDeYr/i52T799rFCAGcuoBhD
8OwTRl16vI4UAyuCrJSJ8ZHnGKnRoP4TXTE8dvSyszpbf2rh8MM2SsAGEc8+6fr3hfEJhs2AuDND
8SZWNNhJhvzPWR4gdUQ20KVM6qaLirvKoVCJaXt8CoJLksezranMw9bnhK3joDe8vgSEfNhCddXL
mXgxJkwmuFPOI+J28vvE+LnKjPEmrM9s7l+Bn9Ly0+N9FBJ768uFQAmHWMj7NrOT6hZEB2V2CpqQ
IQDm/GzFF0tBXx6+lTxYJpH2PJ+IiuclHOZfUiCrJ4yLwIAO3gsr7KDiiFa/oG5MJaRK1qUZtyYq
CcqnpXxs0nyeC85MwUThrcE5RcJryYJyu8wlIiQm3eXhQ/RFHE/DScNSudKENTQzbHeh0ozhCGwX
pEZD4ZS+a6EfEe3843kIcE4ApqWjQitgILvqQT0mQhxCRzX+IMCnFMbHXjv7VkTcsZl4HMD5LYIs
EnrMhhGVUsJLY8iEbDHX5nWvAv5186Xrvq+MdW9qSaBb7WITAxuyXde7rauJ22MmVSaS1PS8g2zp
59zpohnkwiZStEEY6n/3SKhraq6OUG+UNkc+ZrTIvAjNQ36RKvQ3BLVsYxSfFIfZjYqyam7G9dRB
GLLp5Cz5Gyjn62qGtBPcLjgu1jwfTTPRW6s8Nhd244dY2IqSl1YEmpl8Q/EmyFPTVO/7zj3SOA/P
dhZPywe3CuInMPS77zJP6/kHbECBxqNMsSoODQ0JBubcgrqIgXTMqH3/W4ZwdaoDJRTuJ715cuIF
iUT6rrAmrhk2gcge5X8jyiATfzGsTE4HfDzS3xTqcikoXimjJ76lXYUEZWzSUaedsepO1nZYYYly
rcoYPPHP0hi57jap9QpTvic23i8iOECfsVehgIK7VQSFUSRjQjOvsbxxCC+Bi45PW2TI0LxP3Vf1
u7evbZQXqq+Lnzavo6eZ5HPJ8IcjGJTfpuwoDdL57+c6tmHmHOI86w5/UOiu50BntfDsJzRzPYaP
BNizrCiUFrz57mW+P9tytHswT6KANAILTK2fcsDA/vAAwvpTd6GNMKlo7UKpVYWFzLYoAhgxpX07
AEthH6wcaN9J8gBC4OBFUI2wXaNX/+8528y5B34Lo+uYD8HqoOH9TfBPqjRs+mlV3mqc3GTglxIi
ezCDfLPB6iIHsPgeXxmp4QUHrgz2OE19+aHuPXE48fzy7utNIqQPEyECKUgp2bY8LBDPzjER1oLL
CMQd04viJlFYnaiPSHVcZ1ejDcz2bAsdqoczn5ifpaJjiXvXGlN+HUl5ZWSq2/TopJu923Gq8pZo
jqXmSaRe6RDhDpw4/LCDXKNup3tATmwdV/aRYyemUhvpgfCFxQ/gC6UoGKa+SYbNqh+SdzewX1cI
meDPOV5zbBfDLsRIMzoMIdG10H7Efn+B+ZLA8S0L6WuwFk4k1ZUsnDtyFUAeFrc0CNuSNULgl+WI
dEWUq+W1zVXQQjhpFfTElP9BUCCcFgkPZ+7Rjzw2OLkrMFGcEHBN1QvUe5r9aWlgJElWMNyhhxPR
SYyafd/GlwxumI40vWSoIO4z3QVkKP9YgFqKQe0pjKZ+AXcUvJGqOgYcrwc0JasFeSbTl6QLXtx3
yObZsiyGkWlfAaPxnPjkGwW9SHLrHhWR7uD/90RmCDyootgY/eC5rVKgaN3TN0hstypXUOhxnNbQ
0WJOP8g3of7dnxoUTwuQTpojfgsGdV9cAW9uaLWNa/KjTheXUnU4fGUkkS+WFIGRgZG4nd1QF4HD
oAfI34ArL5k8Lbk4lPbfISYt+ncZ3v6f++6BbhtBv8G2Mi63IWsn56HkVo/vHnxR7G97CxNpCCdw
zPc1uOoIthfRtPv4PCPvluuTxtQFE50ua24bBbWtNesls05ZEvq3gMqNvc/uUrDxR6Y8YTKzKCvy
8KA4tg23abnnKVhQgMOKLhr5DpZNS6C4E1Gfzs2FW1Wcr3FkBiKrrJUe/COnpgyXlZlRc8wUWVSz
QxTkwO0gFY4iqevr9lyMzY3IYt4k4LDppSaC6rgV3cpvUbg87s8XQ7TrVVsZ++Mha78xvue/s/cp
jdPXdQy3uvT5X3Uvy2ahz6LxBwmLL5eYVeJvwLTXhgbcsADMA5r/FAS6qILkkqqHFfzXz1tz503L
LIMPsdgi77PfWujSrtlIj2AF6aqUwX94HrV9h3kif/82+sSDcRDvpQ0m9/uLnJ9MiWKXtikxZZ++
TxTiei3mWnvmP5GxQYouPM79Bbwz27HvY1WfMc0DxNu2FvLpgcdp6xHpiDsrHcbt/hcRfQHHOCDd
/nGg61wfN1iMeKnpOwtgKCEFYug00cne94hICtRCoV3eI7N+rmDBNXVaY2gfznQjO90rFrtnORaZ
P0Bv0RFCH9iinZdSLKbLpEhVhYxKw+w6+1x2l10/+fknwpi7pClmHD32MZsk9qmWFdPUpMt1g0xa
RjbFw9Qh9kLeJIOnQ4t2d60LtTU21A/KO6kriw3Z73TfCPlz5yuHOXs8aLd4RMQWi8SntqE6zKwa
2lYtTrwHNh/veD5mLURIuRJlHeK8gzGLRYV8TN89itVnl0+j83/bxOO3+oPUTNFw6e4z7DDgpQzF
/1sMSaPCi2mpD4s6B/hKuLv9sqL7YBa2CcOk0ITMJ42iBBT6JjCmcaGjYbtxSgun1ks/UPeyFFrN
fHWlss7rtLdKoOQaJ0+hAG2oVU+8DcQ0S/dBxaZjTDp2Uq1dygbdwb+x9ZXV7hOTmE0tBO4wqp4h
76MrtX78ahrbijfFp/kzt8cG1SwDc7x/ORePDrxwe/2nqxJNNtHdpFWUl9qAGypRWyUqc0BCeAzt
gs0+IwUSsEOJk0CdU9/S+d9edpwWQl5vJKwK/u3TULzxQsMcbhiFL3kSrjfBpUvaK/GR23AE8V9y
UtKrK9iUrEoBlZmwqwcwR2X5YAfy2Dr26V8ESvfCh4gYDMMU7S4MM87NqBNvOjJ4QAL1D/0jaNse
XxwOR2DDDRA5ceU7jTE4FM2pVp3i6czbkCQMFK2nWC7kws14z+xNyGtV0sTfIdMNqUG+iNxPWe6b
mB/p84OFgsANRynMg4F3/24VC67LcrnMsXlFDLAYwups128M/XoKvb/68AjDQfUjE2+VdWxLuPqn
5rMHQ2nddsKwaL8eg0rdicckRuuPABcSI0NlfpkRzMg+lEBNSsjXeeJRJQwg/5F2ff9hVx6a9FfY
yqHpgGXVWwlH1j52lwGQforCzh8d/zh0CNqxrVRPsWJqgOiEHv6ujdOrPbhYGchoeYN+qKaWJdks
g9PqB0Tz50cdiJRyEHofd1kzeMqNGHoiTVKcq4XslrWKYY05cn6876ai/b3a5OxXuIVjKOA7BIEz
OkpYVtHa7E1V4hQhJFqXUwOM4U1gyEDsgX+EnnJdfHF4cdQM5W28x9Mlia3IFcaLMAjiRjZYEbZl
J/GFJ07TqonlKS6PUoLq0l8h9/1XXoofG4KxucwKq7AW54g/PXCncGD+r9WfFIakxIPT6Hw7/e7j
AvW2PTO7SF2xGuI6euQLfz1dt0cQPv041BO+PnEIUwzPB0z13+4QI9bpeE+Tbn6KndMO0wgfYemJ
X1g4g3e56fEJnicCCejwY1h8QJ9fAPQYzhMvvFJ00cEk8dGg0B4bfDPEe+HilfJRKltQ7+9b2Xz8
3qS1nMiN8apbCgaaCoKhB/38lsmOPgsSQpnUPX7F2dK6Eak+eloAvuLdgeZrOKmZauj7xEB7797m
b3c48aGzy99/Nz+h3+To+T4cMpgiDnqQK8MFDF6seVKl82IoLIWbnVlWJvCPtTz/ZtL+Wj2/FDnb
mpKRbCM9+abRBpA/pXwarPLszhKmYjQKC0NRG+tyv8R9sGRHjtKQzZ9L7lv99lo/wIoSJBb31ts+
dseEcSgDHGCEXAVL7O3uwUgJktDnIeRO3TXRNlb+ThccAZn0/YQHy7U+v23fHvKrn+wXMQuBzTEd
jV3YE4wdX3R3A09reUPjsN/SQE6Z104VxnsnbdbS+4N71Jw4rL+dirrGda52FvJ4HKPelCFzsXvS
7zPQLV3E08vuEie/wGi1SBXXeWxjNaPS/m9ErRxHPipq82nodhYfQYdbk0cn4gkibJN+1gtMGcD5
ox6UQ3yPnDd2saNX05l3cVlL7HXbrUciTOYLxNPQGTb/K+EDVvKNO/54QF9GgeimVHHUCTn3jxqs
aaU350HSuw/08MUQ5ArorY6J2do66u3zOFFwwZHMv+xypPaHZ8vwvr1LPFSheRwUluI0lu7wiUxj
zPduZxITFRnPIgxinruC4YS14rFAdUVZZMWm3IEWQhA9xyHLV3ALY/kMYMnJLWmyczaqqONeYIHf
WT9pUSAR1jXPGMKMW4I4sN2LfVeMvy02c4tWUXP+GyWxy/M9f/o2Lok5qi4cTYvqczXTPeAkbUh9
R9fJc7ARxmQjYM6e48sBZps0v1exJ/pVl40PwTQ7Baj5STCAd3cT5pHgUpuljdGhaUIJcxjANmNQ
FnEM3zyCBPgEuCvxRAI0BwJuCXKRBsGdSYWlUBW701csjOCGtv6edKInP8D5rHS1YYCmUQz0qEjw
U9tNzMkcbToK7pVQOY3kn+HHQCov4AovqJHaQNmeOKg1tn3vS7stY22xNQDeD+YVaXbz6KD5XYbp
p9F6bpAbJqNBX9BUH9qUBiFItNHGkfx55TlSfTaixNNRPxgR4n1MN6ivZXjfEkTZTwShtaq6czpJ
Q/mdvaCZKnO7Msc76Bfx9BYqTLdUMQw9XT1wpdI+7+jDv0eceWkgOIivXp3vZY8EdBsQL63v2QIr
6QHYKs7188atkeg+7+MRXRPsKlsvyD6hDuCNua/yGbr/pDo2V0OqjCXrTxMenPMNBBmSfuVF0Qzi
OA+BXIA5zwMgH4Izo/hxIbhd7T7FJKPbsEfdCz6fa7uMzKzF1//5aUlatWLsAT4SqTplY+AcH7zx
SYLr+1mlbPeWaE7FoWZS6DumlT8Inp+pI708b9ub61qO5HZqZen4QVXHMMAWFbXJA4wQsOnFf/w9
SW2IpzOIwsJ2+rkR7U1vcaEhcD2CPT1GhACNcubn5OIW8SQ4RxYsY31sT7Bv+zWAXs9cWTwDr8ur
l2PBzNLcXTRwg7ngq+KmqFfIPQGhG1ow510bGiyDl6NPw7wOic4x5K2ALx3c5P5EZlUG9L/HVtZe
wpS4O899TY7wCk4fw+RDg/InFc+qpdPEqa/Z5dsvsL9GM/XJsRQifK9lW8P+jzSOy3ogFMjK1Qxu
G7iXKIwbqxYAECzBPGA2Q9tgjmopnqzSgskHzl632FtGnS8NWZOjNvPTqw5JSDLLrBhP7ge7K+r0
a6VJGSJzWIZe3L5TTVlnQU+hTWK4FWdVjwVFcJR3C07ozhrekJwMca5xzWy/VZBQfAFgq0H3H+Lv
i+8XebeI6nqyLqF21SXx+yMILcqZs9+5Q7ZKcUrwnArOsYgmhVCqB0r9EhC0uf2OaU6BghhzKD4N
UgUNEawSWIoNq91AASXmcm8aF0pPs+oVLhdyMmlaR2+jsnbbne0SzbxNAk8c+mcRepm3U9ujNOc+
m9PcakXsDY2VEhB6brs5FztpWGSUJQdwNRuNpB+y8uvW0LTTASTDIOw3jsny3rEPSW1uzCV+ZQbN
iERrBprapHh04ORkoqRw5a3Gnd8o2b96kRubreStONott6+FVgoqUy9cK576NiMBhCgNBxRIap9/
O+FBhjpFK4qVZNVc2Fexw3VB9RATsFjtLcETWN5Ne9LDQKj22jvhu0RMENH0HO/nMAJIPu5DJ2DL
zCOwltxPQ4vI7c1iyhIQufN0ySG93SFLcSQhTDGq1p0rzJB8KqYBM/UUdMOwgm4hfmrX2S1StsTp
wdXVV4pw73Cw0jUaiAFVf2DvJrCPfPFHThnowXbdk786OfNkXUU4MApxDn0JE0Kzjeej6/MTBdZs
vMdrs6UWGxA74vam0xKUP6QoYJCpbDBQo60HB6Kbz1NS3jaLLLM6OhUDtvZNca0guy8FcWBpykiv
Yf/GLwWaIPknS1aDFEGNk9MlFheGOgZmPMFRO3iPubpO8Q/aWpTSWh/KFmIjYkCQcjZ8Gud9EQ2s
GTl9QHdVJML8+waRQBqiMq9nKUvsVvxU/rPyWNNYh5KKzNfJ/X/bkb8vVgR9AVh20FZUp7QpWccG
AHwdZvo+ju0cDA8vxe1HpPCNNr4de2sA/mDMPXZMmEDcIuFJr/QjksqEdkRTMUCpvAjGneedQ1q4
l7ichrowQS9jx93CtX5/t43LVrrPlN9ESeCFMDf0IE8lHIlHqiZJTOY9m3jb45qANdkEfC2ITF18
rbxwtiK27WySTADQxyYWuU8LniT/9XrgL5b838KVqiCpfpz/TZUl/lObgT2vgl4JEjq1SiWNbAsT
/wF/2GiwfFAcUjefg6Im9WpKwFMvhYEN/YoTgoAiRB4l0xjmmbSeYkOb6H0HCxPAAO/aLdhBpu7m
QQj6j84OfnI/scFghEPhMsFeApc7AUo5oBJWTUwX4p1obnwVsM4K1IH07FntDedPfRw4tgKoQ0bZ
sL2TL0qIP5QQ++/RETJzENqINtprLOn8ny4Sq8Tib4Vr7RUt+bTWyGvMDFVuatQC+b0fmJ1UCc98
gkp8EWBQvVhXmKwP0/W1DGLdbecP09reB3IULLN9UPyH6VDZxNe5sgrIeyLMJ+403AXDbDTTCdN8
OSKrKv8e9pzpWJiXYHWDdb1ZGG7GyAJGo7+dcxaxO6MuynV2lizMnGshogLpRcW8Kcyl6QJKQU1b
Qe//sAddkm+ZQBKi9YthmIyX8xtusJytSxWR/tge/ftgHfKlYpuJmyFIyUe+gSMP8yjuttSiR5OJ
Glf6rIVN/1lh9QS4SKjW63SiRhTEuBd52+NYTIAMNINLCCe49/FetVH5OBqjtSO9z2R9+PAFZY04
EHEjX/d8Otu0GcM0iR/VL7xIgtTol8taPq8l9azZ0rQuix7RY5kNVlfueGxB/2veoSYbdtQnZsga
aryIpibN66Ez0nUj6HriVQHiUhH1XW0nkHwj7Rkzp3riUEu7vl/KwI2YMZH2mb9qe5wmRmZ8Pg4J
3jQnhTz+c5ZkpK0alYnnScmAX0XSos1Khvw6pAXBLx1uRHsWIABW9ZqIrayCk4ReEKisnAgduigC
a0w06p1ISxSGuojtsHcnj/0d3PW7Jy4PQ/5LLxlAAhVjjaQZ/pPg76QswT2LCK+ej1FjYm6o2D9t
5uQV/yG/hd8dSKE6NoftekdfKIieLfhtdFJw02CP7HiL5GXosJjxBRikYUO46CMVglyBiJxYpW11
6xC/vtH3hdvEnGPXmXyQo4Hw0NuEit8pL6LBYwAdhVdKxl8BSPPOo9wWYqGvkuAsDs5ZYqmdJ7PY
37S1riSdrP8csxAySFrwwSdQpCEv5+iLvS6IIkVXA4OpCsa/ITjWj5S3QsvTs99d5QxVgfp725UR
09H8TBYvP2HAqz7Ar96yUGkc4Svru4U4Kcl2FytnCbv9T6Qq9nyek39oEsGz1NjfAH2a5m/qyZ0F
wPYB3Z3rhN5P2Q9bbWoTjZxipeMUyiBlHB/VRGYS+fpgXtmZ/QAkBai6Gvc/712u3n8hX0VQK2BA
FuS1lZ+qlLbrqo8UKTxG4E21LbueYvZsOOePKckDE+Fc1+2epp28N5boKVliSv7BSpXyP0nJpp6B
ATmt9Yo1bv8Iu0TUgxdpixbJ2W1oCUtmD65cyK98/qhssYCNlV0FFnRjc4im1Z5CNjqsSUsJZZrM
mtBs1vON4yw1Gc6m/TZFF19vjl3wIF6fDZbliBxTbhy276CNgMOuFXAS4U35pPucrmnFctPm7xF3
iStl9F+SJMvTo72AXTTzW5M784YRm3+BaRTecuWw3YMI57VwqcKNXLwfdNrAPVnW/ltQhA+YhVSV
0uQuvxS+hjReX0uIwZWdv1tuzFERCUihCHm2HQ0Iulo4BTBRvaYpOpz3x3NQzanVhQaHQOzz2/Vl
Bag+/lPQYmRA5lr5MpAgcL8ZxGIKA89uayXyvzv91tRKdeJplxqvlLv6g4rqVpHB3A2SgcHQ0fQ4
1+Ow1elJY9+ilihylEVnsDjDyO6AxBXDZiemdUDf5KuEOjmtz+AiSRWUQs+adLpdg0EWVJoBLjRx
zIzbJt6QULBzWkUEDJ4BHAWZH6FGJl862EFeiM20thCHytzPQCpJ6ZLvvqTuNeXuuvmjx+/dU1vg
PX3pT5gNKcLJlZvbmYQA0nub9J2hWeRIc6zTq+RtBE2faUqnfTzt7LIjDC8+4Oct4w3R2OCNr5M+
8fF6wW6FLyGeHVVgqGqw/IIJ2DEix31zBcmrJ2Dm3Ww+wDX9QDQ/Oer79Nf/hRNeNfWsL6qvvKm/
zncvanUsfIrwvtn7Y4FG1XzKWS9HTJ3FkGopWl93XaLnGuy9zWMzHAkI8ZBsA8TXhzutMqrhNY4F
DboY5Zmmnnh2J0FEMbEiLUGeocvqqkig/V33M4oZPJ4YySdJOZBAU67Sd7Bcaz1jVTGoPb73ulB/
9uos+fG3keSpPWrMPUanYUd/vNBOLd4r5kaHTDVB0GRE6uf6q/52laSl+oQt3/8OSSUd9EWr9ZB0
tzf0o8HgTjTx64Bs3/YmqOzMUL5jH+Ik6qYsxrNL42oYhVlwEAacY7UQymuvQg8BcY/eOBpQH+4A
53XTzbupcOg9tdbIe1kdgtKEEdweh0FODhyr9DBGlvbRVyAtfRAU1VRdCJhSc16fMxeJBgoDt70w
tAyR2GH44dYy1JZtLho84NPKad3+5ZwvAru1YtyUUs96ZMnuENV23/3Llp9iKQQDaVGpvMtVZ2Xv
Qs9j0NU0QgzWO9/U8moYb9nds3hCllUEX51W+789BfKboqk1/h6D/NjxK+aQtAggFRPjNiy2hc3A
eqNyJe9NEhZtnLOu3ubQIgXoeybnbToftKoZfZYo+4+UEzbMyBYVrb98r5uvzuiA7YIvjs58fgcN
rspCqDgJhSR01nbBj/qGRJW00+9gecePjtTAkyh6i3kRrlCLi3+++40M2RwkbmFWKnyBq68CKtgt
4ZFp7QcKReIOS4MAxZKtx26m4IBDo2nFfbqhqXy/l9+YuEMbBxBQjgBFR7BT5T6A66jg1YdIZqBX
PXFEE5HtsGQ8CkfWVU/uTbMIbbzeK0g3zbDWq/Ps9T0CR6INbgL1rD9YJ+x3wE718sIPx0yYCfKT
7SdwjoEKWf1bOWB4sdTh2LY/UG8dcHgx27U56p9eRaonn7M1EXNLHM0BZTLsUsSVD1s7jVXMzF/u
K7XkQ0atiGwt/bioRWCtIRHah0kRNI5Q0UhadTt3JSRQcnv1L9qgnIAwJtuYKLa/MzUnQXzq3Rbv
cY+Y4z80bUODA54ZQW9dgygvlJVZSzlsEXzvSoltAnhMGyNpcmS2fTXRwaIzlsPpfut8ZV66X1i7
fyO6fCoS9eVDRFrjKQEi/97FcNzXdZ/Pxj3zu3Mr/ijy4BnW7kRS/z30ZvDFB/YvvSXG8H719iHy
p80awlOI7kEg+wnbjNfBqEqPTgLa142tARZRQYHCpc5EgCVHVzhsc24Xgrpgj4jJSnGRUvvf1GS2
zxqvTcKlQgDPwoBaq0MdyxupP/7mG6rDkx+Zd5m0QRoQvvLXJqZVgxNTekTqHzQSZyFBIW9sBLfl
5lIJzxrpI3QX+27fPZUbyphcdgGwNVYEhkuaAJe/RmnjzEfwgQmU5siDAGSedHvexJquflGxJeaH
MBeD67o4Br4kBITH7g3RvBzWjSFI0v9zi3d9yec3oGqY6Q0bvNtYNVqR19nYztZjjbbR01ELfSV1
iBVgILeBJC8Ovtx+W/niM5ZdLh4dWnZO0fE7Y3WI4Lv+w2r1pWJdkji7NTyRp5yhLAvNDcWbVxcp
dH7Oi6dnj6s3SDbtoPpTWAFC+WUYJwBhykMbUBOIJTLKRmFMKqJci7M+0LZWTY9QQ8C7/R/NoBns
kuuXwo53WSasrm5DkZ9g6VhBFhcPWXTcOl2c7wezaX0cUn2XIIi8nxfPFQNICXL6e+jh1iN3dehF
1CP+raWwZ59Bi+cj9/BEVtw2kx6NBJO/Gpjwx6NU/Qm5yH86Ab0/RDD2vyimAQhEQmCeRNJuj2f2
7jj1wRTBGTZHWhr12xL2monwzdbrdGxKcHy/fXbVDEQdhrSB/ZGYbHT6S5LNQrld8dEaHiPNKiGr
dYngj9LooyrEYPSpw/TPak7E8wHX6byZxrE4R567QjNaQrGJNx53xiDO97c7uEH2SbjPO2MVNYeS
oZOEjPkNu0fahUEjWPm88+SPjdqe4+V722VHsEjIOxyWlIQzA7OMVbx/UrPMUxPtwpvBT5qaj3fr
YzaBHmWxGw8L70xm3sYCSZ7sDuTkmMjRE9vRYkVLULzU5BPOInljWWvxe3kMTfKHSeE3fhJvmQYR
Su4XtHGpU/JiBplzrMbzPU8JC5oGksZa+a2reMiSvZuMF3zZ/T/D+eXILf0JYbcE+zhP5zqv+7Dn
ZntTBwS4oD61w9+5zWdiYQdQbsUJjzKcnsisLeFgbeSdjH8jZ9GC/VmAsdLbhiSnU/nNdEAN5lSI
aWI8dB0HMDAH3/BmCxUusyxU/heJh64RP09dZzpWQ+fV4iTCpTHfxmGekmhFX5ZArk9gO5aFLd7D
5Ccjtc4wQ/MX03nRL1B+I7JAVadrd9G29r0tAljDMliQTfC4PjRMHS5DU9KjesixiNgG4v9WFUue
E92q9DBFV1FIWrmaDw9I441OsRIfgb6ehUOxHF12yPQ4IAYQQmipuAJrSFfQO4cYcxpqpLB0lP2q
SbfHyR0ECC479t11Zodn3O4ZkH3QEN1eXFENTRxy5+Q7VPy/EFGvziqdyQ8i1awjqLqWpXsAnuPp
XKY5xbfsV8W8Y4GOPxWCqj/mIfuiLi7a/zjhJ2cqzif/YMTAc3fWO0iq28ZmF9gG36Y+Vc6Y/tsW
uE0npxdGw9MnIjv1FfMYMKh2mHsC7Ul3hs0thx5TgaCU27/FWraRNl504JcUxhO3i2XsGQzjLoSb
/Xf+ke33rlei9n4SKhaLt1rpBPeFa1LdQKwaTklyNNfVjkqN2Kt1Ivx/jBCLEsaMXhbhZg5Z7Hnq
UQvZmpHEde+USLv+cNdSzg2Fk+SjYYT+C1owOUj5VjgJasFUkuaN6zU=
`protect end_protected

