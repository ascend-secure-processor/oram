

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OyhpSwV8mnf7rurGFqgbHmhCproJehha5LkqdkYJOPk/qs4zuo2D37IHzW0AL52NINiRTGMs+1sY
7IlJeTjuOA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o7EmNjHUAh8yCt07byLodQMevFkqQEvQX0lRiND2Au4j4tzeHRpxCWBJGrPYvu7aoC+2jwByo2lm
JwJHOKG1N4fOUDK9cZD/7eqlgQx7aNQjZj4vXIqjKAq29Dawz6srru1jwtZU///aXB0UZvRYHSnN
DGuPt65b275Hz+L1sy0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
w09dCKMd5cZk9y9xWhos573Bul+P0/DbboXovqwpyATTzMasgkXBqAHX3jEGXtQmJz1/4f6IkRHF
bMgd+EU7QVHfisrj6ccelt+O7ihQAcqFqG8tmFV+nyv9kRXnHKCPUvu4M2ZYEGcuioA+gsVSo2SF
VorU9uDCutVvLxaR9FSDUHquOgpd18Z3wByjRNG/RXgho1kDB2lNCWeAmRmIGFLbTwGQ/1CPxdbw
fzgsNESHh2x4gjDISwCophynjo2hQeJejd4AY4zEl6qJjjXJaAw4nuPOe3Rns5pHf4qFtcibj4ZO
pQ+KVB9RzsWSNg0lDahy7nrv000MDPlN/zI8Qg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LOrnkqtL7UXfeWA0GedMarggVdzTLYA8EW/EOLwMazRMz/8wC0diegP0ERicUUOv/wpADpE81rrb
Nomjy5BqYGDaETYXIYIJ84Ke2O4VMRTAEkiDONHY+/0ZAibbVTRA5zFLO4v1yPHbhPRrkLOrBtZk
Pzu2NXwfd+VA5pGKkwo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AOnfFabqcs0c+tG9dF35bmVJzDUX0Zs+3PVcMZhdOF/zhgOX0FR0RjG110AKdwKVsbgMWyUKb7pu
+bcRLioWp3YOkE8ImOMGMFmSlbgSHqZj1qMtd27zgyFpUdmN6xiaiN2PjsYdXYAQheRjjTxuill+
R1JSbNF5rWf43ROHwVuAUblNclvHxY7xPhHCgIqRe4KxfbsNdkWpYVNW/O/C87J3PDLawu1MN7KQ
skit9ZJDNoxw8qhTntUHvigYBgWAd4zwUPz4aENJ1xIf+kf8NtjFBf8xD0C3dNpZkPk49eyabkiq
bin5DeDQK2c9gONEoED6rLxAQ4f/NCCReRdosg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5504)
`protect data_block
N+1uBZ5SL+n6skklCQ1FD7Ne5Th0GjC/YhwP/ImcLv9ZwW4jlnqe7MvAqjm7AGmZMx7ifpSohM1F
FfZcR45iaRkzw++4xmvhKhw4JyMywOdyCcruRmAKeLHn2u3EZgMPcua13xPERV9b5p+Np0l5paku
WxSSxYmIT4xMIWHPPlOdVfaJLax0P+3+Qu+lQ3WL8hR3rSYv4VLCkIb8simHzNFhvzmHC7Y3DFiv
QkbmzMhUvcaN8rMIu6o3R3grWREfHKP1gtynHXspVEFqueg/4N6uBO9Gf38JkjYzIu0akO0PkGHG
YudU0n5haCCz9KnPxJZBnFLrP3teDZ+9CtoQPqPUTDaGRPwJkQ+L3/2ZJiGgjn2Ay4Dz7amSSs7g
NuVID4a8PHLBBL2JAClEfgWPzIteRwPlLEcfJMa4cVul/pzcF2UGpC9oNRHJ3vCJovkWIeU6pjFc
RfpqRMiVAhtDaRSq6arSI3wxwOflHMLEDDoh//6otQpQVV5NztqgqlyZ1zScDvXF7E0zeJ1dNMrg
fW4JEu8xNZs1kNsH7auyw7gtV9m9PSBE5GW2dj5JVihuBgn1YgjFRFFIvQABYgOAq30ZORTFlslj
b9Av8PfbOalCJhEhghigb+aNvue9sypJ0/DjoAGFLDjZroHrzIQTrWeQ54XVaDLxqgvHSeOG8WuH
wz4yjFric8QG0MYhEpw9EerztvDSkRqJX89zXiHPDBhI+od2gZXxsaMCLtj8ndi/2BGIZ8iBldhl
8kIMqtdkNmbCKKnaUoT8tvttsnhrD7nRURmTcgBfjTv9M3iRYoktyzw7MKSmwQGdxh2yArpOHrnp
OsHvyTpJWXdQh9F9I1cPepFLh1UbhT9Q1AwjOPxdb6vue77Tm5RRsv01Y9HR+qW/lR3/f2aOf0Bi
oSP+mNJnwfvgeSiJRbcRquWKtDYYNy3GJaqH3HUkbhXE6beVR4TRLyrd3WFc6Z02WhGg3vRJXSSb
sRcwFqy9mYESAFfWP39nIScPP2ky+WxiMKP3XANYaGzvdtBtSm7JuYz7rO5AeIyPs/6IvEFhxJ3+
Ur0Usm78PywoZ4xzDq7cXbXvpDwZ4LA42C3hV9Pjop2iqetS0GFd2xAf21t26DNVRaT8tqt9Mp1Y
2oXIzRNR7kwzHEQA98rZwETyVrE6jPy7A11fLPkoEs6sIf5SLOun54p+uWrl3ydPLnLW+Yy9bHmo
gHsEmy0OBMKmxXYDXgybIqyMWoNI49aVZ9L+e5dtrD3aIWv4HPiqRr4Ka55cMAl/wOD8OAzC64L+
TxA4vMzR8NeKaVFu8AQQowJWVbcVoT6W7enjv51yKDHd1KfqbtlZcWNvGLVQwqAHOBWqQNt7guB9
t7tsjMoq/zysjqnmGs5TC1BvPDd+8clljQzVq92f/jH9njC3ByA5ELzFHtHf7wzjyemVPA56Zk9I
vwkOLtEA+ZVPsIKPP9MHkoXqiNwKwjbxc2AMWm/+HG0DyymY70YVGv3w9nDVY5GAfjJbrUW8Yzxs
Gi0yd+x8wZRHixp2hVDCFr+b3pYpxNzYm31OxWVBO8XHEFgwoyc0HiBNBT1sZxPj2SYVNSCFkr+F
gNGoigISpwMPXi2d9H7DXB5AhOx+N5Xt52ftkm6b/ZzSVnSqKskSp5l1ZYCDpNk54WbXlbjJXKuI
cIXmIwOujtYDwoit+seUPO9kzxWWKv+4qwABGnpWp5GwgeR/nnMTDBdHtNgIrlPEQhhs69dZVTyU
CjyksxXQbDqu+1bbSubIefqiUBQkTm8mLMamsWvkNgKl6xk2HY6ZbetWsN3YVZmuf0gG+lSDnIRu
/MTtJRNSJYpQT5RcvyItjWDd6voo7QKuN5bb7vxNcqkyEzDi1dRdJ1JQxbTKvJJRNUPfQvZaWhVR
GgXlZf07n1xdUBol1qZZcAL64uMSD/mqghjBu9V/KgHY45Kr1jxAtm72AwpLeTFM+ifoxOByVgs6
fWRtMa5J0mTbqvIddzKaN9/8L+H0e9RVZGVKCjp0ZnO68voVWYYsvNTUnHweDLrwgWiqKmHFRcdz
TWW3QbkEnBsiydtRD+9mju277GJ4Z+uh+GOzmWSCuOGZkoSoqjXVayNfam7y3qU50vKi5ymxoq1k
2gKesysQrDMG47bkbEDv+FbkB8nqgKVus73HRTs1i2EhZPV5bwzIj7DtEWFGz6LoglMl72WpWsQe
vBCf+qUv5eYUXI3S3OHXEwWlbM82HYEUiKr3rux9Mx3eh2k28xDlRWjz1zn3LiysaNevlGu8Ydlu
Cvplr8olvXuYra34sDxkiVfZxFsk0PVVRW74LtOt78RnY9tTO6d12pW0BwzsWJwVpzh9iXI6Ajt+
989+vBro25Oy43NO8S/IDQn7PKW9FvDPpSaYxgSFjxIfCWs/wVSIJef8APv9Mj2q2f9XEMJiWjUf
qfwyL6kVOfuAKp2nhVx8HfhuB2+XJwHqSvEWquo6rpbHtqekMnlpni5DLDmoLi5zGlxITbQD9D4i
sK9N8kjKvw1uOPnFCqDTUv+MWbaJo2MvhESR7nm+1CP1Kaj7mo0g/ouSMXixN2NwGSKTgPtB+avv
M3Pkt6CPxxuXEh54lndSnCCuo2dqXQEvVhhImbmuV5Ncbd0unOVWRli67wsHhy5XuveNzE/YkP+B
3MGaoxenUS1/2ZwuUZvKYuchcHO3xwzHtzgjTKlnM4FFv5gKCACMoACySFrkaNt5GzpoJPJZFCvC
hUYbdgDlokUX+eyG1fEzDnlDuYjNkylthJWgJRR9EQ147Pf1iNYBTWHAEJQi/HEqmG5ucJA2MTeM
aTZWGGV5vI/w1qp3LLGXoUfKNXEsuq3aKOwcFjXty/gElCpdTBCQtwS6wtvWIwlgoUbY1TyaVE1F
ltU1nqVa5HR57yN5NuZZy7ZzVWnimj5FXWuV79+vohfglZid1ASDQSi5TGTn2mmV44P9VajDREQ8
7HYHgKkxmzBAa23JJNVMf/g9jaDjqN/SVAWOuTMwHuJx5SrzVCfb8cMb181m4nvf+3ngyPc1bg1g
Y3XtUR/0ApMhPxgYhme9wGsgtzKZlvJ9Rau8SxsM8i6PqTORfReJ3o7/nyiQZMhFhrofDdouzBWU
384imKz82oQOy+E0Me0CzXvusAFInnmrMDYnFrqHtzxsYon51LU7trxK1J7iGnrymUEwfu264BFU
MpnPE0uVj5GtsF10+RWTnYkYhvNtFfkh3ur8olBz+nj7o0g1G82ouRRFZPIe6iLWci9XZtfO9r6o
TE55EQAht2EEcS+5dncAMrXwQUN200KrwiXHWbuoFqD0bJjBPBhUokReCICC0xmBx8O0+8ILXKGr
BtXSaSuUx5zeqM9EDhitE6ykmUfYv7Cx0wazSpGofAeJTY/ep4AOPvBajDY+Qv6GUW86zV9gCUvK
wNhKku5Jq8lChqT+3fDwBpbNoGS6a1eiHOymrLDa0UBaAwcID6WdDIHtkgTZ8M2pcr+Hop6d967+
K4QbwYMeGBATh1ijkO97A1JmM2+Bg2Sl5WTEbFNlgq/y/GV0oCOSu7a50G6mtX7gqUV+4a3NxsVT
oDmofmd+yonovUhuh/bELgGxa7wSXkrVZgXVSEPJUy/EMnDZ41PowknoCNO8P6bSrijIUGKoFNh3
pJc+2zAWB6tQCjILBV4QqHrcD9dIGv8xMb+F5NyOiZdbcxDY6qdJKVaawJF26dPH4sfeShAZGFNO
Sjsm8N7H43uLGq0gbnYmiVqw9hFo9viO++n8MutHvGEutCzuoRjwWCRK6guGVvTPF7wRDyJekOt5
TEg1iU7vcDeKMkx20JxVsq5Y2WgzdRzO65f3iAtpX3c/BfuYizYWobvxotqnX03yCUWsL0dr1XEV
x+XOLN4ekidqxsKuURSEV7AEnoY2wv/AYi6c9I4qKNUVDgfrJJucpTJYAfm3KxDwfRwM88El0Y+4
Z5d5mFICPcsC0BsNU4t+/dBpLUPpsCLvKR1gAqUC+aTpLGv3Ap+TYYf1OLNHIn2+lR6i/lDWpcvM
MUSzP47EcHoB1LyKn7468VWqrSdI95gVydZlRwiR97ARzPaqzfQqEyhbaH4pphwgyRkbpSaFQHSa
3VsjZ916UNw/O91nyf984m2PihrAJarl7XMmXy5ExGtL/G4WC6cYcFFxTbkkmmeW4pqH27jr6dtn
RBoHEDBXsZURd8L6FLXJPcu8/2nSm2Z/b6KNDugY3ENwhZLq7UooG7A0TcXFVYFDZKeDh9x0TKXX
A2xphX+L75h3EwF59C5Agp+OiiOXIHxvRWj4sjkMaDPgBFQAb0SnimHstlhgR+mIXxO2Gi2WZ2i2
9RbdJT/G39FyKlD9udSixDSCAijH5hrXLRqLnin//aLiaWZiNnUHZVv3uXHCfsN6oRUIr9V0AYH8
APwHeGu3GhaX5Id3xEUnC9o5NxeTavmWbbnI3h4hQqHVhUmo3Q/u++4Q2nJZlfamPuEgUIZemHSg
I93ByyOIUXt/KUV9SUJhdvKh/gUPeXhPzcMo4Xo5tiUXPt5iQ4cqKw4dFoxbJjUGsMdIwHJxIBU4
mWLeIf2PnhaLH/O0BN0BVvFuvK1Fz1IyUlhA8BJQDKEjCFJs0UJRnQSmjcKVoqRz6RfJIGA4hDMq
bSn0oM2IDyGQJysovi22K72VKj+9bCGTgAIag2w4k0h7L/5l9bN/y+jORcVq+bsQoz6JwqEbR9Qd
vlTvYlBFiazODtQ06N5shhFxDk4OVPHZ2hfsG86KlVwdmNC5en8rEBRU6idBszaRi61hP9QQJIV6
WykPIX97mpGjCnVoG1NisB6dthSABjUHIG1X2j4bqFrr9eLH3FtdvL05LLtZMu9y/PtNDvP7EfLF
hK1x/qSYK4zyAZbXV+dm5agrBWq+63GueCaJTasJD6A0M4qe3YQ0mkxV5aF0qkJALuhxmE5HSnad
xXNZ7A8wnFt7EyVGmaAFuEAXTFoL14psjTgRgLCGTenc0LsoH7vMCGIwCZdKxC9GoBKIRMdsx1nL
0ZQAqcruzfA7QS3ddvLQzrL14CjqyOtme3xRot4AlT2DNVbsAAr4p2456xBP0P3yKS3eJGxlZPEu
ZqXQSle+LptoXHvKg5z348pW5MOtc2ljvijpNE5B+lA5Jvd6+Enudo5oXJcLX5Hj9AS4VgLdRrFU
W2kk+xuS4lVRGGbUc9/fsKeokOljVN+SMWUZD7OmhmHtfI7+MDHVNK3Rt8sJB6iO35aqlril0qvr
bZsCihoIpTi1N0yhmY4lg1WRa/tMdnNOWB1eE8w223Ez9UJO10bFXBvvXCL5xedBehW5XZ3WOUJH
HE/OLtI8CnK7CGz3PjbLrvFQpUKyJFtsmLRo+7wl8ZLc7Jhgm+FS+CmlWF3KjYgnfp2WH6FxF6s0
ucy7IsRt/5SE1EgHvZ6mvsjx2/dwLlJz7nqyr//JyVWn9LzkHYpaDB6VP6JTiR+vAqGzut2eoMHE
an+NbCFdVkUVIzNGXBAGf728sktp9rIc9od0ZgxHlNrPuCwWlgZ6BlXeeQr2ifjHAQwDdcgtHF02
+fLRx8LhJHis3mm1MLi3k9Zi5M3HylEPPgoqepQUqG7+QmXU8T0cdiSW6aHSJe7j6K+/kelF28Zw
xd9oZhc6ckOEC9T0fE/dfAAFqy2ihpbrItVy8dcgnmjMWT94/HzpBjfFBx+irfvP8avt67xqlzZk
cXMOxaQzFe3k1hWYsxv3RkYwh24wZOrII0+B8e8Fi0W4eDhuUt0zWAlKgnbGHCrPVhfqI1Ji3Zop
m9VtgYBrZQD03Y7vxFa8N1bdBxIxjNOUTvOz5PS7JuC2v7q0ZuCJm1+TDUt7LP9nDfdrupdti60Y
0Dqtik8eEy3VzCfho7ahXNj6/StipTp85futyCRV5L7nuzOx7HsIUQ189AOOVx/Cs7V/fWfjfai2
BYsrdsecfQcPXYhltRJd/QQ2bt75jkT6tzdwg9yOtQr9/1llES8KrP8vSaebFnjbdpf5VqCSgchZ
9AXsV9BYMLJZLdtp+oiRrgw8mRKUXWGIpoM+tXS6jXyTTcUNZTsMtCiGJ984WLVNRaFCmUUsxe9J
gbKFf/GOf1tKQ6yy479Hj6cqpglN1t30/OBd8gLmuLTFlz6/IliEgZdCm6keS75joLDQGXLVfgWK
EhXChlUaV8qkx7lgivZx2WLcXxxRSGQajJB02rhuMP7NIeTOXj0erYBg9LjJD8ETT/dOe7+M0m+/
qAz40gWv+xjhXNSMds5/Q14Vh/Te56SJ6cyQUeWwLL1hRFtuJTgwUWLiCzBiFmQB5Fw0t8dHOq2n
ZgRHp3MSciCQx63IVupnL8X0xUS8C9jS8W+ZtrMhHOw2RnumVKdQK0ytim3QKo504uh1zy/9TEUy
S2HJdldBEUrlcJuPkX686c/U/RMSklM4h57E+aWcJKHWmbLpm5OpabBvhQ8/isU6D33EAWnfFRxJ
8cG3nbQ/xwxhGQ8TACxJLoa5WmHaFWlCCVijTmMdJgRBaluqURMOBeOqwQ3FAx+Q6F9cp3QL/aB4
H+nEsq3Qos1hCTPWd8W8Nt2ktmXYxxhNkWBgcvqMVDXaWsqATvBnvK3Pd1kz7PUmpL/HgWyqrQu3
ExtNOncKSX0o8NMqK904QwBW7k3RzcFaktIPaSRlQSQYYs293XUIOVxSd3mc4mAUITSnUIyL0xEU
Yx2UY5DWwxZNRNOm6v21HTBmvRJKiv0wIW19Zj+RfIlLY35L0F2mrw27nlRr4WwPPx57GtKLtpng
jneDk8q6gG0FGGpBEv1M/9uL7/1ZVDjZCSszFsuMeQ137/sQttsdnd3WmwPPECv8KGSKfk8L5Ayv
RahF3xvSdKkQ3/L7Q8rnNH6xLc9xkk6LQ6nNc2zuSt4E+c2Uc1YTnSQE+e7JCwp1Gd90AhtpAyPp
0l2qZi7B8kdJrE6f1oKGO6aTIkL2A8+YJG7v1VxyQEfTmaJVAOI2GRQTLtVEWYFE6GHm75iszuwn
7LKu7XDZqHmvtefBOBlq30y2X+ZgXajRbXQGRCDpcLa2dSlWTz7phpXFIvakpux+/iwNB1RCkKz4
hn0ZBuYdglP+CA4NCG/4mbGigQN4XRqmR6ekxq4TZd20uRk3diAekiftmQ1gd9rnmCYmDCRV9c+2
DqQesWT16p8k48HmSniIoLpfWOiYnpZJM2RI9eCJMG1BNKFgq2DBjkyilKKp8YfSbgMnc6R2O7C0
hTYvyB4sn37wweu2fpj2cNkkCFtUsFep3lMNNWrYP0c8y5Rp95FMxfI1QnUuAoLb9iwJZ1b1abhB
4IokmeVfJS6MmHNgdJi3ep79an2yfOByN8omyjxtXME=
`protect end_protected

