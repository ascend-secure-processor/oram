localparam  CacheCmdWidth = 2;

localparam  CacheWrite  = 2'b00;
localparam  CacheRead   = 2'b01;
localparam  CacheRefill = 2'b10;
localparam  CacheInitRefill = 2'b11;


