

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H7mWcY7ahHbsC5LVCP0wGD/8slW9mpsbGEE0VMM5jNFuW1oTIAwmaf0Am4MEKHg+pogypb/i4TEA
li0scWnaRA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nubbWcKsG0E3+YHk3ZbneHkztt7pKlrGE85kCYZ4fh6xr5Ug+nG9OgbtODCN8x43wij/24qVCIOz
bFbOLO4yODqUo+L/tBC/SiM7OXgg72YPZploleeJaYccrdOCcxiOJdqrK+gSPqw9RTFyFl7syti7
VupEB0/tS0vu5hYSH9s=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gS3LmOGZLJTSCz8xGeAUDLvxqbehX4zHumKTewWQe+9Vb9wwIqVdMZomn+cDSUQrRrnQ0fHb7zNA
SZxnpb7JaCx8gRX+gPj6uCiv8fbMMNKdrdMFGK0hFfWpduVqsxfeGWoDLUcux4vf1wmR760URG1X
zl/9K9CHVNOEG5ql0l569khJ1SIeu8RjDRaRwoRWs7wL9JE//mDWQOgpFbGmw2TUAG+7NR8Rybkq
AQn9Z8oI77X1erGPpVEBGu+utcELBAgLIVAWkj5xjQFdNyW0k36+qh0DO2mJ97Lp5IDcGGbvzNdo
OOijtD5tXsGfDYE/nwrCIKt75hAPwutW3aigFQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cITIEij2pkbXLW6ox7EvJRV8snJxIrFPEnDh9TxBNs36b7R0chCbyMKUuSINVdcShK5I/Eaw/kco
oqTNzwHUb+OmXtpnMSvQjWYxDXskYxkldqh1fpD9UTsZdJQe8Pcg1XlzcwZDZknfalb0h7yBNHGQ
nNYpeN/lyNLhoBHjQIc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qF/I3soQa5iqvpU/5LP4m8lt9LOvVDLZn20tVFDG4vBucNIYER2tUvTFcP8jI0CLkrk7jFB8Lo51
QiQfJpzgnAUZB4amN4M8+YzUkzL5J9eyIme8fl1dv1Nbk7LD1lBctDqDK5bxLahDi2jzK9n/Ki0i
83TjUHPFuLLAWxh95BjWnojTLyqoLxON9GQb4iWTzglnAmUeHaI+bkw/c3Dsy4x29tvk/zcGBNpF
1PBdlAFOSlyBhTIJ10iBoo89VnZV+PYFV9crltar6qHhYRN9d9kW/0k78teFfKZOObkeIhr8yNe5
jdLWseiubvFarVCcPso2WnrF50tH6SWHtMw7mg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16128)
`protect data_block
EXWtTQrJgB4VXhmWPH5C8lfKRaeUXQQplUKdKdaInKnm5SnVG6LcthOJJy3xugXEN/oVwVFpisk6
jcqOXyp4UqKCcSfsQDTzK31oOljahETe/ANiEpsThd8dzkbXN9Wn5B19LdLGVfxyj4/31swxobee
JBBQAZfxunoZtLMY2PhzL4zu4ajbyYzXhA+7Z8AvB0Vr/8IiWLyT9Krr8qiLoZkrPS5RdciRTstH
vgRCZXK8lPzMOPofTRIdDQw0GtdmJEFtjjLGqKLplXqvDsl3eGu0K4pznJj7rGUONEAvTRuFhzAC
zJtIdWgjqHreWUzN33xcJYmjfUOFwDhJtdruJf2Kr4mGFjAzPXRzzusR2aoysNv6qPB6yN2RBQdB
huTgkq8/X2k6yrWVe++PEIF5UkbqjbvDnXGTDLk8k72HI3T3h3LsWaLnhBqFouDa5qaYGoGgY/x1
i/3M3XDTwOAy5/FC1wF+DUQHuHt8SmMDimUGqMVFPNqAaB7OMHCkW2GhMpLCYWCh99VTlHWtXlpW
syRYVYAKrjGAl1F0PgUq35DlMq4Of3MBnysj+smpqZ3sTU5T1rSOQey5GZHJA7OlBXaygDvScz5o
am13nPkviQfsVnI6pqnq5BvYzLQuKZoQ98CQOZePD3DA1mH0zvG7RBvAJwXb9u9HA4DjyQbxjhJ5
f2aTBCNdPjBQJlnZIU/4EXhSgSv5np8VofaySLE3kZN02xFnJeu8aH4/hW69R1AI3W9393ymaDq+
VfadEROVYntU7w/1VxNOLHE3OYvM1x0uBZ15OWbo99yPIXgTdxxYMjc4YwWNz2cwWCnb7Lwxy33r
9BtheKDVJrTa/btlwjADZKKL291v/zZDyJlUqZyK7Su76V2w9EgaqE/z8sZsYCyraEV2kvm99hye
7RLI3SJZR0lxp/KdARv/2oq6k0kGtHxumd7Bw/0huabfYScTJ6HaesvCBKrzSGMkSY7Jo/RPMKaw
nriAXJNhnZn5ofEgkTGFfVZkeFOAXpDkF+dZaeY9X4VyceqBSILqACq4LuX+2GTvZP/snA6vpWda
Ude+64PnfUjB6HJsmKhHVCUXZZHbuaBfWziu6BoAepXKn/DkCErUmHC6OFI1EGvMAknqW3BDP/Hw
pkAKCr/O+5Q4QZ9Et0NkmvT/poepLRIfo0UdyPauhOpn/GlAK5DpyoNrGQiS9zCKk2IYmw8pXwgg
S96iN8egybXF6WbEBci1BQaXenz6MXq9MGbUO1SMlITupkBS80xSyv9f7eDsNEGCVTYILzaLp6/3
mn3A+ovORTx36q/Ygbu8ZU2SHdrDUd5ydhWIVgOYwHNEEPlDMamkOLE2QOXrKjiG+Svb4XAGfW99
vYWzR5O8MyJDIDo8mISyx9UBqNOE9fYT1U7bqd2hjrG0PRFsvBaiXAsf2O+1MnF2TrtXdqBFcRW2
QWo3S9Tl4A947S5xGyAAVHGsDE0YlzH1oq13GflIPZrh6JYJFLTOr9s8Y6gsVFhDXA2dCZXjhQR4
31DSxahPDMkDaCq/Z4Pft+N5prDsoHHX1a+rW0IAo73qYl43PziYlbrfU8M7uBQR/GIrAgEbwWJr
gSWg/AizLZZlPtBFLDuNtnNTt9qpY0RrQ7q0DIYxbSh4sRTK62yF/71fPj/rjDw0U1W5QocJIg9I
WJVlgeWA83Qt56R4zGhDGPYor/EIukT3ByixUdKBsv0BUTZxVU0Eh77Otps65WWeD50ge6fWmu+/
PQuQ9HEZG2QdVVAKMZNxrZj3o3fbincz4MtWDRcFhJw6yS7eOa+N07SzubaljdcWzV6lLOPDrUfA
BSy3RAnz1mvJGAZkcTNGJyaVg/5a1qGeurlk/vhsspGb7eJgIX0MZP8Qq+mQyII4SOCg0SPRj0Nl
6sXOKX8eE4Z7gixrFp0/44nH5ggv7L5ueVf0D98lh0Zc6m+jEzf7leBYRMh+cZM1Sw4gZGQhVnUO
b722D6/4oCxt2/X6BlwxgJXFw5rhprBriNbe0qCk+I83inC+mvCnHSM7H4h4FPf4zV14O5Cr7DmD
g0Ok20dQu800BZ39DSevMHOctGTbPo4+AMHtnPYPqZ/kuv8vW414ABq+H/1w7dstQhirZNr6IRvH
Fiu4BTlB5WVsR08CLZbzu+A2LasRdt/Q2a/ZNukI8gMkL0z7W89JGaswbGbysv0cj52lpqDhd1jO
b836r4o10BbGnvxo26vgoukRT4sDa9BvNMxtin9kd9WmGagSFSb9+TazGsI2bUXzZuyK12L04ZpH
Tl3cdcS3zl5rYhyN236rcfsjjV/GmaDM2QG6gKJQpjSPAeqcRjkUAGoNhLUvAPkO+D+taRjxYSOI
Lrowx84cC6y9J9Eie0KP/BYdxIZzVec+sQZhJjf4jMtFF+kRtRJZA9lVIc7eLNoXyV4Pr9p4ZQHe
I5Njtw5K1uR5goRp/BrEit5VXvGrNTkBo2dVLBEEhpn644SG94FZ/f9pkLuj5MFtMlRzlyRAFyt0
NridKxKzXsJRNIt61cBPKo1zgP8Q6bjL09hU/ALgHi+kAP0PNN28MZ8PrBkVeVKONUnIod6Oejwl
G+C9EQlP5v0cuOZUYSDF4QPDJnupONzzHDj3yiTWZdb3Ax38WhGnGY4aJ9jHCgM+BbQb58jC2dDU
figBSOpGq34b7v7Y1z1aeRzi7vIlIzec/To1pDpV/k+5rq1iTpRUmHFY1ydJiqqzwN/ZK94PNInY
SzntdWALv1w+B54qc6/0MXLYBKRdp9i8DvSzv5h5AP/Vv0UpuwUjAH/w1giycFDcd522Zi3vol4q
AnLh780PsHfHatlreBx9bN8TGGOs8Q51R8RMCiSkJUXGutzb5p9WOeR3iz37sE/6bQ88XZB9u3lj
80ZgDbQThDiWV6bTfn0eN/Hhq6TZxR/8anE9DBKvvorBVKjq1DukTjk4t9K5L0U/iwZpnX0+tX3/
tjgXnJMipjCL2hXyBuoLaKisgWFL7XCG1rJ0GTIe+RtatljrkQjvJHDw6GOPooJ5DX9T6irZImhm
TtsEfd7RbRT/NebP18PzpVZulK/yRy/vRAsmjB52r4r0iDF1TvziS1dY4H74T4xZ0w1dWOl0XG6f
KfCyrMRnuHKDb9s78GKQUu3H6bEs+dbt4XcaObRISOWuBdxtVVXBV+747chVleb1WxOYL8mC7zVV
5BYLNk0UplBWOrHEK23fihFA3gMXqm0ogTUcEucj0OfctClcTfIfRf/452+2aEbqUsnP65vy/LC3
9ZGdl50n2NrT0FVFmZw0ad2KhEpl6iSbjudxjcUJKgQGILRd6jaOszZT4ESMkcP1qDsFm3HZNnKT
kBGTyt2SRsQI87XhJpC+cJZ95EXA7PqbEXJsCnLbIPN6UIRtKtGBIuUobEFdHGQijq7nkGGpnYWw
K/X0ZEpNpNidAPoihnJh5NiBuPj2/JTGY3u4TfrYUkPe5iXSypOor6YJMDd47FsrINJwRG+3HX5Y
dOnrVH3GVTAiyRA0o1nAYPHqkL4r9wsCp/U3LGNhbfSm1p6DYR8T0JDaobEgktVQAUy7MQJsF+FR
VDFwDR5Isk44ARTtelgUb4sI9ciEnfFpIqdgjCM63CCb2TH7/xYM/8x0zhm4nq1QQqcwPYccr0P7
OIi4XzE219GOcS4jYyX6hAx6yBic+TcoFr8Fz7AMC4oOJGMYcNGMlvgkhSmWAtAtCSEpRoRRO75i
2x9FnQif9XI8ifiEMhgLyr/GFV4qE5dDyGQqo1yE6tM+xEciZCL/qhQKsS1UcccHcoWuacjlFBD2
f+H8iwyrkBSSLHsrhP/kWaj4g2ZEZnABiVVD2gxYN84E9uPrIAw0r36/P7hYRGIb2KT7vwUvfAWx
qUIBoxrB/5/7Oo91E9YVS3MfkigGz0bPYpVk5Yx1jqrIvKvjvHCQWNXUoLBHs0xqkNSL5nNRDrMR
sFl5QqXrvMdPupmy7H1c4lsvUClWTIvgE3Qpnz1ULP6BvOZwZuV8shQdIu7Heegxn3QiVdqMxpOP
0AEwzk3aOCvxWM2y8nLpkVt66Lpa0u+TW0wu2oGWF11pSGXCZZnqY0KVhtElCV6dxF8veqWo9/8J
zqzX3wQszidegDlRCdIlSRLwEXo57rmqb1brvbjmHIH/VAgrYkEEIDq91TSCVNYaPg8f1YY/Z0eh
3UXgwseDIfHpWeSLRVVG6JRQ3Xr5B4Jfe2GIdmVCD9c1VoBup7mSbybr4XE7LIK2fp8z7qAgNB24
naCIV/3UiRG8qRxN5wSqM+DkS5r0BwcDd19E875oJepAjcnf2jxglXYzYZ9kKkbjG7jGkkmdEzXQ
aaZdVWIQj66619U4WSMbsLHj+0/pa7uPsaJYhWRo9I/CMjrTXjsro11LL/6iOsDxaWttIlpHs0ur
5Jab9JbERqASNXIxcwPrTZqKEKNKtoWE+mqr6MKvWgEk4HUwVmQ8RHQD6ATjzklJX/YtXt+mQR7d
L4Bds6KE9gvIJuIykIoDYc+eOwYmHryNtQ1ip23UBwSBYH8SU4N8XSi7acbFRAzWfxRHBfUdT6Hc
WBpS0+WIc22brmSLDeoSGasgkuR9JpYzbh5YJTQ8Cf4ULCToE5hBW7JVMgH4Qf35A+CYejLuKQet
xiUkE9gFf8U5q6n8FG6z1/RgpwpHBFkWmE5AVnqS2SUyRLbyIOk+Qa/7EZ3E/F5iVvJBWDs08kDG
nYy3obpu9lIEgHcVN5Bt/CPkYFkxkCPx3VRnxHKipqlLrYafM3hHLsLkNuQtMZIiOcibHFaGJy+3
1ZD8XJJYp93uEUpSxl83YaC1Wc4c3dveZvNePIz3Ze1+3sxWUV1uujBwu2o/AJS1IqHfD4hP8vrm
r6ojpYTl5tAYADMSQ4u9Sri+y9DhnRN5Hh23HDt8Cm5DnltLyIeq/1d8t8UxPVbiP4uuXSNR/crL
dpJCJojf6UpMj5yAjhPTVT45rRXzi0tF2Isq2DzaIT0tvJC7iXDMDHW2EJ0yG6LvS7c+XasSr/tJ
9FlBROFGPse7MGplLzYYrYhl5/Gs3eecT2kGjeWpwQWutSTCJtYIdXk/ujHgE2gkvCJh0f35jTi6
/aj3vN8qDO+HGtGTGzShlq6GLkkzZDPodDfNsNP8ZbzAho0/YOEoas3wpE8qb0j+G6M/RGOwg4yf
d4rjE71TxvWfyZHMa/qckj5+Xm7fGT3q1XYlwo1sWRnyp7uh/NMcSDPWeLlBjcoo4ZLPBUEAM5cU
dOgfcNQYz9r6AK6E+kn7Wzi7rYQU5OblOwC8n8L5qTbln0itjKiTmLtELTYcNxOfljaSmEsgVKAm
V2QuiCDOtX6AvevKObJIVFq0caJ9iNMHh01vuL71idWSkc/AYx84OEOpDUWiD6x44syUYwAyCUav
oQv3FmrdK79oyzBvKKGqgz6kxomZ6vQHQKhJdk3EQ0A4+UP4N/BwVeOL3+eSVpSTKPIehm4N7X0a
F8n/703KzRqFJH4e7CB7/+csGBrK0Ma2/sU53C3jhLDr7P40BmmsPiHCbVUrUiDn2zLKB1diBZH8
JAVQ2BiQjQrftr/qgOfILExF8xt2l6SpBQC+CT5nsPz6PKbLWyQADy6hLUiF32ou7ZQUyiFKnXh6
Ec94EgQnvH1O+fDYwBDbYncjKHzR3ugw0rNH2Gy3oXsrzTAQLwXDV1dSVNIcnpPqfzTxdkWN+G6q
0/ctNMUxTmm0xj2hRsQAUVukEh9uUXyBiJGzAaOYPF9m+zMlA3XWBsXHEBKcL52SiJrBE1cWNm8s
QuaPJDSWOaNcG9G6G/SPL3NZYm9H080stFO1rKDJLLzgTTeKE01hLKwz4EzRxS5NR60HGV68WQny
yk1/o+QAxAfhnA8waoxHef2uU8BZxuPney9VWY/c6okxwUmq66JcO/2jjOs4YimJzn1IH3bc7GkF
C1tm3v5HYbNJgHWl7jbNCvJrk+J1Zu7qiUAe7NFJoUjmgdaCfX8euKjpcV4/MR7bN4LZsULpY4e4
dwfxPI6DwZz1OTsI9vijgpNwXhRo+On+C8ltFgjr9z6rTv//v+fJs98pdFBjkPnQGNGnn/CEoh3S
tjF+kCvwqTrWTyUo3JyZw5SlACA+qjYd2NQcPvGGao8NXG3phFU+irWmrO5UzXDqGK+Rz9uBHo3/
f7VpmFQ8VNqDLqcNRLzliC05vZypdSBjgMIRkLJo3OvijOAVT6Bnc244jlg4VeK7sTMwZssuys7H
O0zFH0S5I3NIUI1y0e1QkIz68Y98L+sidPF+oFX9PIibwoTF35BIzXAa1fjLwQVmRKvZ1WNB6YbS
H0oCaUyLd4IXIJS54mOx5zr4vaVZn2c6BfSmCJX2t/ndRQmQUy1vnZdzlYgPDQxNjTQl881KLCXi
+Vdg3WwmmxBY0VDGM/rARQJxh7HS839UF/jkALcigZ2GPDxc2N4cSPsj2Di2C/eJXiqIanvmG0Y4
6zHBC5TedCQC1WQD0AGCTGU74gKg38YSP/BFytxyoTezSV5Na77E1g4Raqs31CkKXeJb176t+/pK
SSTEWq2fVfe/PlbiFM1jC2Fs9dYi3Rl4XYvuqYtMc3O72XCHV37vjiq5HWJQTCjOs+4UsXjWAKx0
SZ6hPrseOGMBSK+FZLVoreFchXeDHJTh/eJ2qi2pGJRZcD06Iu86AigWASRw6LfpU+eJ8LYGeaRw
o9yI/10Yp325P/7+2V0ytu21dslxZL+wq3PF3HCi9ZtFuCqcOlaaqKRNfA/8cGNoPuCQLHBhMhLz
Yxo2/wshjVogF+6+oi9C3pm3RftW1eHnOJ15QByycypgCyCqkFeyj/eo2W8b7qDNZ/ptUGXrVTYD
fcNhuHyt98RHVSve+y2noJlaknFtnh+3yZPeWQnyc6UxVzO0lPdeQ7RVhBaOaXlJEE/XGNWqun4Z
WhRaIVwckOhrBy3+slNuI4JyskHqRbmJHj72YsofWsZUdWBScmJUMg71WovIdvoKuzkmlZjhHJLW
7qpsQikpEeLclWKGBS1qHbdbpfYNVH70jsgzlX/SD5UgWCw+yJ12MS0oTlz1pi/u+yiUA3BAnkUu
exyoU0/cI0p5DsviLU6CShPP7lp9j36ferKPYGDB4rDw430Um2ONdOPDLSeaXPpau7XPJmOVjQdB
MdphbAaG7dW9Rw+iAPNwTARmMA5IkBGDGDfzo91XBNvw8qxEt87CaM9jTgnQ0oLoiY5k9ipjxkkt
pxT+YmkQCvi/NHOdueR2p2+RZMb3Fq/Q/TPUOjszlLWjkiu43uQoRugw46Y8g3Cs5D2pma+YiLQy
KGLYfGf0VNqo41FQ/AK4fU7/sbk6Nb2VA2f1FbnnSghwwLfTNfiBk+19p44/GzEeioNGNMfYg2BN
18EwO8/iNZPN3VQ4S5l3DuUXRn8kQ+5VAHKq0hfY2rUagv1OsaSGB+olFR2kD0xa6YzUONJwmE8f
k0IHbTdqHs2NkifdgdbUbYUcvKQbcT1fKllMTGEH7qnuMR7WZwQ/YygNpJdjB/Ayujn37cg/88Tw
hyChWI/tSosCXmyH/wAZ+snYXeAUEzuu1H3fmxFtCxbOwQ7ORJC6el/ngimIhPVa7h4d7Ned5ncl
2jwacLlanaVoEB2ZBCWs8SBzl2QodUh5Dsm8/8NLiAS92q/MMKH/y2821aWmnZodSs/cNLjKWhyA
3V1kJMlcMJYrxG5BOtYTTiqNwzlNR6vaxdlj+XwvUIu9i8iRp5+Z5vCG8KD6ppOjJWM94Z3aoWnU
CTuS8HmxuuxsIzf6qtlllfvHCXktofA/fpvnbA68LRTp/0NX3VncSw7XI1pf0fXzDhacx1tTX5n4
CD2uz+yV8CyE2aJjAORGEOcmdDynRRauQ/PXggg0UP09FWeRc3fXR+s/zvobM7UdRQlNDmMHknEU
HfrbdcbnhOM5O6KZIW5Kw63UXO2ZFtYqZaYrt1pyy4t77kW+HooPx2Q0rAYgiGtHNkSaSycSBt03
mvB2ggj+3iCK1YNaaTafWNrT/PIazbYGjhqh0uj0Z5Xg1YCSwSU2mw98Lsic53xX9oVXrhFVSZ+W
Vb3narBMmPHuu5cNPtVU41P4ra4bLKSefxGi21VWQn1ByU1N5vS1HIPhvaQbJfV7eK6pa5Fc7Mk9
MctluJ7eg3qQ7Qy6+oRyC7RonJr7zh8f7m9WpYvzlq6ZauLFu8ML6K3C2U0gMrNU6896ls3/NKSP
TKNQxk1fqCrVewbPEnfvB03BwMVNxjFXdgEAxPlh4ZcuA+vqQZjaA7J8jNeHJETkRPmPyWPR4TiM
bRv/WDKAJiFoShsOmNCtsEDNqeFwQxl/8yx8WJz3QZEs2bSrSXED/OqlKlNBEF0YGRChJzlIFUfR
+yjuGSAa1w89a8jq40gAKkNz2fyyQufytCpKY4zuVhGy0g5RK2WcqZwmty3Yt3rELyhOZFL+9Qls
1C+slo4NYFjd4e/Xbsg0a3mivw5txDEGGsXOkAuxuIQ63fcLQw9JR+ebxVw7paOdyK0XDIYQuxKl
Tj9xcwbG8Qngw71oIc3F0pT/+Qkiee3s0QutJwhfkxprYnHLYPeflSEp2iWrO50oXzptNdrUE9Pq
y2K12AvKFxRrPOFRVZr1qu5r0voZEvkOPDPHZAmf2eL96XgQZo+sjyy8bzicmAR6wn/SYKmzu9I3
ra6zfBX0CQz2pL7SOlq8NvgKGVtdj1o1+XkSpn/I05cxszdJdbAf8HZke113n8lY2MGAjlwjpV2/
SCMXrvapcl827T/QVdZpJd+JKCA0CsHrWljuk+7sOd7Got84A3M+iaj4n1peKMiv981TJZRRaS6m
vtd6IOxZumeGlZ1M7gntSbBv0JKZGEs7/g8KmGVLWn/etfeBc/M/c78t8tV4swoHvMiG8jrNUwTB
GF5cXh1o2rKx7anA3zE1Z9wcqSGAAAnAgQKHCNsz77sVjL6I+9nBZXM1suk5ASWZrzm/HwB9YI6N
kUxgld+JYKhMjCaBB+vtnprrfmFG9Kqw+oPhtRIqfFMfzoXqxjcZhu4oR43qrSARU8dnT/X/iqGN
IFm3/tXEu/JZILN4FeEdvh13VnQ7l+vfp/E00OGt2ySE9eZt3fltpew3U4ICT5EgoVJz0t4UnOj1
TwRvRdY7WJH6eRYVcSvL0BBnToCD4Alw/Y9Ew0Jiwm+5A6LsJU9KctXe2CXScW/ppVzgv76TqGPR
XkJKsQDfsWzUySh9gTS3WKDbQwU3YeJUthwCnXXOKJOEicbJwSyPjpx+bHVzdf7N49XSIoR757xG
hVCTxRf15SQemBo8kLFdNuWr+PZbJwHWMcso9ZDS2KkryfySsiw19UBV/svqdjqZRuLQSV4pfvxn
xaEMgnh4Brt007OcYW7At5RfH31wBW/sK5dkGszcm7mB7Y1ShMNoWxLpw5C39k0Yx7tBpVW9EBOt
0fkEW2Xw7OHx+FDm+UvH3db9jQsFQvpjZl+jWe46VQVcGulV+AvSN2JNrx6toP6yRNZxJJX/CoCt
BBChubpcBfB5eMXCh4yzPlradZODiEYTmPSRu0hNEF2Kfq/doTowa3JoTXVXOgvwfmFkSU9jNicx
6FOf+ZkcJQeasurK2/ON8+ncmrKZ0pfBPu+7XdTIwsZ4He8GbkQkYJEPZb4nPCKou+VqFWnVdL95
znOhL9opS1DwAdXc68I609hbPoB7OEEueFcQhp2iM70/VbUOaAFYbthQc7J4K3ows9WSb8Dkc1zQ
p4HVRAc2vAIDE8otzDatwu+4JBMh6ics6z0hJJCC7sfpdoivUmApz4+0Mf/rR/TlXU2zahhhzO9h
lT7ejMS0mCFy4QsHfVT8olM8OZKuwXOyWTRHmXFtwbRKtZ0YYLMAt1Pa3BXJenNRBNA4tT01aB9X
PaREgZDQgoEeDzvOWRVXPCWAUjHfIOxXa2JuNXHi4/DEFZUxtvsdhgPdjeQ38qRyXuB0bIk9gw0T
UMvQAwfzGD6Lz5AdlsEyhWW7kiBu2OOQxX4cb+ExkdjZepBE3oP392OuC56OJxL2P2hryuVrZYCH
FxWP3uOY7eIr8Eor1NNHdmEN/jfUtzJMK6YbaNoGJ/hB7OQ0vA0iauwRUGHDIxXdlcmf9HtjGIrJ
5I7xtoscsPp3q9gaXq+jAWBk8kYDPfXv4yPTgHwmjobXGUM/GLnIwBmMuBapcM+LIQz3Qv/b3hot
s1kUMRyuA2gQzCHz7aadCobQB9nmLJcMASsyakKwApFRfjk4qjQKtcqxsTH0UXtcORBXjjVKrmIu
M6g6yOkpHdwQG/5us59cSOQROPw/zDX+of/ElygiG81j3+8qiCJqv/sohIxmM2oU9zmQKpsHkHvy
iJ+kvHLJlqlCPTgJDks549d9lVeorvAWAWw4lYcgf7ohqM/aycrqjcjcTDfPX95lGKd5fydKM8CK
1wjchx0NK86IsokIFH3SWBRIPxzENZ+QVBV1eBkNWihoWvJr67x1physjVyq1wLi/aPfpKzcd5+q
shtun9UzviiByD0dTq8WEg6Xu41Q56stZBJROUXI9PPGVNQr/rBH3QYx6ZsypO8W0dOE4UIYJ8Wb
UL/nFcuM1fLOZ1wcvbXoVMppnGZdw8JqYx9fSck1lVceHh4ToO5XMARM4U3k/gWgP7pD41p52p3Z
7fM6iJGLnp8i+I+v8W65fyiJJecoOlsf+cFZq2+s1H6diBFPkIqRvjkFAEPaVWApZFkMERzGvAcD
KGfo3hVcIe5q8Uq/5oLdpxaKrLrnWJE+geFfuj+sjCsubpQQI2SMhJGoYtHPXprQIaV62taL6oMO
WwN8FoBxNFwgNw1b4dLLhDUE2G1k7/tbkeb/85/nYmMoH0gFENgyA3Fs+22PkL7Z1D0i+xcEk3e5
k2jOJCkoXoe9kSwhHPkTuvGieS4ta6w5tmFlArFJlClXd+zIEZRDxrdE/zw+kwlN+52ojVjpQYv6
Ovd+gz2SJI4NPdqN1VtfxWI2G0jW7YBMVS2EzB9H03kOMECl/RsnsmXwcpYRUbrxj4gxmGd9afEe
+Vur5JCU3KroSLOewg6lz84+Vw5Sn9M9UmKyRozxFMEInrU3hb7Q6DxE53SWk2knpluy1PWrZ7pu
/N4k9WQRZxtrb8e7l0Gfm2sLZkECOzceLRLi7WpnQ6ETKReOdqCyI0MWqvhD37GstPPMNZD7oGwv
B21rYRJa9kKEoiadfcRwP3aU9SRcoaOQDOmAC5YQbqE3eRxQjGDpvaX3zu9McouHLHHZQ6TRUO9l
1bQ0Gc8Iwt4yWBgptFAXfAekDlblvNDkvI5Okvz9kETMjSXKuXOcL5dyDkfNF45NyteCbNBY8OJA
+gzV0kSDyS54f7UxqzTnQn2rbdXv8NmCD+QIYZnAnIUeDSirv5dj6YPxJKmYXhPs8T0PF5GOWZ4a
tsgQ16hc8FnFIJyEl5kK8mRhN94eHI49aaSpPbEcJ22FeA8uA/+JhqzkVYzX18/Jb1WhhN+X2txw
3MBAl3HwDmL0Tt4J1q9ILCI28cRWzTwKCw8giz3lCkPb/jWubeJ7CWZJipFlcVzrSjKZT2NI+v2r
30QRr5GeC7f7BpQj+E3hWyiETpEBbXcSpVK9nY1Xm0va1fyhI15dRkCq4OROAtOiBRO8wfJZWEJ7
GclGdgnYDqvV1qWj0932dmbun9Y8fCW4+ZhJqXOPyeFI8kWyUQrpOJ+/gSNT39Q88Niv1oEKFwok
5G1i318Jiii6EsCp9iSPxXIwMrMAxQ5LxnX+MiraezmSy57lXR7FDkiMzZgg6iPOkM/FLaHU+mac
I1k1yHNxWceF7+TbZ6H02klYX0CV/xEuUJOu2ENtFEdCSip0ABk5aRaWRyzehZipsMt7vNlrxG/c
3eYpsqFE0nC2b4B9dgRQRCEQTWO9D7Np1eSGzMSWrRPznBpK3EyWfrEwhPIRf3ez9mS86OIrhT8H
ZxsvTUO3+bvivmptMF5BehqgxYj1iXs3bjJgLDKSnpbKU4dPCT8+Qy9HWBfbCdDNTPrT1KCAVJ/4
uHj6ioqTxpYbL1GmV6avsybcULG2GScOOaXrHJ3QdjdPJDl3p+kPR3rAY1rMdkOvZPBCe9DCA6hC
up5QGwcm85jfwFWydW48dfO4Yhb+t55tpulKiYpmmK0nrm/SMl4ZQiGN8MT5vpMNKQJbaIIG39mM
E574pmLOigQEl1t6TXQKsvhjcl7Ox7iGBvC8jMq/2A7yFVk9EfLul8lFIQXQ+j5rBKktDyFZ1a0u
3Yg5cKhdTb/Bb4qZI1CLpjLzbASH7H3k7KS5GLCeVGWJERARiW+mye/gmVpCjGj4rAv7zbCO8SBf
DlJnt7G2bTP8fMdvU3Rk7wTyv3pd0GU1RCHxIBXrJpnbYbpqvyuIhKx9QZAbzfnsglVmsDtzjF+s
Z2p87mmsyYOOX+uAjIhbbw29JSAqB2E2BufCovyLfkd80jbsVhh3w4XqnYgkjAmWgvlUMhxZFu2o
9KqFiBxdhka9XyXrqpjDahzbnXDCA6RGwCIdRzILEq3HRso0dO9s69uEWX2BYqII9Qb4TH12fTrB
NX4EgGg/PKYZNp+jJ6auvtdXIyZfiQ3lXs0zeP08D5oko6nGCgdy51qX5HYqebdztrcB6rfpPiau
qDBgHjbqCQhQxn8cQa6kNvwx22GKw+t6j1PQpWEOohxTtfEskdRbSV0zvXQoJP16ckg6Doeo93DV
63DF8188RylJv2psf6xzkKV1n7LewRHLQ5GUzctDgv0+jTYRFVDjlxrmwi1JpKiHnBpaTyqk7lYc
girfx5jvD/84/HgOodgjbj+FNvxf3ZqjDq5C+KQgplJ1OrP9GZer2+1Xk6Hzm7zbaXiytLwv0UJv
o9uk+lp3lb2M7my2hyVQwzpj1BT7q98muqhZmbJLOFFPZCP7ekZ6BXYN8YJKfMy8lM/YsGTWbwiK
qFDgnJih59/MIxqpnVb5NTqF6VO0p5yZxzVhGhHrlfPWcixhLYg/UoEwL46idMGBOjVlgZGKsnCz
5NSaoRvpatdre9JkovcHJiP2PEiGdZS9COluXtUuIoA55VsunbwXIsX3mBe7MVCKWscvTwrWwTEn
t9LSw9DLYeSJxVq1uykUQIyHZcC3QlAHBajfvMHisaoeGmP2MrUZeUgplNPp4Rrzi6VzhooHBSR4
mGlrb54Pt7nVn7gkrRzFfTCj2vmGNvlxac9NcwO29LgKMKqr7yWXrOoe26yN5EqhDvf11vja4Zfb
J8n7RKTlxA/k/hdo0iY2K2xLsztWY8By8uPPuOdXmrx8GSzqfbT1KXrOJla8lhKinFqaaya/BujT
VVOqiDhX5b8C0a3tP8CDO+iU/fCJpzublVVL5qtT5raeQg2pr0Ec6gPe4I/zmqwg47QF2NJx2MN8
3nIT9fUfbi3sSCiNlb989QAGIqoAGUsoKK59+cH4xama7AsQNTjVjUJiMNEpwPwR2QScFDMtmp4C
Uf7yKlwKdD7B7YrFs9w4kVNTtwGMO5SoiWk6UOjmqoTh1VcaSH2zxfC3JEBkKMMLmby/RfwvNTzS
3GJPk23apR0S+qA0vM2xgYGkj7StovzNGMLu4SFEhCU5fyeZwzN8b9We7igpQb43GLY+r9xt11sJ
5ibDK5w8zkjFy7mM5C2faDn4m1dbTofbGrQGbU7y/bJnnP3avOv29DO6CeJEKkG1kWqK6cq027/s
uhvWaMBE3pVndt/q1/dizOZ+vBY9N5e0U16BspJ6xUkkgtRzYV1ycQDxSFd2LNgxe6uiu+5KUknO
vvUdKe4Tw5U9M/VvHqyjSexBQBWQhQcyCSLWziEg2A9efHQFTSUrRE5TlUANwnaxXzNPpXxiSiZu
CekPK4jWPQ6iPDnglWLmmOAnbBAKg3LZwxzYipJBlecuOCF14pfRzsjvZBXFhppgIePw/ApX3Nlx
GKITr39JcH6nhnjgX3+ksn1Y9Bz8nBrqqX+DfGvkW+zIILUFlQhg4N4yteR/uX0aIwe/L7GKO0Ee
aVmasC7YsBtMbs3TuOaYPwEp+05YwTTXpss3bW+LCLRE+VD57shAUdG51TxsHG1JxCOGS07RHcXV
o3/0ALCXYEyT74wYVJWQNKYKKfT6OnM/nYfpwzsInXuyFnoignSH72FoGDL9FwqWqwAiOhBJwtl+
72hqCiNVLc3Y71LKQ+dbBR4Yg45nAkEVf9HgycSpuJSsx49z3Zdi2IxuoMaMKE5lCMevkA0wOnyN
QkxE6CqIdrCegbwY43axDTlaIzqE1Ur5ANbXMMIQ0s4Djvqv4G54SbANeNuok3EipEFIPsx30tIM
8oaV19XiFWYknQBwiNPfkCCm7j/UDWVn/gAf/SCtlazUfE56Rk6d5OGPYB8FE7dNh+lzg5B1j/+d
USIi03Qn/XQt2IXogWCydjERrZqtls3vg+xG0tCzLSMd9unp4NrNVp1hHa4fV9a+0J7Pc38zGDP5
bzpbxU4EVUIGM99JdnE9joDB4+oT1RTUcemBLNwR6BzupuuzLhNDC77biT2WHy0u7223jeJezmv3
LweTHm2pgw+I+rCoJG0sE1Y2zrgfzAmVgIoJaodbK+ccTe5OG5wIHS2syJbwR+fyWC/tM7lknF/N
fAiVUdCluKg7mDuhTS1EDM4knfvtgNgYC0uUXDOXeEbboNepxF4klnLhsie5dh3FT4hSpgdp1A3e
jVQVkNcAWaLJQGxAJG1wF+QO8ilBNX/nNayF92jX1PC03deYX2AMh+bOMWmLIbg8SROquBnmmYda
XuAVRrGMTV0r3btJDu9CWvuTs9EgO5/7uo71+4C1uQQMstgyLa/SeP/aDsgzEiBPx9WfYXdvrtC9
AvIjN4VFqwzHI23247QpBZ5fn8PuFLNX5+bVBxncJKwnIlrELTesfjJV4i/GUX6unM30I8tk7MKE
plDlgvhso/LZTZYU54HTbbV6yqqVVJGi9l3Udi9ToHx9w5k5N2k9InJL1s6XRwbgUrtUpykbk98a
Cy2qj5N9OGE71MB++LFwuDv8zSZhsqotfGitZaA4PNupwmagGtJVTnruI7kIU6siZDivKK4hw/Ut
9Bfy0cIKlk0ctXU7VP+XYMAAWRixvpLaxeF4/ct6XqlhZaMQU+vqn4xn/tb2OT64xKC4L8hNkpci
ogpU5ohkybfsxl9WY2ImO//RhrVcBUisFWuf/kEBtOZOrN9IvetY0uwWZPxnCASauDn4yuyzVy7n
UZyUluTtPZqflCxSsIY6rMEYL69nHxx2+BzPfDLhgXfiiS+hwgbHtvQ8ISX/d/yUkPqIUmtc4FAN
06RuCEX+IjIB1EQbOEVWwG/mohYeLlaM0ptWAj0r91t2rzH8ysM4Gkkj8FCNBMyJyhkzN1BzBrg6
VkRu88nLg9SVPcjaYmG6LPFW+R59di+NWbPFR4Dmx/Y/85cAPxhfwi/Ks8kcrHGj9rNBSN+Bls87
iYLzn20Hp7loXfTbkgtMkClEQXab4IuvnO5yQlZx8Q3majdgscP7jl9d8p41Gaq8o2kWBCLEUAnA
UFQrl1cjuhlCh624PeS8do8GqlaCrL9D8bCBayr61se9U5EhA3rQJHD9/6oe319H+ah/JwuRPR3i
8GF5Kv5Jh/J2mFVVNLMHYCDbxSWG+Fklq1kTmKiXD+MlRlwlEF1I8Q1IHZMvdup/7SjkX0y2bSX0
eFb2i9+TvPyIHUkzeMiYBMjLwPt8Y+Wf8yxVpSMJpcBOnq0RVq8XgrzhF2MQLa9T2cimmoKf76g6
IiqoFsb5eNHBkwmheLFWlXSqtAhjsVsUmxkze8ZwLRfqbC4PosuRxTC/EiottkG0NBRC5CcoSNFU
5+G6OX+YA1JFbkMBu5q6n6+HjrwYIZa80FDEEZCLOVELPNxdepkC+ZVYMF8zr91tYu5M+P9jEege
n8GI8G8W7xifoP8K5xKJ3TGkyWRIxeaGhG381xJt6kRsGO4iXKc2pC93NkmGwtT8s/cuxspUB4Tg
e2ajrc0nR/gkZdkxnZg/yLjNjSzqvzEP20u5ilOcGx33vIyLSUZPPDndahHbTePLkVFRZ89CxIF2
l6+GB+f1VJu242yI4yHiK/bFAySAMwE7UVKsfOQoqThsOxhWrAAye5rXI1YnhME7sNvGKPtuvPiC
jrrLFDq6BKhDoG2PYqZfAi20MpN4/q+e75g2DcCZt5OrPJ8iVhP9i3Turc0q9Pq+N2sxuBS3QHFz
D5hwnorq82l94H4j9k+JKb/iMCA//O1ObaAXsrRMb1vYm4Dn+yyqEj01lSYDJmueA5H0BlCVuOSI
dfs5QFDVGF9tTZdAUNE5w+tOEJIF/STVS8yZW7HtDq0WW7KRItzXSuY1rVV4ZgkHza+mmHdlV89T
oyww6TuARKu4zXzm6khRn9L8K7BHsjwxUXD0sOCpl7qoDcVZmcVJnfMKQoV2iXealLK/oDodGCJL
aS3WVVcJqmkrEXPpPqD53C5yZZoo3Man6d/Fcb2bmTK5lMZhBjo0dwdVUazM7GrKTxelvU5Ds2oh
EYwyaQ43BDZonjY1Wyoe5Eb//cU1nqDSqcXNKKY0jDVAweEZN1mTp08qiqZoWbX/g1LEZO7XCSHi
NWG6zIHBs/xMbifcy1q3FBGR0skNHpPWB4nLVJ7GGbGTi0Ov3vL/CuS3Ut3mSaMVxdQ952QOh4ne
c9kA355ly7By056l12qZtDPSk3mnUK4av1bkiDj6uHm9FpsQuL0sl4Us11d8lRWGFowlBNlRIBeo
OhZfhUQ25BRgk2yrhQv4FtESYJP3bKP/5lZ+/JbsTi/AZsD/pWZmPeIaNDcWQEzLFtaUZmYAYbRj
1NZM9AsqsWxX/PVrbznDj3dnWNfHAD1vN6vVSYINHn50hqufqahJjL1Mma8byUTPmNptFT6Skhe2
xl5APBJICelAn/s58FIs8PDO+TWAKyHrAHhaRZphPJiqeMS70uzrDbeEyomVLMZADaF9pSfY0NET
zt4ky6v1pH75QBq6ZodPpDb4qKtqpEiAL0+3CETYBGjglLgC05PiBPewL1v82vfAOgJlqqxu+LFA
ZEZt6333Os1g+jMrvr0md4ag73CSxW8P5aTFZRSsmf4VusbO4rIoprYEiiT10MixsDprwbkFcgFd
+Cehxwx/IEhhDnX4M8N6Kar0GXaRtLznCL7xVZ2zmJrZ5QRfjg+NnKd2L2XRBhkjEMYUEetzXuP0
qvT3pjA9rGf6dF9rgxbkQuztEYOLRX1Dw0ar1oyHV4Ya+ESr3N5T2tOKpRyionhLk/mTY2ioJJj9
HjFWBgfZKmyJkItK7DHYTVZAEp+3/C5VpWh0mpayuFt/eJ5cA05kChvDnpk7RoXgBiaBFCmNF1iN
xZSru4fL4bHoMNJJqHCkIxyK26HxedkYw6zg6itAX3CXpTqh4n8593j8ohrYxgMFhEZVBr7vzxY3
LLXc+9ZRuWwIh9ZZV7DozCJnsphic5bjPjAU9rc17Bmo3v/EuKk3Nq+3GiKZDTXawQpNioCa+X0a
slaEYHv3ZCbqbDBnthiONWpCMMgaZpvQCrA39CGcksjnYOikh9T54GuvpuT5DyLqM9gfM6u98+c8
jX7mIdbnNbBx6TbWGSpjNXzEnAjujAYdTJhLxVY9LIClWKnDotwtLMB3E3rkLrqiTB6TUdqLlZI1
CUQ/drFc80hqqEAghdQdZjysVdJ43+Ym8AN85JUdI7NRLW0TgyXq5XIxb69ywK1eI8EriKFqlxAq
TahGatSsgmJQV3ey0HNanGf6QpSdL7wzZfa75iVC5FlmpXPA51ayZfZHYUvXyWA0TjBg/ryNkI5b
YEqUn+KlYcn6EYagLqAmiCdAR4MzIym2hTQuL0iafbGSa+Fd2IvSopKSUWyqAYfjb2rv1OV33fkj
2uBI55kfRdSDgctayoJguu628PFUDEgkXtZbm1XcDXxZWghBiXl/z7fW9MXJXvlkzPKI0+ltxh/o
nLfFL9ZdxumRT7nmZAYSam5fqwCd3l3M9s/NmmZcaAv41F3QEOXvR3on1Zl6q0H6pBAUSlH+7Vge
oMvpma3yGzryKeBBAdASMgTVD69bUcUYlUHu9Db1VFxCx0OMfVlL5n7Ao3aV1mBE9/yHf+b+Lykd
2vciVDeD+A05aZES2lPOXHMiXYv9+lGvG/RBXhXMAM0KEVk4nJugaeTiQtj1F+l/PI7kdF7WHAVB
axspOws4yiCtowKh58gvNklcFaWQfoB410aKKnei9gEREjofeT7GDAoZKyxb6TCa4ZQ/1SRzsW3Q
622QgbudnAP0oQZAeQMnODQedPzmWUQp0wJPaEN6gZAo+o7NSDnLfXjbiuhf55dj/l6WGUuIC+AA
Gn/cV1wQSHp+r8AXW9HLRZh8at+gtGfds9yIvvOh1+H2TVG9MaGECnDgtb0NL3a8NXaT8eW+DqEH
9lw9FmSww3f6krHfUkTPo9bAxjYaH1tRBSnntn9vJNu7LsQcgzrQarxYziYhfj2lKbTzgkkaxuiR
0+/Hohf30T/wGyb7BbhHVWQOZqntndgTNl0qCIJmiwxJgOBVmLQd/StpsDRENUk3vFYogEgmYG3K
RHBYlnuKJOmOEIaUKd6uKxtVmf94NHm6oW1BB/1F+Z/D68v2orUF+zb9gvFnm9wRTanpiDiFKYXz
/TT2stKWESYZq5P1GFuQqxcW4kGQsx+KHcfSHaY6RUXQHTIRBF4QayEOgQQS5ovqp2zmNgJ4lRSj
eeUkLuAlmz/jBMND9TqrfR0QY32PkpdUyUMhG47cHVpNckrUYeoW5zJZ6tP0t9cMPprrSfe03aVq
KviKUqF1lj/0ORvN3veR13REKNqW22x/ks9b1djnOH7anBhx4njGVnvUBCwwL/rcvIMFZ7MTpIy8
FwzF1oKd3zVv55FYDv4Pm/UVRTWNC8V9+7yuLiZlGduG3JFu6N8BILcWGLV0W4n/Mr5U2RYeVImL
7juy9pOgvUO/iUJcmRXf2GsNy9MCmHrsTHnHLsSXipjDntySDwW06OasQVzOTRB6Hy2ea73u9UhI
hm2shEhg4sxXI74ilpQhdqFY7UgQnqQgwAbMI82hiKXJ4lLX47QlFShZrgR1tv1XppnaepYS28ef
2na6vVWWp9/oH98COn4WrBvSYnU9oj326BWXBgHxW+Na0uTCexegw2Z45CrKTifb6Dx7C0cd2Do8
mRYl2rqK5G2bqOqc9qfNs/RPJ7wgLolKqd6ft7TAygIX64ZPEOjy997QjtpfHUejVW9FVzFRuOYs
ODfasWJlklmDT4Vxxk/G/sc24xWg+yu88qvO/Pko7/VYYifFoub8FE4+jEmPTMPvqp60IwHVJOHG
oAN7qxHjnKae9MKq5V8TCo0QP/DtZC/SXGVYyBh7+ng2WFA00NF2N14uwKpIbyR+exv+7afXA00g
axh24uTpIew1zueCjsCQhmBUFTjQSfe64TvuyzYuisSlnokLY+IDeJVsJ+BThuo5pwu38d7BW92p
U4CurkPjiQCJPosiBl5BuSdWS0DdQT6zryJnOVuqqfVDQQxALTRFb7aSykk0liFAtIaBcf04Bop5
h75yLdOPfEVLIse6oMdxABKkeXhGZarzJ1eZQMMx7zpL4Pr2HymvmjFArihHrUIio3AUma6NSw9P
+8awX0KEkvwsnXVMCBbmf6w9d5kjGuF5KvvmbPv/U3Tol71a3D09lwHWhoDlEajI22jIrd6kLvIf
gJvJP3K8V1/rdWLDIHIzxyN8UhifPAX3PCWBpQ800sC9QibUA6nBYTuWmgUVV+42XCvAQsJW7M1b
jokFiXOoGZ76Og4ZAAvPkdvINYtRWPnxuvnF49y1HqhNqQBb/p0rP0YijvDVcLt6GE42UatM5A60
LbHQzTskkPahKDJM1q7PaBzIOUmlYDAsWWJGvvNqEwURlmypNhuAuZpT7C5LxZAAeg2RzPALSbqR
ayYxwD0WEABR2RvX09MQaIv1wD7oFknbrIfW+GSuy6SstAcwPIJni1NkP6gpeMXeIQQHqDvttT2N
aiWUb3lpgIiShXUgDZ0aE6OohGsA2yB3NyyxJVFsitt6dWBWBepEsQ4ZzBDo4v68gz/xztFCq0L0
Xt2l60bFqGG3A0+/G6TGQoSo21k3hQknQmHBhd6qRzfoNn6pht9BXsAo5iYVe/7im9R7Fw8ZP30q
iueIxTN+9fMfGZyfHpO1mDlD98FZgdbL3BSK3CM+W++NC0ZJxZFEOfOp34j3XG4b5qefKh8oJ3bc
ECvKv0qeWAHy429aFIJ88RSTxltMfUy00yN9RZnRizO4oFbFlIhzpR951RxW1xmIa7RhMelvfbkP
Ot69DGkwsv/1EjEyzvdq8PmSncDXRbgjmS0xfTUW+YZnZA4N5kCplkc5yVLmHUkx3TffJER0B3Ua
ZU/0/4AxfyvkGBQW94ee8hIxihpzX6k9d1XNJmLquq3VM0duZs3iGTuWpwM20ivQsssJc3i7ekC5
JWxkD/VALScaGCp/7f/SfPeDYtsRK3vz8IKEnWOaw34Y7d0fwn8n/3kgktIr7Irlc7d12lsnqRaj
vGbsj/hSbzPGJliagLc2tHYLnY88SwxfR1s5zQ4pULIzidxEmLsiyF8/IFdnc7EsWk2X24QkyDsC
H+RMemiQ2ei/5GDQs4mnQ3MR7bQhhHx4CS+NrKxkkEoa5pVxtGYoYUkkBbKcDIig8UtnTF4cwtxB
TABBues0pvE5FCx8iZE606jL4OsrBLMZcBbudPj9o7cAbN+Exp0ZLp/SfsLRgxnZ6H/fkKr05ak0
s5Po6TmHgGnjpOxRkCBervOd+1pUs3za795WZvbCTPV9dplsNPaDbCC5QJJHc21Nlm7AmJyyYtKU
cDFsqLY3Y2U+m4ELyA5f7EQaBfXUtF8fbAkRr21CAPbUIH5z17lJBgNpRgwUbZu5f90Vgi4QhjSy
FRubAw3KwO9bwmXajfziVLPhVsM725bh+opuSbVe2kzgtkzPWKmzlaFHT3+X3K8WkE49368DXGd0
3AkFKwF9GUgmWd8OPmfTx90gN4PgV9eUMaCxxnW2nZapeOlDRz5yX8FqpPAVEqFJTHp52roIDRrm
7sVbxFNNb/VCffH9gbZnT8y9PJ5mO0u5vWdTSpHiaWHe9XcPsNDwQOdCZ9m6rJZ3bBom5viWrh1L
aLfTLERemee1Bg41WwHuoUhjtSg6wt7VxhulJGqtIgYCO0aCadXMDfUVOmqcitf5coVMUVpWgwmr
6VFZIf6aMmsMfJgJN1S4fI9W8rVXTmOsMN/6lP0Mb59vVq95an2NmIYSku44w0+jI4uXRmTDm5aN
wVp6UUQHc36aQc6SIPKUTDU7J9IxQiBfjneARWZ9r7AEFIUJIM1MgQStsy9DhkP7LfOlsQ0HRtCo
i4GnRis5YmVFVGpPrd4zTPPg4zcYVTLlNXBO+7Y8C5rqvSGXm3CYPCXwfm6H4eh6W8A6T5OQqBt0
AGZdxemu4ETAMLomWfo0o5o1GtQxOD4vsT2qb5a+ZjCSf+fTtgEKWOvLWMLKOLGSURfsKaUB
`protect end_protected

