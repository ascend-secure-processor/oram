

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T6PLQfq+buTQufAvaN8WB29DzT8c2gjL/f/L0dj1VeorOp+Gl9mRJcXEJQgFrWjpAdyA4O9/Wnoa
OTb7phkbQg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
brK5ahTIZ082Gl88ccmzW0muJP8Pafw/dLpacdqrmH1z91LCYIBEbPKIQw6E8gJvZbiHsT442U9W
qGsq3ixJ/6Qzt1RfiwCXTFK9hKA9GqplcVkchxn7ZeqBYQgoldMZHiT05dZ+2LgO4Yzs5U92Nm30
x+6oR0QAcI8b3VNuB6M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3NMuqk0UTGQPgzLSmiJRPObdLMgFO/ZgDL7vxxx8pEFHg9eInuibowejcoD/oZegSM7d8TpgUShD
G2pIo3g4wA4d5il7qz5wvbG3JWQ4LKnq0WEj0F6Ry/NL/ZWrBsP+HdvSdvSMbVfQkBfqn27Enn4+
No6gsZQxNcGR4ab7vN+V9OXq4Vc3ZbbkhOHUVerB7FuiPKwAqRLPaPPkmyrpF/guU/kg0d3OuRBM
HJIRzTegKS0bvBDbh6ajc6wBmM6++1hDdamk0PhJbCNPOgUc+fTx/fN5VhaJY4kMuC5s3u/BlWQA
HuDbD0q63tRa+UAFhY4CL1JxQUmUarom6+lYTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UFMxDEmVs6+P/+ConrhPlmqzQip98IuOEG4GGMZMPoCVix6bOWse61aw4O+z2BdEEdCLaj+B7VQo
V8aRKeXzQCi3H86jeq1nS+UgrTMfiULyfJ/6fAYve3IYbNeNTw2XQQSytFgvb9yWJKWDo3o6LUpC
L6J0XeqRYCwiZpnNhE0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hSN5Z2bXKb9T7e+2PIQMhfaoHZ76LX6JBX88xIV4xE/X0OFL6InZRGDIzi+ggI0MzxwwXye2apxj
GDbej369DrZI1Vr6hwfnEkwC27Ktqgt3kXnWSnWMgg+xNLNLnce5pYpgBDwQ/RRVvBuqzpA0ztjx
brgrL/bnAzTHDlB5/7uAqtW9DOW6MOqocbdwocA2/iPGlz6+rUXUa/4kpTfNTdL105uxhZj70a6W
0G/ZF5nbO6Tpc6q/JL2895l5oOlVdDarYO+obLGqdWMV93BSLRjDJly6jTYoSCAGm8KXn0FSzXU6
e1BF+MPo+KXXvI0CXZ66yqb2fPHG7DVrvFLdhQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
FS54bezHbHQdQeJ/HRBpnG/FMNXC1M5pZsNidJ5u1/LSrnBZSYkdcglP/ZOx0yfGaAiVvxnwcvkg
BZBAs67jCIdmp8I6QC7/Ve5BKXoHy7QN+h2wj12i1B2jvzWxsBlTyIMvksSWAcgdWoU7Uqj8Uvd/
1sVkIzX8YrVSgGJewwqsGQyL5wibF7EWhxNVhjed5/+loyNCGk0ndKUxTxHgfRnJzgLAk7veMPJa
InML9eyB9Txzykl0Q38I0rb+FL65ShlJraVClnZ7W7rI28nzs/RoY7OdROUYqcQFmBfiC+uLrdUs
T/iXJGMq7CzlUeupqSb9hDYhELnATMV1efsJNZhuwE1LXfpoajkiJee2pHrVEUfcNn5vsVhI2Gmd
EJdPask43reQSxK7F6klRuv7HWVA2JZbQGsbKtbhVS1x4zLAkLvJFJSUrkiEpSeISfgbDa9AayzC
OFLPpEh7Px2cBrbDtMsrlW6HjdlLEk1vr1SO2w7HtOEi3c2yR2ltRYYi+809hq5VF2tiYjAbd/Po
VWEK4kbC/yxpaqrqZC1A3hDbdHgIzXQTXmL5xOlcDBypM1LQ29EgA/My175ilHjmv+MmZCOfnNvP
sC+2hrMAMuWRB4u1exoirj6Ig/t7r0DH330LkodPuj+6+Cs5R9xg9Ylu76C5EMC3XFaKYWyViqt1
3jc32bwCzC8Fw8mrOsnhOLkY0MRc4XaU5FMMDSsvBGv72PALoSUOh+Kkaufn2x96Y6ksVC36xCl4
mCKHoqjJX63Po8mQCGep2V4l0kljnHqtgGZzROqcicialg63mAVV7yyfAViQUJy51zvYRFIyEoKS
1FPaDc+sDcCyNZhklhI2sZw6lnbarQCG8Ra4HLm4h99h5KrmTFPyj+T4r6e7FaPodh6AExYuzs8Q
0n6OEDfCjXmzgWKlxHTBeCFBWZtOLdgu904r67Lj8mf6xwV+QRvINkScWhnzSSYFJ8USUT6Vmnf4
l7HDAmmzBfwUsen+q9AbgvD7t4itDM8JOOJ1SvRhcIzDeamnRU2app9wmVwMO449RZJY28D1VJwV
jxSu2MMnja/HKzwALU41IGOo9jB6YYTerkApH0KTbiOtqoxrA4qOj9DAjaUp4+U4rUcz/4bb5S7a
iQznXAw3qDYx+AEUikZQVL22uDjjwa3aMbMP7FkiuzhJegeCevf5Rd5sY5ED5QKaYBy0c69EW5jH
K7sQx/3S2nSP92xaCRiYIawijJvoSKTzCGcAmdnYLBljL+3m5ZSti7LGjr9VEfC41dguWXBDI/ec
89mB6cegBIKmQwqpqbuS1vL7bUdefv/owE4aZc1wB4Gddb38ySvCM4DgS3yeCLSWkBZeWQ/8Tktv
1wIQiqUe5eczmO5ammM7KsK93wAKUpGKExm76mBfJbjtEJegP2xE4Y1v+ZIU6QHWGrTRL7MOju3a
gBPWPVScA6ZoVSyMnkQwUJr8qZ5HSKCqqGJ8CngR/sKnvNLudVCZZW+GV2jcfm4DBKnxJLVqSdlh
b6CbzAtqeptTl0Ucgl/Fk30cQ3H7tpOogL3sTRxZxM80eDRcL2Lz/ZIqVUknU2A0DlUkAbAkFb9K
EONxE4/4EDSrw7N/QFpQku9+FGP1m41Z7Wj2vOaWoq+6yOeX+djThVbzf6B69aIR4ieAMjoxNJdk
jq4fVms80YPC9+jFSVjwoG3WBWtC/TZAD/64RQ1dIIN0eLLXHtxHdVEZMDAovvSYTUaDe+arwiGA
E1sDrPd3oQkMvAPxKGpBpGFJ6WC/fBk17Q3xhd2D7j2wY+4S0i/zjsLugfL+eTKqh1oxBPrPDGnh
PcJpc3Whd9OyUBJaAAG+S4pPQG0WOS9zdt4Z5OcXsG9TstzyorCcxzYI/LfWPHuxTgUBOPWAVHTs
6HSuE+0g3GRmoy/cyyWSAaTSrDzLXNt5a0euY3KQYkwhdbmfUUrnpYXwWkwuH9L14i/w5jioJtdG
9gWmK8j1fw7Ugy4BkTm4Safcf4fC0lGghPtSdj15cB8EfZyFMHos88v0iUmpmHEUB0c5Q+XXp+QB
D8yG/zqBf7gNrff+95uJzsNyfKvTzV9td2MGtCBj9NpAquE0VrFNGG/+TKpN3EAZg2fvk5tvVPj5
UuwNlB3NwuPD9fvF1MjEjTcr1ui7Ku9+/sNm+1vVqTzwoS0JcmP0slP69ECEsDBQc5TjuDdZZN7b
0lG25tOC36ZwybeVLCBueIzsdfZwNBK/YsSu+HkOJT68DJ0vFfGkl9DqgZlTyJxc7/oho7fZN7qW
KuiWKtJIShl0W4yf/A4eWNhSf7uaLZDIMfeTfIcQH8P14tPAR8qD6ZnLc+iS6QjqFN37x7TfDIi1
zuz+9IC8wkNcsdTQ4n/yU8hdxX/SxOrbqxj7Do1wIFcB8UrI2zDuXbl2B/DTEuGe30SHhGL3g5Ai
xhJiwAw/bIi8TarYVe66AQaWPr/AsC//AfT86XF60Alr7wUcgonV9XMr9VL4M6BX+82WqM0S9osV
uQT/uedEGJiBTDqKpuQIClixsF/tmqGdur0/u3w5a6LXKq+EknZEr2A48btv9X9GvszVMo6wne2R
HBXy8FkrAC1iFf24aU6xssKGohpd++Gs5B2KQDvwfb0/+kdqdxSensyBaQ6QVg8IGr6gCHoWqQuP
qHOWF0PfQy+rQ0he9G8Fn0aZ6X9QWPVojaXfCLT2+aReq2HYc9lVEyIMx/W3iTQSGTox+XuHFgxI
Mu1XbV/+SzQ5D1mZ6Nmt6MKCNmOJ7+1MgmD7Npx0OUkzak++FEMo0Dphgtd84sQ7UzgV4jKbeRyI
exiKP92mL6h92K038sHyg+5P4DEQKgMMdzsh+GEbsa1p03ptUUYQfVLbHt2+loUtWX06v4HceDq+
BFYNUoq5mWpzzKTIgl3Rd5e+GFfpXksmV34VFOGuRf4cTM1NZGsB/xWw/y33ZOlM2O7aOveNnh2W
DmtoCwEWH1gzA2TMQAdEqNdkDyygulJnuA2mAwCTjfydSxWTMg2uBhfz0/xG6BTbk2/zNmB3HhR/
yt7LF9piFb5cv3dMSAG3bCRBl6Gqf6eDgnSlvSspUCuQjYKvVW6RBNX+Ae+NRYvrNZ+y3KLV1rwT
iSyTolmBmMLJrWz0JxiK9nHI+GRavv/bdQbxp3s8WgU8H5uVipYeNvpM73c8fB6LO49n5snmbU+k
SimzCK5vfyrOlMhz0WPquRhLWn70DDe1+2fH5qdMBYbMxkHPgQPgzHvNAVSVFU3yRTWVB051ucw4
xSvoNVCAFtisFGLqPo1fIX5Glhz7LIjrQ/JTscrFAqc5wANYRs36VlWgS2KYiDmZvENpBHsEV809
PgBxy/JWdhj23Kh9lZgT6c0CsdG0u67KOH7vUmaHFUQ/d+cYzZWmdcDYXBde9XNL5P5q11MYi98P
3kD/tL7I+XSCs3p3NRzCk2nv09UF5ghXRcQzb377ztwjKXzUrL4enviNLGhKR132iDTmC0fWp5Ia
xB7LONTtANxO9ZEN5oLAXnqG7y6xKGLmf3W9uPPcyRYFUEqx+7WdkR2J1D68dFJXhPS8QW/SbSyG
kOuFw7A5SRguYYMT1rIBK6YJaYGJ6qdBgW7b8pcPYKd+RY1/bObpux8VZCsjoBgEv7Tayv67Pafg
mzbof4A+GNXJNv86DANCzG1r+k9D3vNM98UC5fzd/OaGQHB5lW2Ee3HRh2EuCP8QJWyfC/KDpWjz
72F0y6b9Syz39f49l4njvQ13Mk3L0ZDQZURIXZ4+rGuTs6PjySV0LdKfKAuBIlH1nne3SUReCiHI
JLbN2wLhLHmlDo6pDr9+o1Rc5cdGVSqaqS0nyldSXKC7aKbMoWV0sJp9tHgPEbuS76r7nvJkgfu3
LbCI86tfbYpuOGXvU5i6zVa2/Uaxbq4VGINU2zrxQO9KGFqlYmDx5+DzAXxcSrkHsP7A3p3bJGBH
Z8QiThNZ2221BZVc+uq0RQA3Kk7rDY5iyKkqASbHpgoOojaYQowS22H01L6tZz2d00IAN+DqT/Ud
VqMAynpvqibNfA34T0lhq8ptpMI+kGxzg/pqHuzt21VLeGJBQk6NDX/xedIvikEEZzXVkBAI/NUS
tlgTKODWWmjgu0ABv+WMVhJy/wzjBvF13GWUH8j2FtX1+J8p5kL3eXyK/YW45YgwQfeKKmuEPcMH
bxqE4TO+KQUA+qc5v6BwOsHjAdLKLlQF+eg7A01wvEoemOxB+g4XnAQ3YjgkpydN6Nfblovsp0bs
O61NRrZSXfdiW2T7X92hBF8sMNgjjd42wADqQIka3hQ9biyQ/BVc48S/3MFnvwVgYKsfKKy0jP/S
IqvD/JJe2YNgYqGgW0uoVzEeG8vYtU8uC7F9qa38ZR55dUBTDW7RSWgKI//999orgf6SEuma9x3r
GieFGJqvJe3XppeC9LZzbIS9ck/qzYiXk9Jz26JIJ2Ht5c/gl4Qr/Z/TthvdbdGg09qlJOUS1+KY
V4Fa4GVMQHLeiybZYKqZHMSQEe7g0jZPd3F5yPLbF7Kn4Ehbjdk5wy3BsqINIfnM+1QZeuRVBEFe
kyuvII8kJDko2Xr+B4PR2lL6kOcVLU/eu3nSKjGMeISGUUkoe2nQ2pKR7qOPgwiMbdDZmKs2T2xE
OIVp4UzkvJeillEcqpkkSlDTHsTqM4WvctXJLcBanIYkqLdZGGwKorqhBVwsMIr3Oas4v9fJKBdZ
2gbr/N4s32wzQerqHG82Tj8g1dsUGGs0UXvbASyZN6kyOh4o/l7fHNbrRydhA29Qlg5RPuG+Ea8c
CeZuUMHuPiQ5UCQJmBusfUJp0PPIIvW7wC/0p1fgNDsqQLIWvpYufCbPKspQp4fd/uqPWsKD5NFJ
MSApvc6235nvmOk6/x29w20P0ZjkMtOO1yrVsPBBFsmUrLH2H2dhoqvMmmJIrzKzEL/5XHRtFlyd
nQVUr9aT0q2GOG0k5oPUycEUjnmLvMJLbAUHOo8iDx9w20Xn55uQjw8FES+Koj2IjHLEJBO2BtRA
0yaKx2QGGM4bIhjIX+ndVj01+udLCCcmXBUcpb/rE+LbaghnnyMoqopVLrdBKYd+yT/PgXCjoeEK
e13Sg0N5BG+WBlffTh+zyq8gMIhUYR+R+28wv1CMeM8dWMft5B/LvVtLfoJQd90Bkif+uo9XjbiA
W6ZXd9/ZWlGsnVTboYkeViWL0eCcSPV5uUFLnZK5cgznY6LOivo5WIw/JbsGsWyI/C6c5ZtpxOFZ
AY19Gk7xFcM8Q7XM4L5AgAj6uQ1JqfUzoI0GFPUSUED/F/6mjLeukEqybmFIiYAJzBFKgW4we5pF
2xKljmCTj0OGZQ8Q7PoO8EhUpB1adiEvMXyiZBO4VBFYv8eaxSEt0XW9KOeEjLmRlAgFMTpaMGTH
0AhETt2YkEhVIP82IjXw1D0D0bhJNDuplgPG66/AtOK4KV7dFPl3VPQrd4mqbkrWZTZvorJ/haHy
yErJDWbm7ASkmr6aVvrIeWF31RJW5e5SEgtxEJDFHAXHrQkmfK8QI8UmXhiocbGpsqMYDV8dem4k
IUfR9x6wJYjG7z6h7AUz5vlA6KwTIAO/WAg74cSgK0no0MiJkI64CxBIwnFLc6XVWnYcqfKaUON1
RwubOfU2pSvCVLRxB+p0JHRbwV9nehjPOhLiEE3hIRlR8ToQ0s1PIs/6nQwYE7fA2YMo6fXu5U31
glA6TdvhvBa2s9fhIBtW3YJlq9AZ3ICrYDq+WBz5wga8TaI4kZ6N5ft9zTAL9EHYFBf/G1V1tQVO
91CPo2CarZCwRM9NR717aP52A6DFQXdh9dpx8AvhWdgm0Awpnys47qiFucErH07J0HP641gsYyPt
D01Gbgq8jqPWYf1/EAwE2gyPvj8kkQgmZT/29lbdTFKBUYEXITtA4cphiMU8P6y1a7H93e4PFGje
g9gce22vwNTzwyU2q36QnUP47K7EvJCvI57kVMq744mmG6z4xKBkpC7Zdh+eNlkdbKUtONxEldZ5
XT/R21NNQI4c9lTRKhPE2yziibcxsjMo7oymZxhQ2TRfRbD8jkYCNenZfbMVNSxy3bFEFL0dfZBL
ZE4zr87N+P/c4sM5lDSnjw+rOTxswNSjrT8V5ID/FmepSx30aKX/+FivPm49QrmHo6GiRsWap1YI
ph5HwWSFBd2G2B8YdU6IexA750movtLgJySLu5H8qpFn93EkiGHTobCoXgCFwcxewbxEF4Okr3VB
Y790dN4/FY1MgGeCKFCnkPI3Qu7LGOcqZykUUNErnqkMEyzJXnio2aBCvdECAf2ZLK3EMkd5pbkJ
ctBwNPx7Fyfh8GLwQYuq8++0uw7LeXkJ5PsyiCXePXsnwEO14YJEjeBY/9ftTGcbpHydYgFXhHNL
D7NCIZxun1h+6/Hda0AuLQymDAHC5hofEFrVE0Qr6EFPE+0YeDrEXYR3qTX1xRjh4g6MqL52Wj04
ho3RkgPn7M8GcIIXZvTjPFDZ9XFHqATNjda6lyopm6IJwjPRpGZJQgYB1z34ae1M423UBrYVoW67
TqIrpCQGm7aRG59/HiYePTXkemFOpwVp36sbk9YwoN77xpvDOaGZec4WqAdBdLBHgIM4pdSG8DPU
4GojgbwI6a1U/6pVaWjhJvd848XFhuWFkWVDl+xcR0E58Sl2bv0QLTXyok9ppeoFXCij1qzaJHdz
Asw49ljEmffP6GL0AOsXveaPpHcAEz+FdnI1Rc2VBLmBZ3ZwoQt9EKDMkq2UdLJy0h+LNAIqMrmh
i2BYmwe+1sufTe6tFoTyZj2Qok3FBdOff0zTVYHKVDVWaJyfNju8FBWhv4LLttJ1eDLFFVsf99Uh
x+gVpv1e9x9fhcxOC0X/1slKYeCB3s5AfU3u9ScbNrcJ/IC3K0OHHAQgas5kgQfbUAlqw6tYXyJr
yxR4ywWndC6drM5R8/NAdH9r3gSLwl/dXWLaQiRRu3m6zj73ED7z+UgKXl3C6AqZ2ofZi59kdrCk
MkYWtGoJvqVIfYoa6WY4zOXqoG82qWF91wiOb0AGVeSmdobzNhVvJTCeYn8+8D9mFviKAz5wmS90
+7au5D85fZyKbv0=
`protect end_protected

