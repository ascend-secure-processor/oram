

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QThqPKBRcQM6ReHNSyBTL0WHypN/8+2ouX0AIlYyfTx9mWsRZ7a3/D54xJ91Mj8XTwfvnUK+YYWz
C/Rn50C7lA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f2VoagMbeaGX9is2SGnBkMtzzgfB3CSZYOHpJC8Ji/y21SA0XjJdXnSq3idfy5/lKkeQ8DMIa19T
9wQCEisqOJxN6nheLw8RABTn7fngwjMYeMDrfwN7H1Dwm96WADU4sAHHR8hvo6tMU5+IRJFjlq2v
aMIeAMAHVvR59d0MNqU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FVQdKVlLn5qPCMF8wXSauZEiaJ12pC7R0OPIFgTItVSn+07mCwYUMdGZVSQCmg5X2APGNy2432r4
m7jEqc/xabn3Wha34do2XSrZsXW37eVpZSlsXmsGnv0xCawvShHjIeRfLuzgPylZPYHba6apS5Cq
BUCF+YowW/WVCuljv02Vz3F5hdDjMNjo+aI84LgGEPuaIGvNuQvgOUdRUmBThOZwWHjrDmJdaUcE
dXfJ/epWVFQCvRdCPYUyy98wc8shFX4Ea+ObHvxy59Xun/z7Fykzd5f03KPheeogSKlYk552IkPq
d0CCuD7wwQP/7EY8vtwjQUY4YRVNLwsoBsbgGQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cqgRBzbiww1KQZDgiXRvTQhROovLKB68+aC4vUtWgUYKCWTuSqZ3E8XW49HyvytGMbbl3DqiUdDz
dq4JCVf2I9QiG/BrLlsKYANzwRn6rfT5rZdtBIsZheEMxknYwN2qwBp1wpBMubzUUXRSbZj00cQt
Wt/9hVs5t5J9PRw0wng=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
beCZXfYsgKeHPTUJpDoqwpUoFvg/t4K5oih7T/feG5pQUFRf5C/GdCiTqNyhqJAlol3c4RiZjac8
veYZUs1UgdQZiUv5/kx2v3CIUe8X0d9U9gvIPTFCT/o5zIEYz0Wap5mygcl+DjkYgQabQHFn21lp
YKRF+8q6ARAwvSEgDfqmRr363oYhAitrqSOGIlzKr18h+sudSOPX9hi+I17RuGyqNoZ2o8dt7fIZ
7NJxOjsTDJ4xPlMGOTl1QMx0yLDm3m9n/0/NdVzl0yN36GHMiEnP/jje1caMbwiRu6lQBdbTlQYL
njYNVDJNSgfBbJ1LQ8Lc5S3ZImCbriHMaEMBHA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24704)
`protect data_block
MQaY45BAMCGBwRe9py/XXAXzpnk2mpEmWml4vdi/ekggxbKZ4fzy7kFPUw2KMYiVceyfBbLEif2E
t0gp5hLiThpRauIXJc5ZLjwWChEg1zoiV6sUoSTCC5o5rdftKK4e1jnZUOMIMiKCBMCgaYnw87Mv
CWPEksG3slNlQmM0OXiz4s36YKARDarjebms1k0FIYeR4O6tbVjGMUFEmbUpK1M8C7w8h1C9EH0Z
E9S6yNyicGVVLQpZto6UJaPqpQcwrRTRxUCGzfJsO8Lt9gJ8SES3Pt7FYe3EoSWkoeUuQ3rnta+Z
N6U7mfaTgFTlXGJh325wpPRQeyQV4Q2lpTgJYUJD0awF+TqkigPaGAQC9y819441C5bc5wWqd1kV
dmU4tT/pBuXlhbRKCIG7h1saUyfqJYsNGRZu+OeG0nCNUm1J/qr66wnxbiq08ugU1iSHVKw/gCwJ
JXTQNi9tAt2Ftnc5C/EnBCXRQChmMN3b8auoTeMdpasXRH66AUOScqSIuEIPAuNKGvuwNyK1N8Je
bQuelJjzAXrfOJFy/s2REmt20Ouo2wQniq3d3dr8Qz29JwY2HaKWIXrda8zx5SPWoHEMr0fek9tg
BCKw9WO71UwmIixtxU4rnC75N8Izx1tZDdYFd1ysINi00NqIQaY2/QeJEE2nf1tXm55Dl34LdQiM
oPeYeTayw4fNpfh9UVOxMU+P9AznoBYbd/gB6kg3Wvela2m6jFhiYa/B7niaDR4ezkQVPO9oxX4A
NdROqOaq/fFUcG83JHjvxK9TZuZ/oh1928GiVbY2fhPOGUHBKUDWxJd2OzqSdB/JBIJLJt3gygk+
pJtIZql0SOWqufMkmv2PmoE26SFS5ZnAz3zTuaka9M0v4AYjNslRD97Ka5dxTNLcE4aX+OphMGbu
u+8xbAxQWwe9m0VoO1M9cOnmo8/TMMonorg17ghq2y96xwXkCTzUxM5Z5oTVohcHr0KROgy8L3W3
Go6Fv8GIdk9JPKMfjd18PaV1UGIDD0jPodCHmx0ASG/T0Gq61aKHFJhv+BOnf0QrV80kd6DeA5RN
vI6BwUiEEyT/wqiUfIhtKs5gIQo8pbw+W+vfJsMdZku1EPFBJdlOq54Idk98HdPiuVQ78SuaqzvW
x5+gzLZxujcF6D1Tk5pM3xjTvIAsBZQvOXSuwUY+W8ZExlaxMDf7uNIoj6v2QWsXndzZtsGxB3/Y
1BaD2qK5cKoNfXIbrI346vps7f+NQnQAPPtR/aQkxCrae5Q+H64l9gAeyHAmLlGvbnPjnncex2jk
DjdXR9IVwCEa6j5wvWHGEYlZIgslAonqONDMBsHTkH8K4OIijgOI8mE7SVLfJ69OI76pkLZsBgpJ
UHi+I1hfPvO9kLUdN1kvSf5p+6kcGu7dvmJNwv59CJO7cobyUKRORCay373rKHr9q7cnblIt7ijZ
UIDBnO4igymSIfduwv+7u6r0Q+RenSNFt+ncNzWzmndPTA4kSVcYSEHCxV95dxTjQiFyvuqU2lCr
u8hM/SDknt3DnHSmGPJE0D+g2QBeSLIwlO3wT8Nw7tw/Mg2Tx+F6SI4WLo6GFHg/iFHcNBI93UFZ
R9KrG9h8qx8ScrM+TKA/ViIwdGBebKBvq6TFSydS9DwM8neKIBAuKdf9YkCLXxhVUh/S0l0uHZ+g
EVUkeK0IrfMe5rjxaSfKDm5Em8CGaz/s2wur0LdRHrQr4IumFEiLKqTMZPSVgpQmiQoAQHg3527p
oPLC/4ZR3soQ3jIx8HrwYgyaVAN8gv70/bLngJ/suxbmcDSJR5vguJrw9ycuL+ogqbY1uTciLrpC
+g8xdWev5kZh51QHU5TTFwptKjOWHQ1mL+w36+FZltS/dDDSgAPi8g/NNRgJh+nd5ONMff9fMYkq
hlxerDpLi07O7EI170J7w0GdDgnb1aTOa4+U8m7CHDsytbkfOTTltiy0sqQlD+0NaS3uH9w035fP
P7UExvLK5GYtV6bXjj40ensLT4dAGf/PE3DLtkk5xw1JXXDrhudYttXagZAwr8MXyJ/tSpUBUEJv
tmD7qDTVHbu/wp36/0uSHrETmskZaeGCPwCU6DR69CTCxfa2VWUUHRJKzS7R53NxO7DReK18rJp5
wvfxn+NajIMvvPr7O2im/bvaE03HI5dTxFF60Y6wbug3WcF8EoBWdMsCm0V/AHNZKQyw1NoYv9qo
IST2g3MW8oVdKu6iEjM87jUn0FwMe9nL1X+lyKAjKy/rjNZheJVLawHSbpv+ADQkEIg+nLk78n4n
wt9R5Up6iwViu137kdbOUZPQrCTj4wQjij/5JlBCaxS6IRfdPKUe6ri9Op9nstV99qnIM6dZoxKj
TQ++5f0+7ozVHPB5FVpdxVqYUgdUWCAjBs/8IY79eQ+9Qrsa91fOWLed953erQWGuuYeTThxz9Df
EGk6ansmfgIpbBIzPlu49EytzvbgLsTs4mpXXtpXkDFYMdy1dZcA1QaMmlb41PTUUlHZA18ziKUU
tr1TJgBqOXnoo63vXmwg5h7e1Md7m7BCyEMnyc4wIPEeClnTsgdx6qGMx35PyUZCbjPdtafQCVgM
DTlU+Vh0x2tAg0lFVehUDvzby7vZipgPZqXOmgGx7d4XdtRhM3hRrGfx1u0SMhsWuwW3i4/7I8d1
7xR72g8l0cHCEKE+H+zdwwM7MJdW9C8XjGBYvAmc0RmLF71/aLsC9gMJIQvkCEg/XQJ/dam5yWYO
g/fMLM38sGOaHYxwAxepoEQha0jNnxbMcLarQZ8mwzTFZ4HX/vCxSBFG4d5eb3eQfLW7HtR5asjR
6tjNhgMKqsKRRmbIWSVt2/Q/ujK6rYilaZnFK7zM0W2KhVsc7lRsuD/GaUULSxc516A2NMx+nEVE
uDnPPNvbKRbayX1UO1FA8lMZIigsqWOk9ditWRGO7dEU1xbvrDM0tbAYX24fkzuXbSMYBf1iz9L7
xjt3PPkpOiPLAfkbDkq7aanSUZcvcb1mB2/qR3Z8+F5+nCRcomo+LxMbBvRVd6uIU43MNPkSXaXw
1si+dL8Er5yXwQFoQfg+XrPkQsR2NIjp/1MTBReaSHZ0TXpIGjwQ8Ja5M8lcolw3Qq45vXqm8yAV
RZ2bpUvx8Jn8hnUHBdG09V8Q99SE7726gE42iDJaXjK5ggbdPjlCjiWI4zzDKA+X2pWkD+dU/M5U
RkqpJNHm0vyisB9Xn98F/dfScokcRGo3W/gyIiOVplqsgxHJ2pOZBlzn/sByXOWZGsa6d5uGWlvH
HtJCHXZcm2sWtENVcRu/rRbBALMKSutvgs9wnGUPtB5cSKtQgVIRhOx3C2G70+ApjN8pyoS4lXv9
BrYi1WHL0bB+22YQ3VhNcMRoEpOrQfSl4h6XZkX0PXdpWNtgsL3x97IxPxtNpBAFMQ38utxHPc5x
dzTEuEEy1s1TWMZebROIuA7I/29h9q+9rk4EZRgqsSnvqBEmgQBWCpFGxRiHecpBAOFq1xd3wXj6
9bA0IGtYC/7/CSubcsaOS6A2uqg3kASJ6R+NyYj+Z8GFu/LwPstiG0sGe4aV9wMRjCiqdss4BhDT
XFsDvejStw4BobHxp1TWaM3iXI5d7US5+WhGoVbGxeyp5uk+I39Wu/oiEWBChALQs9fazIDsju2T
FPmyIKICeIe1qsGd6OroHAKCe7U1OkG3e8mDoNQBnMjsEnYRLh5CGWGUMLDAH8kXQ3xtzFWikdU1
IXhNLy7iXMjuJrkKW92EwZ8/vIXxAU4axGbmE6fj+a2bs4LqUSh7rKxfsSoY/fiJueql19ercnUj
BaLi5bDo1wDqu2BW3avsvPrcKtwjfIJX/ylk7N0539qqG8/G5GfbHtVbwG3P7wAYM3HD/YbxuW0m
hbyxliME0THhkVmpDFoVwGnya1XO5oFo1Lgj64EBrBahcKX17UzNCJ3WDheqYxshT/hxmRiAmWEN
jcS56MTtMQcHVTaRQONCkszGM84vpozTS5QBbeEt6D1KVuzXdkCJjAc6bJLbL9tDHoNDX76pAL5U
Yndp4YgFA5Ew8wIUoyY7lSjYOwJS3TpoAkj/lOiRm2YOz5DAt4jnHvFn5Kcqy82Qg7iUPW2hwi7r
wY3UsZZ25o2r4omNxbN3pMQfsZu3Ux5nHdrwLKN0z2kmx+D24C7lGGbVop0CfegRj7mqsT5YwTIE
AeDJ2UnEdzZQBuDr342fMk03C2I+RnxA/VztdgSeKg2j+Udv1fMiQ0NbpWamm+w+EkqdAgBL4mN1
7jex8QWpPZBZqUX41bKV/apyVD2ipySJs7IHyMtid7f2fY5gcyTBx5QR+/Na0G1/XCSFV0lTd4+H
DjfYbz2sUTvEUVi990Y5smR9NX7ToPRXDo0TOcIaVa4TY0P1ifGRfOatgR5+t3Pg5vRGPybtP138
9uP7Ao3rY9bb2mqOmCn7tJy64jDcs0LpTpwbEKP953edWk5sOLKQp3uIShQ3NvXq6hd0cZovI6aG
isk5NfjaZ6+9M4/qxbPuZQQQIj7W3TLhfGnbZ1yDAcRbvYtwt4sud202IdQc+HhZl5zAlB5yPz4A
RCpE+nBGjo83p09IpdCHcSt7d5uEVwYwc4Vs+tXlC1znwhufkBb39bNxl6LBKoeL+pTxG+1GxJTF
D6vqA/rqYr6Y23x4NKgZA5sfyRf85zw8DIa8knw5geW7iNzCUCElWeOrDJk0Xb/FRBNmbzqKX+v6
nEvY+JpecmrokDujw818xLb6G8IKodWI+dmLdoyWkZyoswOpTWpaiz11cPSxB+rwnMMC8bS7JW3b
nzCojtiuLLkmTrqvoCq5L/KFdik75ZioFvuH+d/wCQwGT4ApZ/PWrOhEVZNTaUj40q7veidGscP7
qiGpkT2uHse97F1SqOgAxa7DNHz3elkIBz+nGLf4J6FiZwvavwnaM+g87bOlFhL7TPL5rPkJyQEE
fiH7KcBYjLvV0Cu59Lih4YtfvMROB6mN+sXz9OTn95D015Ern7UBV/fZTLpXYLXfblng0/QWq7Vl
mE/P+E+cKhkbn08MzepokHixOxtLe5XGijkb67MX60DldIleGbmjwnHaDrglQOQwLhQEsq0yHWEU
Imo8h2EfyodCF5K1n02DMDXOjpQSj0qu1C48Iv2Zgk+v2A9AMLdpUiay1cWsy3CbyN6ARpVF/oAG
Dz3gXLKi2KNbJ/PooJRsKxbDr87S9LZsztPq9DYbld9mmOVu3PAdv6w0oC4yfhngNxisAW2IFQri
KIElZ8dHQOptCuLnUP4qTYwKV2/Cz0cqtbGRrjgM++pAQmT11kdXc9PHXR1CjqX3sM1k6WWcXxcn
27Q66r2ZwRTAirw9htPELGzWY+nYIUwylZw+Er+I7SA4sVn1gDS47yNgRLOsMEzUUiON3XqD4ar/
DfpT4RJYXieeHmKVSQ3nwtn4AQTn98Aud2xGp6bVHUDnDSY7xxeH2N1wTgPcg1Hkg3IKfr6oTpme
DtBsaba6xjQr9EpzJPIctwlwIauT+7AeMmhiO7yDNL76hL+s90oNMNh2xh3/YDOGKedVsT85/VW6
y+FwrFaEOUP0nkpK33ZsucFBSrHWcDb4pyOylKg39gOIg48r8l89K5bJRDk9cmqgK9jZHHuBR2+C
lR9u4uNOI0jUS7f5rvK6kaoK9VSqHQLnKVTM7vx4GmhQ2T+8fqTSEjP71hV9C3tbOuXE4WSHsu90
m7J7iW9DsQF3uUX0omznhCDfKST7XBgPG03TqxkNgoaMUV2bxZq2ylQ0dHWuhFGuP8T/Rx9mRLnB
c6M2L7rXEbZhBYNHea0ImQVytFOfi52CXGQaE8rHy5gvXf2YlbDnDq+Isb6TiL9R2V2Lefiql4RB
jx9MnK6jCnQTZQv2Tstbgcb4z9+brURzGmrwhCvHIh7OZn5IHI1OX+CDWwc7WoG5o26zYW1AxKPN
aL4MkeK6YSm0xFIYAzg9zf8Sys3dbemROY3RlqHk/XUAI3geMCey7vrLrt7FTZwJ4VDKWbGkE9uR
51VFVOHppgDVA+SvuoNOM28byJs36mo8QWWYUlaruZaVToV9IOmHFM+8Txpyl6+tBwunbjvmuYVU
388GjoEVlNOOVxgsrDR8d2+rrAIkLPwzPbf4fX6wHDqCJoHM/vAo3VFSw5nSOhMCvmmWDcDNbQgJ
vlLc2Ru1ZXcmVnrLytgNqUGdwbh4vhpVaNGHXztUp8XMzVwnE8e8/xbmVm3VNEolDqRk7OkQg0GV
n6EvP5s2kDRcScqNjAuCWkhdbo/xrvgFKCltfxs6WAmzLb9xHOx1aPbAoRcXmkx8gFHTH+rVo8PE
iOCKzKu1xANy+NQOA2Lp3TCwJkXZZoR60WbhsQ8UwvT9HFlaDKE1d0l4MuPtssuVKrmt+IwTnR93
oUVDWlRikiA8GTdYdsaF/0KWBaB603lCeniGxt4y65vA0T6bjloWY5bExFwWx4W1aizw4uax0BPx
AOkUsML6vYaqvXwF/EO4llqvAEgDQaxMR+h5rK+fj1UYEM2WTEf6RLisEUWvgwYtDtNURGvOSuwJ
zfiCWieOuwu9q+SrEGGIv/MMhKxmdH0jN4L0yarbPT4om7yfWdTjptoJPzq39C6xKSmROA73igio
0uqGgwDkIRv+B0clPT3vnCsc0tpPeqUmhpc24E7TXIdlYodWm6iqZ1yymqDL/DDvY8ug2mTOSGHO
g5k8tOJIKx7gy5BsA1bSlPog1F5bmoGP4MdSklYpyyaEFacRyk0kzrh8FrI/2PU5uBroTT+dhbet
2W7NTrVxpD2Qew7XIe8g9gYiXdIkSMdjKV1oDsGWWIDyNaxYZENoFcR8lmlu9Rb9xcvzwHx4roMr
bowwZ4h9G3dbHnnvKUf6PCtIzkQim5W+bgD0pGHQxUAr326T7Qt81DLaX20pLul7zantU3w2rcPw
gh4pZT4rvgvQYJS4EPULn1P6VQPpRreISvL5DWvrapscsIeYdCFWD3BVT6RY9AqC68iMgyuONwBB
UaoHrnEXC4vL/lHHSlMhe0V7wqg5ozjb35btP2DN2vNMTxpR85Z2c4mQYbPQfSjbmITWH6eG8an2
ITZ265DIWXhx/xHzLMCfPerrh6wsF7ylQ/cm5rPyeJC2dFwRjTCZLnCsLlo+fedjQNutSwLVakfA
nF/iBAh174gFqpf29JYDg8k4MmNvp04nSClbOR36ydw+b0yUdY/IP2Una/B5F24w5UIHW/8oIJZB
2I70s357y+gSmR3kFdQscZeLGGeIRrKA8+OJV+fCFoX9hq8l1DF14aVJ50TSUzFUqXcsn1pGgn+x
4LSuZGxfdAI1lgBdu0HfNRP06OYSMo7x6YdRE8sM3o4MUL4v8KKADWOoGoiIU1CK/fMuxuiUBex2
lYv2sGrcd2M5Kl5mfIMp7Gj1C5VYsn33YRQlKSVTK+7xZClXKRijMMUhNM2fMl9ZaLT+zBZU9Gf+
0D1kFf3EE+vRdxC3ql9jX//N63woMOfuFObmsgERiQk+5RcDF5oZQHV1wXMQW4eniNbT3tkdUfDn
AbPdWNz4vvrxRJ+r6Z/mp5IaUsX3XG2QobcBqM2dcQP4VptMXYnhFIwu78WkY3NKoWEyEzpiY+9k
2tpQ+pm+c0UAtyoGvmC80adPaHzEYwtJhPKmdQ8cESmhvqFPBm7yTms3gsmB9hFSRfUaYBfTUe3I
avA72YH4qr8fyDgcsoHM+4qRaRrzSuBto3Gy2riA+P6+LfqbFI8jVSwAaIpiadPvjsmnUqXNmspp
XOYXsRFKPMGMPr1SEHHzrGUYuBdBOXbZHcQRzRIpO1Ej9iL5DpVMbaIqJLR69wljBx6pqUGHY0kF
bgoXPR8Ps5emAXDqFdJ5VxDcTpAw2w2ZPfBc+lqEY01B6bad9Qcri5H6D4uS2vnqTYluoNAkEwuK
FJenL0dgJgSe8Ujies9Y3fePOzfvSkdyFv7ouCZJSHcan7RWxx2zuBoPus0Djhf7rtCqQdgXWB6T
r4le+tHRZmD57j7fj/clbyBakuocmpQgL7Oo8jhHHXGPL3msF1UjjQNt3PrgpFOjTZDt2T39LbMu
zYHrCItxAn/AoL4uykyxqCVkN6mCDNzjXgha/GYCV65ZSHJV6pGlxISF3JlJ5tCY/t4+HQiBHze6
bqOQlw12HUGRCQQyJRHhKD0Tf9epoz8GSV4piCxIualuixm8pwwqBLypsrwG5t8MAP1Rh7iG7FEk
0ST6aQ7oOKUaJ9SAhBcXEuQbnX/w2JmId9o1Aun1ieamKgaKQ5A4no+SGvBIvkGDF6RMrviJ+Mhm
CUSLV+URx9PsBSjmoxmQibkJjsCrJxvXay1RjgJos/jV2PU1aNskenMCWexkUaXAiwIPCRWRpX47
W0UmS5GiUPNhwNIWdKNtSMv+gPCQ0nFuacs40aRw9g1lk/4k7euU/4SpIoZYw4nwhRKe7t/t0Z4j
cmSXRiIx3ZIlIhMxJzbr9O2UgvclgNadEI+UMJJ1UZxZU6oTlKZOCoITfsH+SjmfOsMEmslTbEDX
Tf/Uos9ZmmkgGaMVA+INLaTP8mLs6lTN85mokE8QWHrm5vl/OM20s9t3HRVPnjLBYNvvqGtzjcj5
hLr+oEgeRp8h+MmdyesKUKvzW4mjQuSMKpP26l0eA4tak5OFen54hsemjJk0mB2EDnO0DrHmuqSd
D2idI+reKMNR8AzyRZofy0TAyj/iiKWKA5pWWvkyef4HOgMdA4G4s63Sap3hLzX84aOladrplAcd
x9PGFsCrqTOk6Pt7/EIwnLgx4ivLAKe8Jxk+IbtSRyD3Qlefxr6UyKC3Rs3UrZ1dPJ4USScL1A6h
bzYIpP8mCPhH4QPr1A7fltuAoPW/YmRPMhQ/dwuwMnA6oSVxhPN1OMp/lr0FF/BPn1VSyvZxLkOh
AiI0ko/soAJC12XY+rDyYDVJiWN94ASnvf1I1V+aSrXSQ3RUt5Qn/D4PxQ+jmjYEdoTd5GKKpV7s
xe3JpFncna12JnjDWc4Mw3/cdCLA+MUKJU7e0U5B/tAj1EoyO6C9bFwiqtbMZTpdgjgJzOC2VpQ2
FG7oxkNjvXNd1+AhIfcSOqtZxYuu5XOG9oj2YJY6AS5b5LN6Re4/F+0c9ri9+bi3C9GCnH4qUDv4
EzqH8U3exQmbpshAUL5EhuAoQB+/cPzIIXqXTY1Cacc4c/QQIK2q/rlTWFTtVgQ7zQGaCR44aRG5
ceK7Nr/qpP/OmqiLztbX+iEHlfudGmtN7B/70rrpEmDC9fMvx/M4ogcHzZHZnsHqTI133cg2+WJb
6fzq16SYQSK6PdPfnQ/8+j7GuqbDwz+Mxp8ISk/B4iaxbTqC+dqsdPlUZG0nMHqxLpGQMx84kKhu
LpsVoo15YcKb7v+ATmCHBrJO1RkIsmmDsfd+5i0wu3ilkAbPT6gwbCZPPQ+OknmEYgWYB44t2cvE
QoammwO7iksGfUflKCp1JtNjS/HX2TZCVyaVGZiqOXcH5x/vv6gSaf1LPulcDe1GaLS5WaqszOVv
TpYwEvD9v6+24GLr6yrUsSK/Kt0RS79X90bS5xoehxtl9bSVM4hZI3klOQ8W6JO2Z0rPMk+wE4XW
er2A1AUgS2bk4LFkHIYV1NpafguV3Ylf5yNB+7VfhJ+PR0VZaogifFggtXuTJYWDzzKMQPd+xg49
rxnDnNxS5aBlvS8r+fArYp9JI8X9RzdWI2Mmz0lTY0euIGfpwvaDqwVrBzcKy2t7JYik1543of1s
Q8m6fh2eKbzTkLIWl9/YVEZINUgHhgQCG3EIzPl7jKOa++QaR+GSxJF8XloaJBODTkuFZX4C4jRj
cr+g3otnPOdt8wiW11Ijnl8Qn6WtdDuk8i86fy78gx0I1cpyM47uTL6Je7S0A1l5kkSbFarKa+2d
WvHkw3nmxf/lF11L8r2w8/CKdrac/jZzuor8immuLlSJYDPwo/QTSNhBB+6VDV63POB29cxALQVc
Wz3MRBplfDty364P6zaYY+EjEoBQscPqiv2OPWTLdgdeGT5Ieo2ZoMuP259HS7RH8UETCix9SKrp
BD+WLT0TffKuXlIpGSbtd/lauNpirNFVNRcfpGgcMJc6qIxZm4ZA1GbP35S1ZOq3tNnNtrulsYWG
bHeiuNrzHZ2K/nPzjr3qkGi3L/AdqOOs88yFwfWs4sph/O4yUbvCVfOFZX+XWXy7Vh5wQr0yOEKP
vtCrSnBPN1z5h9jFF/zL1WIZCmCKCdYJWmak6Z1K1LJNWDlJgDLK0IbhegOcvbPLMMYi8hjrrpCT
67+fPTstv8KlkpI6LZXDAX5VzJ3mExSgqOyPSHseCptC4E7f/EXV44H5lvfBFxKmm74BbKlA+ZNg
iVLI/QCqltbWmaIrUGe08rVSrAjiSPwBBJGiAyYEBw9MicCrjxsXEcYhkdw/1QGEoEJV6IUHwu4d
AF5sAjzTbN1cW32ZtA5ARZn1QQx0GGNHyt5YUqlbuQkkkiaKmkJQiowwa/zagN8arOtaPVQlg8sl
lThng3TOdUgwtVv3lrhg28HZiOJ9+hNyK+aZOIOCubGoPHa7LqthSEnKh0KKRMMr85zxrStmly7/
32YXVFxkobw8RZVx1vN7oPVmV/idhoF3ABXrdXabodiBjPK3QaoZs1wK1kGANq6n8PbcpZNBjiqh
aTIRkmG1cY5FvWJsmXkae+K4WuNvbH3r3AdODXziC1cALRCoXit3UOwB4vxMkqfkPFlDHWFhj2Jn
Bc34lNClzczKpx0jqDH3kbSOlXwcdo0u/1mZxk0hxgc0djON6To/Th9fJGSjUlFMqMl0TXLdp7Q1
reHo6ehKYPso6FTlkWOIeDng7LuR4oKWNqKrjqxitglHzlhbykTdDlDnfk97UrsifnP59pEs0nF0
TMYYQmH4Rwf3BctIvxrRALNaxxspKrAjo/nZGv2EFevE0JiO2AF/RblrmQ382Q0ZKmX6xbmbeCtX
obLMhzcDTVtt3aeJ1ojTLKZmBg3W+X8A/ctyESj0Hb4zNIJj48NCLSQF/WXQLRzvbXoxjOH74rnG
nl7yQBj7XFurd+XkgG+jq4whv+B4zQtQbTiE+u9m/RyudjZj+A5ZXTdwUYFmKr1BYX4ITVePqZzn
CNmB3zWuS75BW9eHT1Zl+NzfmJWHhwdEjzbmkXyZNXwosOkDe3Gsg/ylTGKABudQ3EqjuPGjkGcZ
QJ/TM6kiHHMUaljONJ8IdFnToga6CijFsCGVFxIV71KRRE0uK/rGfWUxYkntEQKSz7yi+lGlRDGA
buFfflVorkmO+tqaLibdx0ZmuzZeNhDm+JEX7vh4gn5GG7Ivpbb4cV3Z79owB++h25zjx3jM3vz9
rXaie7E8GvPBzsaBuSrS1fxnwsE2IzK9W1e4NHeR/qw3LJwrQWSgp2B8d5Dw7px+K6goSkwKOjXm
6EFg8jRyeM6Abl9mZYM213k+fuoiz4CnbqQf9P7AbI5s+Ea3MTJfhj6JVsR9JmWDo1nBcUNhbv3k
/JM7V4MgNQpKBm2C9tkGOxtNXxQ+Y/LdZBEEgcHam3bLr1ePwlmyxcLjEDlFM2o65nJxwYxpJnND
T6KE7cJ5f+8TFiwQg9u8VKQqZinZKBoVGU+C/SEbBWTFgddKh92LgWrRrpdtBJQ2TAFd8wRuvsym
nSgTaogtDye1INB8fEQSufiIZ6fJ1zSgCbqwX4Lu2CJgdK6zmVp7NMvAWkUr1wRYzV90mFYk151B
hHWytg6I7b27KfLjVhPOstBS4LI1Q8do/vuRfBPirKzYrBKTmgFQsX+e8Zf2/24kKvLqSwOLXZCq
QFnxM3VOSH4AQJMc9G7La2NUbqfPz2w6MVDL90tZF9XvZvMZnUAatzL6BQegciifnTCu5v11Hhba
PxJZWPOnrh/S5KmjeD4mX6ByrsdHSH046RZ1VB4hWIp5SL/rFpyV684l/Y3MYCBCR1EzJyzmOisc
yX096OtzpdgWyELlwAEsiwhYxC220ul7/eaA9dCnE3PVzhSb/u9pW5gsxctAWZl9LI5AFOs4zT6J
rfBI64rmCCiBbgFqluC2Qp+C/y8hHHOw8CPYEHky4G+hYGhKe3DYbtft2vGpuM7s8BVEtgHuU9e+
LbfTvH1MRFQQlBBtN2SR/gZ8mr4xxwb5sN6xa3lwMx1SFAjwSIqCsVXAomjmCHyBpP2s4szhL5el
kYiXKko6jevoGsbrSL02SP88wlmJCdJzuIeTybwoutu+7KDoBvPHU3O+pk3q5HVV/+ZdN8t0a0D3
4rp2SMzTY0g+KtvUmB7lr8kPF0K/1fZyqK72v6jR0zA7ljyxf61SJ9ouA9RYtlHuUZ8PK6YeP3TF
ZkSpHiVoEln1o54ELTE3auTnFobI5QswfRUhLTgAaTeWPm7/BINzSM9/fu2tjveWJtlx9OyCbA1L
M2+FVFHa4OgHvmNX+xB3bHEP1zhHWgTkmuVTOPJrBgcTUEk0OD/WLq6hPKrH0SUPvBRB/TmdkMsk
z8PEojQp3u0KzI4XUPbiAQQUuFkH82qAnHkDYV0RLoNvPCZVb7hydsq1YZJwBTtATKiXKFqIEEb8
K0jCqZZHRo758EbB5oT8zL12aDDCrgj5JuentGTSVD24X9w0WOp99jMSI/dBIw3eo91JdYyjv1mO
PM7YPhFCsLE5B4s08uKP4bwzoyi90cYqfIYexoAvz/XTeZ8NilgTZWkCbPJIEnz9Lbd7Qcc8LL8Y
r13lcHy1lCPDSakfCfmbjGwW4ZMh3WrUkxWLVDytyyI/kjfhBt3DAolJcmsCJk8i2k4h76ttGQdY
jo5/oV2o8nVYSDaCVn8nTU1xs40eNEsUfY2F7dUDBtvVH0nc/+9HSkRh7Z0tUQOyYby9AIFA/PCu
zFQjvQt7L3TwxCXxKBmGDM7ecGwxrrxRzWyPxL7GB75oB3/+PlzT8rwXv5r+g1vf5EK2K9e7Omjw
BTCyA6D7F6i2Nj38nXwgkmivprGr+oxNYAGQgIvy5BH35nf1QSWwFSEriHco1UhgiGrEl+T4Oyue
s1mknFCoWLPa+jME6c7Vxop6scgmW/7hBTLox4YMlIoqNCT5Nc/xgNwiRKG/wA8de62wVVIBJOmu
UcuKt+oMaJPHGnZpbmuHd8/I+ylKOKSX+vqe48VZYmabIRTtwMT3udoD3Dw/m9XMWman+WWJhDvr
pBOOlWJvrl0cqUsfDdjbTmx7Y5ecARLIsdltNVV/exOAMRjHZFBeEhnYqTCTLBDEyRERdSnOadL3
UIeJNGIq9qfp+xJFUvZ/Eg8KBY9Sar/JDt+HGhS2ouL2cc0gb+UXcV6wxkEer+Tlooe7kOi8N78B
+BJ/tiHZJX/z/QTSJitO6aDNYTpUZDHwM2nNFDO2KJIKpvnvAxtbacknJ1eWB0gBDAs4RA3ixtn7
V7nE9Kt/T8wTO1Ro1+8JZ8svsCGmQRTbD1HCi/+G2FolnIcBvV03TetKVQpW/lS9s/WTNMFuRL+z
mErm/jfU0nEdrv3lU3RrcclDzRIr2MzGRBHKhuxEMqjPRsmm6Ga++3G0qcx7ckfCZPSrsQc+8d69
iJjurCfG8P5zl/2t56t38t6TPplmdoHanKRVvI2FLGX3nE5uhu+nSnwF1bJHv8NwkmHM9dsAol63
ZXv/CkpneBb72W6dcWjmi9EdMAJv4B04Nz+7TgeQ7hoxqDPU3UoxiV7XVSnQaK/Nwe3+LWpxwm8n
qm0neFqBcfMwTxsO53In0BLS+HFZ5yhpLP2K8K094pZ+b0FhLddzhxJVahZQoht7BZzQpkneU56I
UBA0Jp1gmhwhf0CtVCBAHG5rnfZsEN5JP5aNd2/9Pz/Ws/9GJtD6MEWIJyE2wgE5zklDP0Reg6SM
XdwQyjH/u96uK+C2/G6GClwzocqPtQ/eMGFJ+h5psTZtmUC6nDe/zedhyUn399XdfT2P3AQQykRI
V0yNkSsswfv6k6IEhjiBEcfU9vD4+ngSVpUorZku4fAwVchzEgerdZZk/ElJBkU92bnBh3e7BbZu
fXBMIY+8c9r1IavTKsoN8+JTVLTdEdEwJDZvJPwbn9i5Wz+30Rpft+o4BDAX3vx+NqmrGQFDRHQr
NgO+crb+7UQJj/vp03SOSsvJiQFdHUq5toSNwbqU0FBQ8ZbsFQbySViK9yfuKKxVg08X4yRNLxRY
Ssv83MGxDpHpRxmbvttBHfnZY4TVXE4ecTL0uhIkFbBvD8QYNZI/oc/FLmqjpBiAZdnS4KKIFIS5
loW3cb9XNG9OQ9YHYmuYZ2vqPprKVNx+8KdwEvC2YaWkmqCp2JOik61GdoaB1E+97nDIDwh3tZnC
US+062HRbOfXJ/2kdfFdar6ThQ490ufTqRwc5tu3IUL+SEpt48JLyDgsQyzWEbmOX9TQCiSHx2hU
/xzk32FEZwkcUUPIzrk3G7H20aB5pc0pfUuEKOSxYcj540PBfRiQROwmCJtJexaiQbkUC/qrFETk
6aBnjWGK5xtZrRAUw+YBEE2rpHhouIvtgbq0+lForb7RKS5JlTmmSoTjlGpTcFgtTvJvyES+5sKF
zTxHwXs0BycBRRPyPM9kk/2OQAeSb82Ggg5i523ZhFGGroGAZiUik/z+oXXlG0IOjpcTX7wjKtWz
n9h69oZmXBhUegqkIaD/t4bwC+UKUBRL+Moh75XSGd96UE5KXbvyjfTrS4pngcGmRSydoiMwhLlD
Vd1LF4g2MvB/ih/YkYDjzmD6fQ5nT2BPXG0szIaWzm44Ps87PfxMGEAJ+vdrWvBk68DMjoYMoKJn
KZPUyxBRCOxRGyRHBZTCmHoW2wp3poLSNpqSURZqtZdfx3phVRV71xzSYxgg1DCNTNAfRjK7OWSD
0JMHzRhgFFb545kfGwN75ZUl68JZar4rHp5ib9LLHb4JsT2uDuQi53IQA7MwTm2JXfQDsz3rFjQ+
gZ/9/aSXVz+vacsigIi+r2U1hMKLpPfpXlSKTOKDKDDfDVt1uQ8g80X7DBiaiig+zA8CQ/4Ol61X
JjmP2QTsMt9NWuDTwGq+PZKWG5xXeupfTHFoGPvR906lu3XiTgq7U8+XEHB12mS9zTHKyu+wWY7u
czgz8YMSVwjCFJeZROkFMgfMDEa+YIyXmyKpUCs+RPQ2pogtVrS3TRYX/Wlt/SrrFgRZS/E2u2qH
7MBlFaaYwC4TLmYkHiAGqzfdRgq7Sw6qt2NY727oD6w533SVqWVSYC6P5E4vJU0YJjtKn5lkqmwd
j+11s8O059P3D3GvwIzklvJJIATAEf9rsNkjoMP6myJ8IihYliLbMhc76SWnsH5X4P3gkUM+EpAm
7XNP2PU895UZcP7WV7RO8aYwX8eMy0e5TnkIPt0Ppyn5EMG3bxkCcwbbYShHu5IDPPgSR4ADUdIt
L29zBnonxyW8C35sSGWm1IUWV+dfMPu++Af8E54FMcHfQa2ZEVZy0SssfgfBN03R7x9eBdakHpDG
FA/gDsn9sCSg0Z1AxKQr+PhSkGBFSSvwiB1JnP9RblIbADezDBKQo7C1KYwXCUcJd8DR2ZLY+BXa
msGkL8EXTmyCNKo9crcp6Ik5xU8NTccEYa9Byk5Q8v7llzHJCbRUl5HBaP5vuSZHD9zt7B21MEpi
ORTDJ7q0sjr8NtzDMlIMB8GdpKtQ4uRpt79TY2L0D+6YdN3tmYaPcJd6ZDLV13wDqRP8kZCMFZzV
D0NobQu5iZUoAVJjYd5zBqO9tjecbVWtKsuY+5QyESGaEiwowAqVqFfDdMrkWXPPgBZE/j4ZTS+V
u+JLdrdcQudJ1PnxMxrJXpj2Q66m+Y0WQC8dnKdtnPTgFdvovJ0npFaCW1bCXhSgQd9Ap8qRP8wf
JAC2KozcLvitmSjtykp/DpN4xGUXWslwhWKj4mJ2a9q6OOodYDZkcHa+4/Zq+Oj/SPREGV6iPcFa
M1o02ZgaSE5DD89BnIi7E90rsuFZHpFs7zsyml0TnhRao7+7R9rj9hkhbPYH3D5w2ePtkFTdQAzs
m8I6Z2RZJcvh8fr++/n/0evWka+CbVvvIgy32fV7Evk5EJDDnAcdmXz0Yxua9SB8L3u/m1TFx59S
5UWpa0tMmDGWkxwKElpj6vSuAtQMbGUAsCOBVNnPsrFJXP0tAayA45DK6WvcSCt9mAHBvZL0aLPl
UisfWtMGtjvcV9L91G7qz1RGJNrbt56fztmx0LQuV8GCqRhA3D5Uy+yb6H4MbBJXJjTLwbO2FwUi
R6dhv6C02XYACATfwLwmoz+gVoAuLGqaE7rlzksjblg/IwTwwJ0Y5oAQ+cPTdXtkPRSbZbszh0yE
80VsE58HK/JRuHZ2FzVA1Vj9in4KAv7C57m61WosQwrlqqJp3e0xa5VV+rszFnX0vlarOTeE0970
2pinTUusnA8VGJ/Hn64m1TqGHg31+4xLo5XiL4JBlVMOz5xa/J9B+xnoRrzca/AN/r+hY3a4UclG
hBijZnkv54Si6rkSVolKNNSi1a2fZkN/QoKb4uslRzXsQsaa6AI2n6AMNcMI+zK24aX5iEVjLBex
CGcT5cD7XTSpnGX414KgFjo72+XfkwXDVFa6n6KneojL8iCNMhHZPjkJ5ntK2UwRIIecfo7ngay3
pLnWLLOZmx5jBS49qKwjIEkaVXMYyT2/ocOSKJF8IqwGR7nqTOibUjI/87bZ4erFjesUdMG2inNX
QH6dnFvLP/wtRbTHEpy+0EcX+fi1fXwaio+HyksHW89moO9PMSZtvSHAbZUZNeozojhPT3O5/Rwo
h33Hk9nIFPly4PCHMMnk3zLc/rKcO4rhRo6b8gHiJ+bkHNUg2m3d8lOCJkBiwrQbgkBhF4/oFIbt
Geo8OvpJC+yHgTPXFaMEPD/T/hRoUEtUppck+uZi4Y1S0w3XMAujKdjvL+et3KP5t95HNisXTjGl
+9c5s8xMHSrIeKu5r7TRCnvSKsz+ob3by4lZYbbNDXsOjF4NDFtq+AtZLmSvRDfYYnCjVt4aRuxZ
C1UGPKpLTJ0Fz2lz6QQ4llMqrY2seO9FRKLDuzq2e5hkLo8Q9asihHfdNfdvE/1yWm9hNlMIEfIy
DFkH7RfWGHtJ0N4Qablx3XVXnj151tsTIKayLuDRfD1kjkUE4zSFzDkf8Dw3eaKUZEaS4FDXaD0E
56vNYO3EjcbxhWk3kT44bN/wJI1EiFeIBtJidyl2HTne5c/I7jpsDxjbsnnLmTkww/mJ5Fq+JOxf
wa+FVh9RCsIXriZqgxNczd2UIT9h41nJ5So5DIVnmXOA5O8tmGa52rTmLCUBNVLAT+n6uEkkTSI4
SlfN8XK7S8fPD/npsaiKPODFxtXi22vkR6cIYuOYBa1l4AN5NQihsKZ4Enkg+M6ufVR781+2JdHM
VmljnFeCDGBfZEjJDhLrEnRE0/zAaefcRh1lGwuFWRTRlb31TyHO+Bbd2wpgRpEJc7EFU9NQI5UI
7NYnGzIfpSToSZIO2q0CVxO8Wk1YOY9OpTvbUmFCBGj0C7zMzDAeeui0ZU1jYIvyZsEzwXNx6qOT
AiZhz813fiBjt9shh/nOxhM0sYkG1ic8sTnNR/biP3T3EXr0ydpiCObCGXes/WJ/4pL0ERutg9kv
xXpcNWS9UQ7Ppa9OYv6ecUGxXlnnvtz26yXYmTQGEFDQJv+WunacijBQ5Nu/m/IlqMI/tFq4z4OW
yW+22dbu4koyTMzP4bxG7+j9lJO2E9dpyoe9DrR1Uqes3surwm0cJ/8XECvY5ZBjt32eELJCrwSA
M1aBkggCIyYeUejlmtBY8ba3qQ2Jk9KRX/h7ZLuwLQc2O+YFCg/wEyEbvYoFOsiewYmkpWDfVJk1
YQ619v+6V0bYr6aYqmRbbcgr/WKIl4Yayz81Mmd1ME72dqqP270Z7QjV8jTsDjJbNJ5S8Ocecn+8
w406Y9yPuZDaZfZl3/BwxuczSLjvElUMBg4RDkp6t6SVxwooA6MDDPOSF6PuRTBsFPlVRQ0qBi+x
8mgsTWCU/BZfmwzZz+AaELd1bTP092bJLrGIv2EMmxTj7jDadvapCzXY2VXd/ixCjgp+CX6vJ8nX
oQX76Ch5li3fLbd8Jm96tR+1c5yLFsGgj2KvDegtFmMTltNH/SKFeD3a+nu/t8nSNTI7CRdGU9De
TCRqBJs//hQiltDLC3cnC6VI7qg+RTbwAV8e03MsbpxOVUK49dtasD2L6Sn10R0CUksf9rT7Pr/A
InWSxOQ8NI4gsSJSG7CdjN12LJgx/dTCdTL6wcxE4DajMi/2mCzslNz0VpNVW8aVbft7cGKGIi1e
FQCgPR0wNB06+YtKLPYkuc/Xg1V/72W548Ncvzr9tSaKlZ1lJM30swFa9oktYPEv+kaCG6LyXwik
f17SNIcr0eZ0OYP/fbzTEJkhUo+sXCzwLPEaPZuO9gJR/Po9naqELLQfjaphalkmBKa2zUhvCUYT
9Fhn4kHPIVRu5yoYH4D2bGTzvRFtq8+OC+T/boRS65YwIlftkgbzUpFogpBu+I9wg6SQyGtp5Yyh
HEPouPEkc5srt4mMvK7mgTc9T5G5mbfqowv0Ku3P2TY0HMIcRiZmJz8zBQka9EXBAeCNAGERvgmg
2s012DLUpvVmKixOOg+oR3KX+aPQMhOQmOV1FQYfxdoyTng8w2d4KbSCApyGW+Be2Z/fXJO5jziC
s4Kvo7m7eC5d2ClOQWuoIKqrP4M4Or2s1wyOHUukV/1LDyC7xDPFunC0EvQwejvJYXHoYxHSsaXG
oXPc3d++9K+NTe6qEzsEkxOn7rt9E7Rw6P3t94MZrJAx5tjCrcOC4zIEhvjNWzXK18c5tCfg3RcH
hW8RFEORYaN3uoLeOJJu+EARUx40uWYCz/pfkrO9P48ohyYT+HN8FGI0qR45RW/rQ2+zxl7pRMNk
2/PHqzbUR9TLY3falIk9uDBsltzuQkZbHSu19Wwcp2mdQFvMocH8XzDsIc84OlH3v0usCCdOBQ1u
foJYBEt0W4M19KOO2R2xWQnKrnePtzuPAtBS/WFgkcy9UTusf8o8UZWXAbprTVqByThpnbvZrw91
wKlxiYp1AgRp0ccsfGFuOpT/Au6+Ts3wdzqDZQrweGR1m/VdII1s2DfVP1mYordYzj6caQnq4dkn
QzRrFebopu77B2OP6z6KPxOHGSHQXBcrPAqVq9LRzgH9WP+HCZSTwYdhPzd5IdMgDx26yH9GL3K2
BOCGj6vHbAe2LwvHCGp16bVO6bOyMjtjo6RXdX9qyHp62aN+JqY5CeDyNTZ4OqikNoaWz+tOkruD
wM73AdWv4ZZeEMk2DHjfrvaQ83Pu/PwZTKrOn9wMw9XORPI6T7i+S462/eE0IPvfldtjTcmJ1XAl
vL+riwqrh6hgTppdOCzr5QNi/7lzqgC2dEL3+Mds2c5AiuCFxxMHoNeh9S04A32V8K2goAo4knVs
wFXJAM9Yai3sxgRWFL8cmrjBymyyeEdgfGnt0papur+1gLeFFfBSlVa0G1y4HsT2SjCMYWUGHFyR
+frMeXe4wu8yhifqn0zvDsKtQ7UVdoSZiQ3vtoTXE+H13aGggRmmM7pzAHSZGE+ipO8Q8NX5YidV
KkPsBA0853mY55zn0ZS9wI5Svowt5pGa75IEaddHFv8J9Ljk5OI6aZTengMJ/W4RzuBpgIVZnMqw
EaN9E32u8mNsyvmvXfkbLAhxJkJHa8aeVRyhIOSeTaol7YOGceySfUHJEs2Cumi6Xe0T0MVM0FyB
pGrD1mefiaxti1OLqy0ZigWUb8zzKRz3xAhlpQEnEsCbnJ6wv6k7geSeBvftxaXdrahVCYPgM3BG
8bL0focRweDdbexL+IrfVj/YMV17Fq9Z/driA/R/CQkTx4zM6BqbEfLgF4Ta2qffmhlbd93l48mJ
SKtZQkR4s2ulJvX1wJsZz65HiI2F/QG0WvCoNO/OhJOlec/CHV81idC5viW+JUicOFMC4fDTx+D3
YzyPHa4wtwnrtkQhI7JJhtiMq+h6+siqwBz4eFNQrtT3g3ZVEBu1d+sxmO4gUb0KcjGCvtYzr+jW
yYTMI+erIB5IMXn5FFOEUscM09SoBuDAFgK9TV6btVGMsS9Ak+xzYPrbxherzDf0g4x/QXtl+tZs
m8LOcc0G2NufUpEb+mnMT24T/rkszNGpqZWagwbaXVEFRyJN/dcpwNNqmdDlUt+qclXVCaiw7sJ/
TFFMPpSf8Q3KquPNCQrsFGlBnZi3DTvoYfQtGEVNrV9steVpjvgySS73rIfz0VqUV4Dr4vR89pvn
6OHo5KQjvAghaL32GEsC1dVbfQkqv7nEzD94CfVmxDpZFui0DVZZCTAVGOF/qtqfncpkBKOguufF
wTUcDLZ6lyaNbm17CoVAEjiKarymgLUpmwtxCS+KhSn50l4ejm0UUBnmHocZZm65UznJoqXEyUaI
vAZgGuXFMgx3oR8RceXGEh+lQXx2TWG8ytkbSVNRoEaebRNgP0jqr7OGBWHBx9D3ZPpvzJsrmmQ7
/N5XFLLVckNpwNn9PG7jAb53VZzvCCEtTaa/XYnq3eNHuuNevkFhBfR6ZFNuQ16nEecZ3zJkTXGW
bOcaJ3+AxmsSHfbdAuwWtr1ePZ899vwKdbEL1Oq9CNu8b+GLJTt63UcXFXGqk8faTRacGrsfBM6m
T1MRLeo+96M+iBpj9Gvv0EvEbkXH51d2VIrolTCcf0gu2ZlK15VlAthF1CHjhmQTdSr1GlPPDiDh
bqPGCfMZj5HeEzQD7V6lQF7SnckyVZ8GexJzJZCRGmYYGoJFGVNQnxazNbcPqeW8104yUPISe8at
1LYw7hhlGPKH79c4keHTRyJw9dC8pcmLW2UyHlQrP8EDPYII2X4Ft535bIFdUsk3/Ms89EpGqVSc
F1v3S+mZOoS7rSemen6SsRqzu4/fGd82d9VhvIBEBUp31iIhLW4Q9UMLmB/nYzeY7f+9+OMJj9LU
4jZ/VnNeMarrSG00qmA11UkLDGXHZO+vmhgH7mQemKaygaF5ChONOW2pkugWYfGaHdb6YBFhOGjI
Rt11dIkDqEBFAWyWTrauMBRcNioS0uBA3YF0nU2BDUksqv+UarR8UQVgiRxoINjrtMKo9kNJPp9W
hCIP3FabvCiVz8v//FX8Cnv9oPfQ1BLoS7E/beksdOq4ca0nD+M2zyBTGLLWYUvzjZsxATJFHKlH
s//lTnMxIUkpoOoRGN1wRgt72PLL7YbcXf3Adm35MMVrWDmnlSl0lhPkVXSm1cyHptMq0TZ7xDUO
bmAC7GS2f7E7ew+e1DtjcDQxUVErz1IJTOUE0eEZtOM+5sAUZyheHjTLVE6m6BKZEwUiFC+TYVR4
8vD+LK9OHc+ak5rbFaZP8J6rwp1RDKRi75XtdRL4pKXuB+xdxi8AijspHpS5D/fdUILj3fHMXzoN
dfCmKRoLOXwArkAqB/Lym+EHY+tLBUYb4BsV1u5y31mf2iBAy0YW8Ccal5sl2Zq/hLR0HCLpN7QX
Jjt1xJYsdGe2nSgqCz4cyAZATCoYYSnzznJO+PwN5+BT3YAiSp/iqDpyKQP4Umm5yY/x7va430a9
DBjJr7Cg8UkroyRZuCvUR7VdyfsSKCyxuL96cLVWVCVj6lBzj/cf6c7Y0HxZXnCzfzgaXO1FJSoT
LAbKL09jP6Qrce8XsoS39oxnXE87cVxLQaZvP94a6+5tfJHdleofkPpf9QJJSFDH9MDMk9ekEGgm
/TTuqza8UlbGEJVuIUSMwjIW/HevT1D7CROrkQ5UXaYOwhlGK8A2ZeHV9LYzjfe0SMxlMFOAXfee
N2VKVg5HuSzOXJgW2WmgsiFnqY6Yxb79y4NUdpjsJzsWTAvauXLH18cwthSk3f5zwaEXM75tdYKI
+D7uDN2bExfu5U/veRlUOV8bXVHuMw5BOBHnIsRMtN9EM0HbVsFDHJGetixEluHTqdLNjioctkl6
O8ryxrQQkT1HsAfCLERTA74RK3HIcNX/rLcKSRKvPBt/HMC+hbMUbbxD2vFnYFJCvkHWL0KcwBYB
hYww6Ix7mk+a/ZbEasEZkVFBYC5CLPs/r9V9rWLf/TX8GClHYV9gC/aJnc+V5cKg5ffUjVOXuTmf
tusUo7eSpgBiUbmp3onANj7AGxGNWchWKRi8y0sGiH6+25wN8+6N4aarrItuWlhYnk/xYIt26D5N
m9yhr0O53asK4eSmlWVUwRwhT7Uv51TxbLjVX41P+RJe8P/MHSYBtM2e+yhiMfhF7WDjPLCA6Z7i
IxE2iaolAXBVe6kvxFYMysrhdxgM1nyTPNDShsTgX8ha3VlPnbknJNa59e6/AkdFqrTYOoox9Hkc
TAMyRBDQLbpX1rydFTcCkTGNQc2LT3S2W8ewFGfsWdqrc0lL+gbQVvdTcKIkxJ0/HLyS5mr6QdWw
cr85bN4MevDtEd/LG8G6tXMDx+KFWrRD8/tAUhD+8GADIYx3E3nt6pqyL5ejENv9fbTyOjQD4oJd
ONMhXdUzTJ+tiLYQSp3EamSB+/iAs5FIh6Fn2TaZ6RZq+/gOJqpbUfl9RElayjNlIJiEvawWx0P1
lEjQkokdZTGBWv0dsqnrgzhGWxlMfDnHpOFwnkAdXUXq1/YSa2+nVSmN+xjDvd0opC62gm8GwWfa
/UxDcz3uKKVziGy1pZ2sVvbKM4VmuQTkTtMs8TPhP8meYfyv9+KbkuZvmsVXCwQ82orOQD536b3P
XUksjVKLyWmf9o3uPumKnin9S69JHJvVb+gybHfV7bvT8QxOXpSjXTOXGf0UjMzDYSnIyeuUCNFN
7JuFtPw6t7cbHe0KME0pwBJ/W11mVHN4zhPbAuRKynpyPr2B6E9wX/hyaDzSHsNpeqWfjiqjjRmU
5A2eLn3yhQfnwCLpY/zvICJUEwEe9y+r2+V8t4N25MypEYIW9bUZ7rgJSTB67v5KsonoJMFFEvnx
5qZfTQcCZ4oILE9VoVj37RhNn+IKf5VLc+lWd4V4K2lBClKgYbqlrXBHLC+cNAd0TOZiEkpgauqP
M9VGJKoHSDJdrB2r7Wwpe8VIIaVjtETet1xQkmzeCHzF7VvDKr78ib081CMLdIlyvLT1TyhwkGVP
eWgLZZ2xwsAQ/kdHF3cpiVeucrdbD+EGuZ4J+AX+ZZwGmwKMQ+lbj+SpzZUUNTH499rE9VXcbPCM
SDrz0Ub6jZN71xbpcRLdAFROWMgJCnwuwd5bYSZ9mRJAR77JiE4rO5XZpFrJbSwOaiVW9EXVV+Mr
S7ibxy4NE3WfRpod6dZ1QFYuXTqfCXTI/kuSDIExQTjqMDybuZtzf+va2f91rGUI4ucAzieOMUUQ
qEFIQTnHYCJI1w6VLsX3DCzUrRBkCNOGb32lFpX/oQOCpgyKv6paqL2FGZNLNitIqsxK5Im3UwOo
XzAnw2um4/aozgfH/kx7QgtgdRTH3Kit/Z7DDhyVa2OE5IAaAT7AyMYZmaczz4fGisNsVR9dM4VH
nMf1HjUBD0ti6DmIiTZbOqRRzVFILevblI5gPXxK/s5wxXEVLNi6G7JwvDNCmdY/vVDRE3r0RGBu
cwLPsmfAW1qpYeHgrP0j349tt9cIPUkuLGxwSelWjXMe4PUdjEnhQu19uPbZUTmcrPV6K40ODE6H
u0T/Ga7MkfikwicFuzJ4LffFW/zMD/PSBfgS2YLHwJ/8GVEXWBIKuC0igPmBMX5ZBCkBFGh9RXbc
WserVZGE9dBDtrbbbS0hNIjCHYwXDYArgtRMkf/Vat9oK54a8O6iXEhozTWseY/3HZEfRV4MDsTW
GOAUlnkc6AG/2DkwBJRRHa8G86c5/87nE2jHhuv75S8HQZ5Fh/I15VTo6bToHNpe4Vsg4/2CY8zy
mmu9AkWrPpkHaExErw+lPc1vPZSN0FXpB202SQ2MmmGF2sccj6iIrT2duDpyS4svdW4115ITH4H0
bdZ3uQtWFsE6WJ+rQoNmnHV3ZJZocs8oweZm103cscI5b6Pjr1ttdUS9XCPZCAxJwvis0GrKXxpR
lqKMrXbI2Mh/aaZwnGyMBs6Ixz2Qbz+rT5+8SFHfzW6z5aP83yJwr3TwUy0Tg16W8MZ0FEV1ihFe
45GBbJNieSFXw1BY3ELtpg960V6EFH9Kr/Q3Vwts8fWH/FAqNs9zZB/pY2E5/2d+jaiiVuJFWOnU
nApFBQMwsIC1PBsELzfulwtiVm1ADsvVREGovfUPzvLiOmVvXM135NwENqNgRuC17ySw72NjKszQ
eUR6k51zAO0i2coV5FBlLntHwDSGpTZnOwsvxlvk5pN6cFqE1/JI7h8jVDAKXsA8FUd3Ii/kHDwb
9R9BNmJaMSM9tUQ1dlW+yjPtQEla/ZluHQq7RG9dUUtb/1/rx4DeyYg3uQFj4PDeeeeHyF2ahFV1
K+kSJpWVcQGBV5tEuds8byq06TmsnbsH39fHykxzCLHlh5O0/G+Xti4D8FDCDkyEARsyMT7V1aJG
Qrx+EfglNDUZaKgSBPd7roOQM5slUJzbvdEse9SXoWjJI+ZU40CnWD6VM4SmDzfL+EXtpBxjs3O/
Qk6vWAFsIsPiflCAwbROTBMhAqwHIrZObtfUzIoi3Hn+mClWXqSNV5cRu8lshbS7RecJ05ECiwnW
kkX17Rb3bFxKAm52tEN3V/VimU92Q9ynYoP6LhDsAz7ir5mHMPgdIBYJevHzD6lwZPcNhhny/B5n
54Wo8+ArRL2txE352dA5Asc9r71AQjuyWOIDohBAHhfqOSM3ZkyBWixbEwm537Me9pZBKtYf+SLA
XrHIPJRyesI1qJn7wRM3C+oO06YFZScKRWohNjJEQCGsFyHhMY8RDlxxeSIU5+z3eCUWn/hMG3f7
QXscpRl8uA4KNIpovMBbCwBpS18Q6FgDUWjvD0m/3QtYf/sQGtSuIUU1fFyK+fZtpFQsx0yvXOkc
57eFI2xaD4XLM1G3HXiElXiPao761Enfw+uNbtIiUX/nfuNbTe0HJ2aeXmMTEB1fE6bLORXn8rLQ
sQYTMHRpQtVGUbjt75m/AtpomqUU4BKcjn4KNaLakdl7yYM6gu8SGNkYTK2yz414wir2xOQ8q6cm
PHCtjly6evuffKNBDZYCBVRdn89sTKPfaMe3+zua9oo+raMXuzIeF0zJC6f0Py90EYHThYAY/RXF
48gFEKo4h6F3Sd5jv9xR+5BUVz1HxgXh7EMb/Om6KVEj9w1V014jatyn75LbaX6KGOaE4YqjC6hF
7ncRgVbRGRaeI0qas2CS9uQdCvbARoOxiw8suQKxfLhd+GvwLys6UjPCh5UlXg+2s5cRrvcVe1Fw
7f3bT8aOEzwZASt/y6pBWxQ8wXoMyGKQOuRdC3/hP/DDWBXJOjhzpWncGFDzwd84wpptD9HU7WUN
zIYmIvtVoLGAwGnjRXei8d6WaKrwov9ZFgaHLwrDs0ihnKggYvQWCcpXD679KOiNOSaRNDOSp/S1
yIp301nxA8eyjP7U2xT3scJtAWhbOv+cIWvGlClN9ms/HQtc73Jl4Lp9YQDNjhVwoTkMArf+iwvs
P1tdzHkYSAIS/JuNnjeZf8k00ZVKNmhp8iyEynYaGYWtwOP8eY5axYyg7c+vjILz9MnOX/NkDKU4
h7NYUTF077kUBP01/+EUtnNDX3qQecSFQfTP2/tUQg+Hcbah/PpQbzEYAiFP3CFLXdxMBMs8cXIZ
ho70MVlaENbIe/9O2PgpTyFHTUrd8qF4gzAFZ4N18z59E16IJjxJrC7/cYavydesFYz+D64QJUbR
tZCdrIthK0uFccm0wOVArMxH3Scr54Bx752tqnodwFVqq95b3QgUByR3B68z84oay7dq4vA1b7GN
0gNnEiBoFBPsgE5LzO0+6SPMbMBLvtlap8T4cUD33VFS/TIJqfDdYT8ykDyBaV6dtyy/puNm/DVw
RDmblIaDRvDqsi1L72jeZpXgnDxXlTUXG/RGeXKlmbGQWKjcWctpINFd2wUetVdZq0xnKK375154
uA96W9cOcAZmDTUYRLsjBWDfMJV4LO2D1NO7Q9j1A14duacX24mg/TZjIHqRo7S7Fy56Eiszh21j
G/wVfJC4npvbtJOsAqTIcEYQzfDpYJ8tIsq/pS7FMLjXvVZZTef+KvLc0ku6VMu4eRtJcrF3dVnx
09tEoEdKRSOQrPjEr8jZhRqOCWh8tZH/X8NueSc+xbt3VBKTZTI6qSVpDLdUJT3sHxJLHlF/AQGi
HJlPwMaTbS0xghMYjSEI2qovyhBmr70c5HWktDjaIC3QtbHy5NODfaAthJVd4QJD3fEyZpNrf8DC
6ha6lXUMOZMXzAOv193SubFkS+IGyUYrrNyKgWiWbSruAhxgi1toNPZ4Mec+vkWfs2cCULgpbMze
ilEB5WZyirkvAOUc+oVZAjeAq2unYGhyIoaEBKLyS2RImFaz9krZMkXUthzltmW2L/clAQVSxJHk
j49540BsNxASSsDC9CKb2sQsXY6vWoVyWIsMKIlSXVw/0sqULZoIqRZCxTuZwz0CLAeYSkaxQmoJ
uGBkqO+CAAwIWStRyQIsBEw7WzSgJZqzQjUBiOp6s21cbGgftE0hU4gcOKeDVDQWswlVTPcd9Ewn
P9YiU6kMY7CVdshSfyCnV6fh3qQ2m8XRkk+9wVr7D6dtI2SYSCBrd/M7vuWZnIrUvFb+k6hHkBKs
Kvkj4t5c9yf8Ew+J1GpKi5sJosvGUCB7BByV5+A1prEcopmNc8evjEYL/RPbEbS/gBMYh2dERpK2
qQ+o1icR91R7zMv2JlvsQUjxxHcrdaYpW7j4km0fdLfRo0GPRHhK2ZB6v5UCEy9rzcDo47VeeALT
QBIbTrAaJ+8x93QsJlUUJeQMo4MG/ZAvMsavS17a+4F3nDuGeaKtvRj+F2Z1cLHi2RAmC9XBkMxV
gdjMXl532UgYXtW3+1DXNiKy3iiAmjFqAvkJw33aNUQuubl1A6Bj+hxOzpnxAptRmJaZPLpJqleg
EnGmpEfLeNakSQ0fiZjtniohhYoYtfccf1PN2EWGR4ckG6LQZerYkCWeJW9zTpwvqKRMwFb26cyt
KKD1gwd2NGqegiGsmbdNJfoMgFJlMNaV/hAPoLyJmthPRguG+0FIiX4P5cP1MQyqrL4IZqd66YvJ
NWas+qLT1mTK8xbsRwXEqcQB88dOBrYvHarWCPQCEvXvVpCL7u6wgsetKgFO8yIWinuup736nDR8
1Bx1KtkWGss9CbS8iEzYusiGbr30Ay5An/t/ch9EiaPra6Gsvrzx0315901SSzAtUHxXbeLt4L1m
LG+Rh0UXl4REOTskoi5WYQE5SVWyBfZE/4FdCJf69cyvLUw7mWp8WbFFLegOWaSX8jjl9YuW4DWW
1tRCYCGVX3BfzKYuT2HUpPktIDCuV8EDoNQIaSrS5rVp8y4plACUSLag3KL7AP//jCnHrAPiVcMq
CJLRr4HFIEtYC1z61pe2Lr0poIZlchlsmnFpc4tprdhhkEm8+WzwunlCvxqr4rjmlh/PFl/Hn036
X0JjK7/P/IS3Eb5/5VMRfZA5lFP48mhZGpGak7kgLJMeC10HCJMYvSDeDf6NibNRj96avKWfrFiY
qvIeMdOhTWFkVeYI76fPwDWzmD+a38wPOQ/iM7yF+rB3und0nnFZH2Z1uVJLcjcTbW5y5byAKTe9
M5N0sbECEoXhNgNcMTOGihzQ/kCVr0zuGq6xQDc9jNvrC01p9tFczHPcUOESuE6LIXdNjzLgzooW
vQ3c4+gmJeuz/GGeGOMfGHdSrlt/6XkMHTJmSS7Lmr9l62A/AzF8uI2UfBo0/Vsksqtz3EgcfBRG
kJcLeFPD18VssslaY0osnHFSmobCjCjYvpdIhMMNaRIbOBL916NzJBm2ZVlK8TuDcWdu3S28hwYu
Vz5C7oOWL235WKlCO1cr0XqZ15sxlpIlFf3KNt9qkCCo2BmUaEUYdpS/sJYeJguOlvDS/QKyFirR
8qQtJOd+Z346rW0Dqw7jXzeQLyGEj8HPUZzzrdjBhiwv9nyO89y7561kFo0OP6Y4VWlsO6RQyeMv
Wre4f1ZnCCpD6AqzTMM1R0E5PR5P1j5dS+EpSnTXwbt3MZZP2ddb003tMznqkwWw3xWuIBHTmOq+
zgWaeQEKxHQ0yIePNCLkeNrYj+rICKH/uTXIAMafCl8Xf3jwfBdqPGLViQO5jFi44T3in19dMNXZ
rF4XSEf/wQHEWBPalscfNf0QeA67rZOtIieTy7PI/oaLOAqAzvTmBGi3q92nnC8EnpVwEc/gczgN
HGrzM249hBxBfvlUs51S+CVUjWiWAxkVX7WvTpV9NZdlTRvh2pyn6Xzrkt4ajK9dj22Q9AQyI12/
wrsNlCoO2KbTdNq9n71TG6lk0lExRSpb3QO85m34kS4AofYcjFrQ0bqQkkoG2tYYbdE69WngF/Bn
wjXk0ya5ahgXyf/hKDAqlKGC+hbeC+IVJzHIzCIAwoj4xQSR7l8pC9KnIGEHVrcP6ZpxEp8bVX3z
1/6y3l66AmE16ZZQdL0/tZCXVkiwf6ULpbQ1hOvCwtI8gWdQ4YRTV/yh0CtDJyVTg+YPLYtX1H/H
jeDQ7ZBZryhbKogGGU9Yw5+X/Og3GeGiR2VNwr/xuozbGAfTOf98WohjUZfGebZh9m4lLepxemwK
dkQ4quyeIwDMNBU8aBB6zCIGo80ZwWLnV5Q1sbjKJH9LQNqXIX0jjUGfg+FshMv2YSHqHlwgs1k1
P+2QEjRjm/0H2gF9lb6ynb8S5j5w/VSt1bsdzWjoHW914E1fDUjjB5pfke89WFCjEwsiV+gAzsih
NLdj4J2198fLhf8wbiRkEA32BU3UpVqwW58t7TCCfiXu0bK8Rso5Kbie5Q/a/ZX3AQUG17KwiH5a
kwt8iCcPqY9V5Mi/AaKnwbwsOi8hkzy+1cYjNWedFgywSANpzh/YM2VUcV8QLakb8QjfRcZI2KVP
d0ZfHp1W1J7t3zEpi2EnCay7/snwrZIVQuGpqK1kxGd0sWMc6zt0IppbLKACOcf85T77VVC9BnjS
+3q66R5gx8Do7avI4uBHfQs+WwpVWgzuxwFnUTHa9xbxEorMHWZQY0rZPsJO9nAIXaIr7fovFDPT
YoPVSZbVbikW1NMwHrRQvF3ReruW/Bj7gkR1t847NBUmBu9fK4tsr8Fp0UyHokaui4dDACbXMOTv
XRMKZRrpiMWtKFDPX7wmFc5IgLEhf7PDAeSUoVIDr/np+bGtkdoDv00bGU2C8nsc1lM3f4csbNwO
RrAtdA+uuPQzdvcbFt6tG7tpCa+oaZrdj6M5wwcvONeBQzhsLexHzcYp8ywOuSrioo6vKPdiaj1U
iVxcc2xxwVEihzcrToU/GEMYVBblfshUOuoOG0XaMlyCkUlOhxlSyClD25RkrnAQBiaMuaEFuhvP
c6Jgnjw0c9rpr6ae0cS6+51t8iOLgy0owIhOkctodjLLxo9Dos/f7rwMuM7d6x+AdcDUynQXT4AT
oJewvIkk+T1joW2pLau4dgOubvKwZtfeYs9mUAC9rw35LAm5hRLVQ3Ur2OpfEFTpfyiY5+cncEKP
2yKMqw/G7dSjVyUifNOQOXWyBnP7P2TdbiIaw3aBn0vbVxASd5Fxjn5qHQVr6dF0ihNMXu48aSPu
jhHT+ZpASCZqOVBTnJTmVQDWfJEjNvAcLt3Z3fbHB86Yn2JasYeaXpcwLQLZHT+brrIVfS1MRH8h
yCpzYe8FdAxI3txIeOeRZXbdPwC49Pzb/UCet1y7wo++9wM1kubV9UwcwB6RuI8U0i8UfMRqUMFm
+U6vSXOq1a5j0f39zuliV3ypccIrC6kllDwgTodyRXy7BXEy+CxfoqmhdbeJB3QSjuJtQSRH4Acv
02mfad6u8zsPy9TQumL3Emrz3VUoo5Jsvmv0GMVYY5ID/cMA+rBKvW3EJq1jltScnbXn4t9jy0zz
+KyLULXyOIPJP6KhmhExVY75rE7Q6nnR4tD/gBCALwKChBn2R0ZkaVwXE/39+SkaE2yCNLvpTEh1
p3KYnnl78FrVgrA+KaUppmDIE8s7QFxYXZuDgyAKED5ZLnbQnQXuCdgeCWPSucULZ4nctaoRpLaE
sHdQ98za+kvULi15nAAuyVQ3ZfTYP0xrw9uvnhMzMav5B757ln99G+7nEYDplkeJfQeblgZ9iPPs
1SNsE80PmqDVcyegLCczK1+lHckm0n6BjGPYo31tv5T9RRVqmV2oZ0xtwaUOUXEVGgH80vOoVfrd
wxTBYOD8PuJAja4ODgIXonuA+FrS2kEhjGeX1+RLUNuh1ZqfLQ9YEI3ZTKyCsgrMcaNqdBJR7hU+
c9eJlqTdRb1JLJ4gpGxI3mRA8vEVg4bBSsCXlgaq0W3Ch6M26V68uDA4neFK/o91FtcoaH/5kVct
O2OMfOKjCKej06q2/uw0E2ill0UVmnD/HP4uBddCmzyY/Vh9N4MebhZy/2U1TpvesbmxtTT7YQyR
f7Sc93ybPe72P9tkQBTxLSiyCEqv5KD7OVtbwwtK61pjvaBLgBjpjLo6LvF+q3ULs/4Wz0bpyF8H
fXTy9T0kSZf1Dh0kMhOXSJWh7g+kjEI2oZbIeJdds24/j5X1SagrDVeaw23P1BAplh92VNrwQhrv
ApurDdRVk971yp8x11hNv5gR1FXOZ2vIT4QCPEohnDidhEpYWjGYlhHf4TY/dmiZ56WFMGK6ZKKn
wAepIQo35wVwVMB5oPO00fNOMgtIBxNlulL3rAATMKEnrpgsXVpeHuAQbt+UivRCf5wVnA29xmDW
733UzpVVsn9TMo6JW2GN95VlO0pUg2sAMotCSgDl/ZyOrIS6zqq8qo+lZRMNc21mVKeI1OKE4lHw
QBuGJgZtJe0xSPWue/WKwd0XLVPOco4AjTECUMoZkYgkXVS2tCUKFJoRguv/m/o+sr8KuO7kZH3D
V6CYU4h24k90mk/3Ow2iYysmM73yP6hNPNHLgNzd4BOSXoy8l9WIWLMs5WXtT+1yRjGOzJSrMpx0
ikCBdInvVtHCFS0LhnjluVMdCr39ecyXTRZd2yyPSloKBFkMmOk3OpaLYGPMrHp2t92Amw6u9BHn
GN8im8i0lormmOy1t6pBU0u3y/pPJDcM07eWU0hBI2sPqVPn4UDJwE4AZ1Ub2URPrLfhk4LXHOfm
X4BZeuNOGJ/OPqBrkStStFPTrsy3gcbIKk7uSswfu6lUQwVgXMqP3AIJ7KOaGvrainl341G+2ILP
UDCtbFD0j466i7W9AXw5dVyZ4xlN4ax3vuxOnrKGzRTkEnt1yD4FvvVsZCrOtB3X2vu7k1qxITIT
k0vg6aj2ZaNSADpmRlXcRSqqX0I47kwwslLSzOGsEybSKZvuEVC6nQzUe2TxScFSQwF7pnwXv1AY
pokbJ5UEi9LlnXU922tcwuZ6F6uXZ+anp8WuIohJYaHSu3DyT9gkd6ONG5LboBIR+KhpNS/Z5SOY
YBs5vCMwWivkjUv2D1AicSQgvfGcEj2AjLurXs1/madIwm933Nl07PZ0uMnuI2j0p1S0WPQaDhO5
iFkN7lOTVJARrR02Dd8LZvPeb4TfaVZw6mehhxf9NO4rjI5dhGrvmtt+Ft+LYKsJ66IGGvhrxYmy
FAPooLyCWi84rHNljTTkvSC//4FHozyZug18pX8a+/SqyBlwzuf8TuUtUSO4DkeybsCExa/lGVtM
06G6oT91xojszBTNVaDieyDY25Q6n39nJ9TsMib+MAZ1KzwQmvuF5t+sYLhqxUgrZa+80ptPiiZj
ohKpdUGw+PGFm4Y6AbmWvnJ4tLIiK6K4JN4Ken+ePJ+NnN/0TvMvP0IfMc7TNartaeKwh7Bw/jfy
6AFWNrvpcnc9EdfBTPCHW3aL7GJyfqgnaXXGWBz/kO/gZMFcqbOXBk3d51g6JD5j5E71IyNb30Nj
xhdRqI0zSwtosUUcy/apgjJUpQY+LLdw3FI+Zd4n1w/bT0Eu9g1FT1twJeUd2QkIrJqog4ql+6RF
/G4CK4IWAzxc6TztC9beheODotyaWBJDP29pMwKDioRnpOztHo5LYzrFgr/wk5CtIEmnpuLbLWaP
1M8ItfPIUKI1i5JctH1qn/BsN/Wl+uH/nYG/RDuHEzvXCTTnI6OwTyouJ7oyG6ZCBviJL+A8u9t+
EANWLYwv99/FvQhEunmFQGjCYRDIMxmjUjCEGNJc8LMjf8Xo6BGaVRj7aUrTqO5cNhdevGWgJ+BD
aBhZTIq9bAGIphez9cgC2jP53qNYtHCmbDkmBIN+NoOAn2T1MVxfVGG+qC4mr+Un2/ooFw5prd3u
U4oKzOjhZLINS3EA0DvGjqNd1DaqVf0mv83Km5nwftuBi0Vp764LyWg8VoPCJgQ21jHZLKJy66rZ
lK74alzzNLLBrChAKpIhkqzWvnxlARTFBoVoScjVQLP6M3n/rvsIy1H9UOJ5NSsFwNflgrQ4JOul
2Ua30jAFHo/lv0wncjiy7vBNs9CzCU4nkhtwlZQyP9AqxvMtSCo5BlO3OcQ5TwFHcho2frPCoZg7
Ltgd5niMq25MZmCNMr5212ivnOTOxFC2EKDAF9o0pNSs5aIQfYmul9tiawgZ6Dzt6h7g0nbJhsYJ
4ml9dmR1OuwWITlEq8Keqw4gkAQlb5jQukjRBsO+gDh6xElckI0emYbdeoWRqTDJqCmpnMVJ1MoB
uO1UfaPr87AOZqwfaWm+rU2cqUdqPUBBH5ZPgr1neeL0PfKQKsht1TiCjpWg9heq0w5EomXTwc8g
hGhjNoO+4vOGAt4iCfc1EfzFoDJnatxo66T4cgEWgQ8s6mXWOGhwfQEJpsHIr8c65nQGEqkzHMSR
FkVLwVvYRpDGKpI/xZJGBh3WmWU/6pK0PqZB4kI9nyBev5KR4nYyyvJ8H//Sm8kDITVHe0W/Q05Q
3Mfxa7bLc2iBZXMKEFQUSAgts/p6CkZiNnnaoLdFRZjW6w+IIWAX/FdXqYLr7h7bVffn2IpzOW2p
g/yk+YdES7PqMljo9+VEr+GnepdqBVg=
`protect end_protected

