
	// algorithm-level ORAM parameters
	parameter			ORAMB =					512,
						ORAMU =					32,
						ORAML =					26,
						ORAMZ =					5,

	// internal parameters used by both frontend and backend
	parameter			FEDWidth =				64, // data width of frontend busses
