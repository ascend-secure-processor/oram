

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GN5vam8l8CIgmRE8dP5ABoryDSiBLV+ADgZJSwS12QXLKJa27h7hqcxnr27D3n/8KfagQxPRTpSF
/dKmuNEWbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l42My/eB6v8h0gPrHev85RC7U1471f/o1uKWZ4c7u6i++4pFBKbtXtCjx5BOiuo92A3hmYCKUeLB
NIbfglWmutNJKte7qLs6OVd0eKQDJh21ZJJiRBRWmaC7g0YJBXxjVdM9APka4CTcHLixFiqxm2eh
82guMoxL5N14vENnEI0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I6VNXBMIxLCg22fCIAqwhvuFROeL/G+/AyQJ4EzU1sP7HdApHWNKcMHN2jGFZYG3OG1W3TQfKjZa
Ytk6hf7TioxsPD8DDpOt6j1GVO6YvEUjyn3x411b0RRGfnXWFdX0pxn4bohIQBOBF7o/lYsHQ75S
hLk3PKaiUxtTaxqt1TcU58SNfy4eS3TT+tsQ9XNNv6eZ//zNJvMLiWeZoWv5mQxASOEn4iTePMnW
eLcTCPajxwj2uQzRrn3TNvm8No8HsaMZ63yXpxYvRTDCVKxzpGfJAU1SKENkPtloZugRRZDmm0yd
500vWCOQX8IE14c0ZwMC6ZOcIINSDdSUYZLdTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7+sgpzjGGqGDl2uujOuDUd7jLioLdwcehjSP4iIQO7Y4Vs55B77ry4Oba9rAEzl/M9hWBP6FQsO
aIB1/HIepGR7rb9xPexOMu7DNfuOABC/JOI8QQMeuCMM/MBD4dRaiIkpcgys1HjRQMLt8VOLFf+v
vKUhrAE6RpDZ9pXhkac=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RtLvMG9HTn/rrueV9md5B4obbFsTMpnmFal/D9D2BdHub3Ql0guCZc2r6knyKDuSQmb3N4LxrEPU
66RIEb98VpDnemcd3LKdz1U6DtvmmAgNNLA29MhxL43y4VO7ZhOt8V6kPwnIxZX0B2vGsjs/M52M
jRihLn/LfnQT/EzhJmtEw+3rMHaDVODs6fO1UkY6gUYj/3iem+N7HSHYTOHCHbOQcbF+6ZHI/XbR
f7R68gXt+GQpkWCm3BpKC9rb0E8SZf7vtnsqQG+cY/RRmFKRAVCwynlZmBR/BJaIcUlliL6H4hmb
OnL/5G+/cQ5LL3iPmqSwBGVFEIjTDE9GuCy9uw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7456)
`protect data_block
PLx6doPv+4g4/fO/JonShi6piupiKJ7Qk0XQ+Q/GL1Z8LY5RHi7M35f53X8XuRz+NU8iikORps1d
BeufBbBN2lT8G2bwfTIl7Zel1UkzuUZd4RGt4v9BH/k2CfHHLVvAr2qutRsMCHRiRhJzOT4IpqnW
vXF7D96Q/WhEUl38A2SC8TD/08wQDBXVcI+X8mGiqIJUJYOfqs2mGdPC0fco4lKzn436FHOVmZLu
DBM8n29qSBDYV3TqjZDYR2WPxV0gPG8wByQYbxE2dejHqMDbxTOmVFn+tCOHUOn6GcRPmqF0ZCBe
Hks7IO5qSAjLOoOBQX3PgiWq03a9CktXErIgeAxozlXtCYSZHnJxizjc3eSt3gN3x4Iban7AEhhr
jDj5PDu5Dt0tysi3SJJMtRKgCZNLBIFk0ETaT2VSmHOwWn4ua7gQnUBt94p70Aefs5HaFGEkVWRy
0+6Bc0FoTk06sCmE+0zOrnwKCSRe/8uLDZlvqyJ0m9NSPd4unuiN+Qsb0EKnWDElJ/+g8FGb/Znu
VICfzYZGzTquogHTllpwIZ4DEYfdcpJuBC1FZymdAaJjJcWCpf80pMpZyDjak/XhI2nJXSswkV8o
vhrkbQGL5WzIQtrpOnfedp/MEZ+qngjYJCxVvAkKHhIUPL5i7XLw+LsGT9QPdUAPRMU+5A80FgiJ
0ZjojpYXPhFeK+GobOag8PBPByyK/6gBgVJlTlaX4lY/dMMkfvI2G+C+L5eA6S35rTocudnLs69s
4bl33Prx69FTPGWBf7CoVYXiKjmf3RAx8bCuw1zl6u1wkws4p5k0bvsEfsk80C/tKb4uPXiUa+7v
njthw/8OXnxi7XU9URdX2FqSULjIQg/3rzJ2bUwZdDXPK5xqi8DpIyfMIbQWm8NiR/bKaUK/unw9
k4PiQJIoaU17U+MnydMqoT7gqNQ4ae6DOUpunAJJFdbQSCBSUeV/ARIKoG7sNd162NhEB7pV/T6z
LjVxGFDHAlM1iTwj0X1TpV3gKnuTFB0wc44zKKe+3n8aaAfffoTNcu9hQgnrIj5k6ySXKoRlvL+D
5sNWlU5AugQs/yUvna5i7ZoDTIsMkZ8FPH9ZqLv3hOxpGDa99ua0ZnabihD4yfcojykjytQs4XMH
tCoGu9qHp5Pe/hHrW6HsnJLBzt65KQEjTUfYO/OtLTQxX9H5qgZRClndbTML3U4j92+RZvAXHATU
meYaZ1LOHGzVR7HnfyITS/Cenjore8vhsZ/jXNA+u419/TVJfAnyLR69ypmD7QSOYIIwddFk/VLX
5D0LbPcG1pTmqG+Yi8ZW46UGmfAaRqufc4Pa8+G/Ehobusemc3qLzwXMlswcG3WUD5g7ivQvOU+o
OPt8k/UgRlKq7stLC9qhgyxK3hTVyuOKT/k2MByVDBqF1WZp2nqEPNvYQxuYd7yOwpvjNgUbk2V7
RzjlGf0RAtVlNUH19nowLUfjUT7/nnGr0Qp0N9Kikz0kSoL4fZ9ht1bwrgEuCGuaB07KODlvqiuL
wlXE1FEfei7KnVtPnufgtHH8SrVFydvWCJVe1EDY3VvnQ7kbVf71ZelDemC8iIqSg4eBF42Jfh8b
kLUmIKd3MzcUHLktzLp/MG+U77fazO9ceTHxHqrSQ0l5OriQzKCYJox1Xy0IdyTALudWK8daN1Xo
7A+2b5S9wTNTiNsz3pk2PxGSh8zZCljFmSNG5IkSnfmwBLXR89TSnyUy89ufqphuEtLRakBMBGK0
qvsqbk6udzrfFkLIDTJbEj44WNtiptX/PbNjwKucFDc2ERp+hJXaLWVRFQGs/dedWXMij2pvtxCp
1rGOgxriQRGVD7wLXfEpwyijH9IuRhYp+ATTUDlmrgmmrj1qstn+c7hJNMPsPC6okij573LbArEo
JiJ+wJGEgy/ythhqo2dm7HmS4f7ou88nlvQX8YgYC5+9Hi1kFWF9EbJnvTa9zFZ47BifvRybHC6F
4TIYBV4853itIN99xoJ3BHvTMxnlkMDsJ5HcLKnfbvNjjd+X9G+e0AZbiSWEw7jn0Mb3MziAJ0kE
5DaqLvjw1F5g4CpT6PV6dk109Yf3iHLvHbq8VMvnd+DWwizL9UFH/aDeSM8tj2NUKhXzfzDNljgq
SsjNHwovNf11APLy0gOm8ORs3rQ512JzglTpw7T+t7flr/Lq9/r/w9lgbeKbyLLvjyKSjrWGWrBI
Z84jUv0rJ0VcbXXCHdTbnaVhdROjlskp8Tf3MMbA7ULqqakcrRoi+G6Rjdk+eeXwJMI5T0A76HCx
rd/GnA3iAsdCrOXnVxvbLKqpEXQLz0KI4QSShdd3CvssPohTIZ65Z94ySan5XpRoe+E68xo+sYkc
pky1WF9P6OoHC+Pvv63dwaFq5jjn6OPVaUDgn6lVUZe0dLE/6oxOS/2W07SfwF2yt8dbpsMF+vRN
r9IxQiXcOlRY68PUc2/dj5Wp26vUx69hfm5y83RM12o+3etqe6BBkA8heIflUVZN3KfIdfeZl2Tx
S4+M8mqcSI4bgf45bcmr3+VQdY9Fb7a4OCa0Tq2EK7mAVA/EoLP4AWlUJS3O7cmoBC7ItwK0tqtt
IugPTP48DkkyqwHx0xxy7jOurb02WI0XsGeEd96ILZaANJn81e/ANckRRhw6z1DSQ1irTmyRLhlW
m9tGBsqPdf8GftgiQ+6AYttlWcfKp1ZWzldWjEy1NKy5s8TYC72m1/Rc0CJYozvUC4nO2VEFq0Px
fqrm3vK26aZdGE8mTnk34aJxwmkXjroAHKxU7wz+s3yq5Ny+nyy/RxN3YzzsQEX8MIxHRDwMdl5r
v599BWmdsdvXgxWb4B28sfFUVIGk3wg4dD4ww2CtLKBWQMsjd1QhAtgGLjdSPKgw2/CkeKZ0gUMC
AWXXt9ftJeBvEeTT9+uD27ZQOyHirtyT8/b9sAXhC0LJ2ExGEsLLUg6iY+pzH4o0Qa+b/i0Aba8y
TfaSULHSbWAKBsvkolRCqeTq+TuFq8UF84M2+dF8FPTRZWsxw8vcj/yvFH4ZrX2UX5IBgnPKK86h
jqYPRhhmotVz3UzDtc8bZQnbg/qkFDab1UwRd8aVte2490dldooaivNAP6iaSG1w+YcBm6IVNSQg
QUJu9Ckz2Pvg/P7GAEFLG6BMA0gn8SA2dtS7pYuNgubh3tPWzZy9+NP8u/e3DtIFkcHBIpmXa6Ri
AUZ/ywGVr+6gmS01RT2ZM4gXOz38i+YyRupige3W4HYmD22suO3sNawGzoHmnM+u3lAaAqyxj1ot
GMB+dzSmAp1KhemG0cpw2hL1yjKSMfjXAJttrzb7XZ/2U2J8hZM+zjVNC/qiVI67QZdkhQC5HI2/
91bZkTC6Tx/xpSE1KGOpJ1aR8fLlvVc0o4KdDY3Rk53zC3MurlqC7gfjoNBOvcyjUrdqto9kikf0
mo/DpstSf2g+6R7g4LHJ/b4m6LV+u8shUqA+6jhES+FJ0KOvx/NwdXzNf7OLEiSmSQHRtSw7Lbgb
LoQEYD4ZARySzaeEzbEVMz4ORWn2BVWEgQN8dvc4m9VC7UMo9dItDS0IQ5HlHqLl5uYVd7QgIXw4
kEeVkGFo/opf+Qo6+NufOm197BoVvaCqumoU/TbsVbSm2VbIWvum7u4tYfPpD8qWMEVN1nDl9uJh
EdcUgSMB2iw4fU65Z9ycruKqFiQiHzps4hBguxJL7EfeW5wvgzSG6+BYCQYTDez/Y8vUQfsc6izY
tFKvOQxYJKZoOi+fBN0lOpeqGdOr4BwMN5oJaAe+vyRqrI4ZRS3ArGkttcxW3yHixjGkJ7waK66G
mKEbkiBIinDcHyF4ReZC1D9nmXjQDmu/L5z9QtQYb2q2R+bk09XgWqdCxB3yuNsV+goySAFkGLp0
Imp648VvfGKXqOI4WqUwG7McIYnn+2dZuae06X2SqjND56KY9YvdbmLvzyC340VDKZmg7AH4rfqD
aMHHnmLbWTYpfOZKyNvPQz85muLAlMwX78tGO40JU4IqGyHvGpa/yafatKg3fTjf2IEMGqrw80sx
jgreZzHQn1/5CZQ5m9kp829cKz2Rp3FZ2VUEmPI9hI+/cQY67WEwrWiKEumKSACiGf666E35qYtC
reJpOpcR1De7rL7clFsa3mz0O1m0dn+izpMd8fLXRZ0jcl1UCVEg9d9tJlVoctopCb0fTB2JfivS
nJD/QQHeY/C6Fb0djz1sNqLMnyjhtk5n8uZ+ju/Z0Ow0G/x2uGmWP2j8H72LiY7pXzOg89KGI5X9
pqkrtYTdu2b/WDW+pGTWN/zIa1FrEbaSzH6rYD1XhEV8NLeCNMN4d9ny0Cq/Z1flCe7yL+dZBiV8
uBJpHQd+WFUBwRqbmofCFsNmkbRP4YOyKbD3AaxSXIslbCHbAuwceczclZe3lH1J1bbleOHPgn85
iSJ3otCsA1fLVfp+W0uxaRUYXtoPDGXekJYmm6D8LGFJaBfgVvztsk/6tq/fice5YqJ+bl1g2C7I
0fS06Ho5zwK6H8QISSibExZ2wLT5jqiqsLQlglT83kZ018iI2+U/9g3S7auEpMsGHfFlhXvaD8EY
Wq90LvC7aOnm4nAeeE2+bZ/yYa38OiwIFGBznoUMWoHAiL07Qpjh5iS11WV6F7F0jzd/2GQDfpKr
N5T0HuBvlmb6CGet+3YwnEUr9663zgSejaFZXWcNhtYrPvSt42ImPUwxrJ2BPhZ16q59KOEYtwfr
bMWPVojlgwzv5beUgdgDVxW3r+vUSZ1yDE+34O1I5Lfoj0H4xy7zus+WAP3HjGvY2NtOFOiHbvkz
vet99azEJAe6WYNyiuRiRbzQIIqkFjoGBAMIMEkwuPKMGnsuigGg7hEDxD5f+AqKSEg7c9xkMhmB
/Bc29jXeFH/8I812qilFRn2WmGexpk1BVrjUBMNNFK7lpkQlK4DOn0c3JuIu+lT3LtWouHjAV0RW
JuqlMOIuGbTWNojnHay4j30x0SGVFldTclHIs/hNUI/tT1bCH135e9r3Voxz1ilfrRuiOruw5YlQ
A4mN5CX8f0dYlKvUK98zp5BaKGUKYhRNwC4Y0Zpn1zyEz+SUIKIuy3AFMk2FvZd44HiQ/j14WBIy
hdpBCkQfVluP8WZzUynsrurfGQ7SKa0OeV4WLpIjtCaq5GJWtj48Fu807wNaRRln3A8k3QET9gSm
AdD68rWuWQ9SwDmOc5R/uXN1t2z7sM1OOQ+USV5nTrSF9xqhAI6rHEoyiRHn0+aKC55kkcr8KHqC
18rullVHPfuFLPZCeY1265HmoO7me13qvE1LprfAyxouSinCgjEbHXCg0+GiKUAUiSFX55lzE763
lxTL1As3ZmajIrrbo3Q4ve9dz6U4Gxnyaf0CKI1maZdeQ3yrWMzXW3hhQhktM4r1h1VshFUd0ub2
DdKSN6znh5WP0u0WLk9zzqB5xt+RcxcEyW5bbf3BnyKGf13dvtdK4POM5IR+Zdqx1s1lJ2nbkILi
U/Y2+fEOHad/0a04q5T0Q1v+PpIcOUpoGuynGT2+AV8Rzf+SAq0rYwShathJQc5d/Fix/whnRGut
fMFgPEepMGhL8bzLB3ZOgkHbNGsr/r5UxqziG4LXEKAoJR9RcX2HmNvAqhlk+gqlHf6cOARkg2kh
1uYzFcPJ5cOmyvc5KGNaza0twD5gQAFQFY9qphGX01gNsnpJKJvK/fjOUH6fkdiqjWps94N+R35k
Kj3I4SP1RQdCYCLanY6LL3pMdbhjdG+1JBq+Te9btj+v4VQkpzS/26+3oWFhtG9OuAZxq9eA4SaG
qahQ0kcat3WRf+gT5fwUqUBr9qrkTZ9YJQ24+z9LUG721OX6YYycdwtlg1ZyDWrIdstKR8hOtBbh
dkGazfFrol26Hr//YNfUFSbTdkZ0KhkeZ7Dm6G0rMgNm28GvVtRhDmAdLotY2y4NiSK7dN9vs/bc
SigeSJEQIXRyGr0UeWysCcd3GaehfwW/uG+/uh+4+E3oI9nJWCPZItt/wra9/O5+SxErrv2YaIhu
Ldx0W+XqGANtShAwHD7aA4S+W6mJ+pMkonCl/KBDkUEkwvdrmjyfVDxIXq9JekT/PjG5rXDdYwGg
46bfHjV2N3rTecHr/Mj9OY1rvJhQ/P2VMDMEYcarIhBqNBWr+PgmDaNZmcRSF0GSlrE8+KeMstoM
kW6JOvlD550MSli4axFZbNgx8neKqbRwH9WhjDtza2bfAV+OEXk5AhfYFlCzVram4jlHkqv/bz97
nUA6YulMrqIYI2naCFKmeF72GPbD5ehzzL+KKSHFSLMn8/VLMe9jBaTwrdEgJSiQHCoykMFUubLZ
vyuLzaT97HXjrdFS5IsXCrQkOBI9fYy6ts8GT6aem7NJ1V6V5eMFAY95p/vy/yoHEqsdGp/d5eN6
vqLj+cBcouwjT9J/WkN8mJ/+iyoc/KVyO3RVvFa35y/KstVS1n5zyq4XYdnuvOGEpb5TQDT0sW1n
SblisRH9DsZhPT2HfJkEDb5UFL7JiRop54prmnsj2S+/XOjtye/7SIkNZhPLKnVWmB/mJcK9BmlO
uZrKE2eaK+nAdegBGhUGl2cRiwUK44nKhsyG9gV5gR977KE5cu1f/oI71ol2DU9HpbGzZVS3ZXgm
vT7ISKcuMNkPQ4Tpj98heAMBww/ajsXfiLEWSgFKDdd8BqH5zmq2fMdlUP+ismt4SICfIfCoFSey
1UBpZyJDpVZ2CsoBCy8wRh3flFITs/VEkdHYEGif/UFcNukcQIHif0ofaGW8mOn4HmbZ0mPNUDbz
uC05f6e0QW+NI+xNO7d63OBam62rQgALHg0dlxTbtD4jzMbsj7NpOif/PDwqOkeInu3y6rsiNVVi
qwF8gVkkLL+CCBMm5WtsDoMMlF13zdRt3rPgWcUzTCcWgKo5p9/NmbCteg2H8KC3e6rrwYQOS26C
ik3LriGtzq/8wTEu65XrVCQvQiNcUlmG27NjjvIqqk7yafJnh1L/1k/OjMaKSgrtMzbX6UAR5U/O
s9VOPGCcK+4ytI6KAXzX/SgVQAt/8AjvUYDynv0LeMrzJroTpYAGARJjanhiT4bePBsNdJET9gzZ
sylHlIArsSY8gmRcsJ7f4vPafMjBvS8iRRGvYodm3d5iBahF/ZQyiN+qPJUABeWoaiXzAJreVkKq
Bjlu6GVVPcF/9Kc/9SvvG11/C6NffzO4JlRrFZbSyVYPWFgbezYNlq+ZpVbLEwfdBSLKxrmuBZt+
Tj2rHTAsoFTNSr49213JNSlTozHoZnGr5Ck1G7cnyZMHXCilmk2saOj7RsdlP4qBUoHt0uzd7mu1
WvsICsyfGFxLABqOhx+0CAW6RipZfz4YYKVfMWeKV5/Y086tjHL6pU32iPWWwbiYub6h6+QYOZ/l
eaBn0L1WIFTjwROfcZs+C1snGsYmlL72cVa4FWh6A2uDmLY5ZnE3n+zXqg8ViIO7DaqF6uUe6y3L
ZAoMX1GTnRtT/aOXGJfY1OeJiwNjjH5lWW1lbAiyrzBnoCXveLkDlO/wwuhYLMnmJQzWW7cSo+gW
exfjXWksXJ92ZBd4g6uqy5tvm2XHwN7ewRoCb93nuiINDmlnWj63uk6vAYG6tYlAoZia5aD6ELfJ
PHcMwHpRMKVbjnqgyas4QfRiMksZj9Qh49GDEZJ+BPBgaqFlHKaZkEeMEspZm5M4yDrpSaRXVx1a
63o+oa/FR4g7vP2Ons4+fiiX1dUgm8ZaJUzojQcQoe8LnN8F7rd82VHyhhIllC0yUbI4EhCmlGyj
Amlb0n3WNVkRFyzwvnySbP8GyoHXAv0jByEaxgiquNLqI+e3nVpreV904KVYlfLTblurp1lAmP4e
BnuuqGAtqVyQmV4avyt980xohSKZS4HpUTO8hQllyMOJfotVtQ4jgOAI20nnQKrkFRKSFTNl3f4i
5eQd2AmLkJsD+yXBHQwSJNMi634FACjoYbiud7VVJQoZtzUb8NuL0boXIu3HN+cYPYFcaiksYPQj
3x9YVv4ncx6GrqqhdYlOjaR8uJjoqWQPBOjlc2/IuX1lJfVf/ms3oyhv02H0gWkk9StwotFF0y0o
xcFu5QPW5Spwln6YeXYQ223uV8EA516M/4mYzYc+BOKl6/8JEzFIq5cwUbi1H8Ta9zjSDd2zceUS
Gjd46KxxxkmJEXkPrK6Kz/A2yjoHFlw8fan9Bn2oPu+oVspDrQFZBJbeVIVEy/DugF5m4xVsfMeS
/SU3ugb+gOmzeYl6E1I7D7/a/4pfPhAdRko2F5/BJm7Qnn0yi4PJnrFerczLuRvsdTeM4ll+Pqby
9SA+EHi1mFjqR4QpgUWJHcgf5AdNCTifaMXjjPSXfWxrzkQGjoz8feb/kKmqDM244RzyZe+nfOCs
bS+WHfHlJtmrFcPBPg9JL6vAVWyTmPU/qJQ4m02FVYGuiLatmSxnyaOzP21Kl6D1yeRTCtFOOPQp
ZPP33jZWdW0vVD7d0/X62WxQyKqS2f5367I4T/h455EOTKjsK/1QtnoXDgF81/I0ZIbkqYxTu6o5
f6szSWDBAKfxegmLMbdrgoEUVPT4jQESMqhtTpAIZs9XctDqaYMgN1BuUaDGrfDXDG61nfl/ncGV
dl6tvSNe/sAzT9IwKmjd5998dIZsNUoIQUpVKxHyVml0zTKJJIihVlBYdtU9w2/EOD8DGdpVwdV+
zPLd+cpF4h5YaZi1eFM67E6DxieG/3IBkGz6KNTxgmKp87acVQVK3KKLHJ3lUEtS9q5gqWRl8VXk
zYD6O3gVBlpjaa/xnDqXNd9JjTipAYlLYfL2S0sHEPUPqg55IRGoakK+vvnA27Rjs1DxlfhCtlQN
F+ALIcszAbVyR1sFFCuDMSNQJy4JUu+p/kJgU2Z+vRruKbb3rtbGy+56LzFrETGS7/nNbiUfDhZK
+wPZpiwXUMTT9azeCADWywGp+XAs4RztjQdz4H8hJSepZjlYEW8GcbGBsp16M3yQVSnaEqiQf4XW
ZYHZ7Jar6jq2iDpilyglqcTWMJSDGI0XDVC35qx0x+iNtFb9mFxiuol+y/PhR7RZMjVnBuqmmBrw
BsMwhvSmFF9WO85MW4zqSAauHOK/7Uq/B9rUyWaCPrYT9WAO8jSRuXE3rD8wo/b2aNGHU+kTRyE9
TyMJDJuHE4eeWrQHICdARuLqFBjzoXz1nNDvmQdfUfiBg7pYe/kXSK5fhYQNu+cy0cpMQHf6UfSk
ko6ZBzuIlCJszVMjFoIBFHwU4ClZkn/zobRJN0y2MPS3mqIiY+wlVN1UGxm4KRWjRz6Md0OkJ0bD
GTczV3QsV+K8TYx+CA9H3Hp390zDAm1q0IWb1mOFiFv25TDspafGtFZ9zELW8EX+6UPWui+d1DAZ
gV2KQ/MPMLFZZ1x6FtHpKay7VkFsAtWP4OhSDKHrSBQMN48TFKQYwlh2mRNypenj4LOPKNinatAn
r+GHOuO4D92h6FzZLBflyCOxzl4Lim63GXWgXsTv2VLk1hULGYJX4r8HSLgcUil91DL2Ng44q/hR
TeVKRJxbsQcdi3rSVN2QsnrYyI7S6u2nvJdy6wKZySxWbDA49uRWw5MLvNBo77AjoMdyNuXPBjZm
9UFBfGrZQyfbvBNXigl+ewFHaEDV/DB/O5XKYTdKaBKh3FPv4g6xFtF3/SMps4SSWsQ9D5tIgUmE
qK35p8sJ2dVZxixKgLW2QAVJROSi/Ptn/c8ekYO3YDSKsdjjz30kRQDHFj20VS80IWqRMKl8t1Ou
ZxntK+BqB08UC4BHANnkmbmdTY5mSDcu9BgHi+9u1zavWje+xOHQP1tPXHUWzny0DPpNVajp7AHf
OQqjb8IJTmjha/ymc2meSas0EJ9M7W6yXQAQUJY/RDbQZgfXlgKATOwyNt1GXZHjDUv/8KSXTB5z
3SNB9AvZhX5JE2sve4w5DXijGdOvWuev1FWsM1XZNeEPh6XE0fxb0ypx+co7dQ==
`protect end_protected

