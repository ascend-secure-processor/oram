
	parameter					IVEntropyWidth =	64,
	           					AESWidth =			128;