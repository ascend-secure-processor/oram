

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q0JRSBI6K/erst4ec7E1gBkk/sWBoLMapXFfn+qmQF7kx1qpDSZ8VnrlcR+hMW8ziQC0Kupa0wcW
nfmRHMd3cA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eooqCjb0IA78gqMw6qB1kV6DmvBfEGYJw+6IkPeKaXbNlhvCOpPNqk6EqIAF+yWOXbq09g+w/OH2
p3xrIyEvCEjtc4YaKXZDQQCQF+hgL5wOi34WFFLE18XPsOzJQvLmN5XcafupAsBnJ1sbC5eXYxdO
sykJOcMKSYqe7yHKcIM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gxcn1XvhWV/wy5gu2OwtEJF2KTfIAFGSvvgZH0bIEWleYZilZnyuiWKrn+K0Tl3an1fzyEiUBZdU
U3RISdexp9IWLgzy1CM3nXrX4B3+0IeXT6ilQBcY0UVkebxKUak+Y/V6Ux4s6nOhZuqPm4TRQpcs
3CuvH4/4FT8DUBkQjA5SvlRx+KxXgGeZFpRBbxXD5jcaIpBCIZl1jtKTXMXL/CFDr/tEdlLsQ2+q
ZIGkgiNFywU35oWgZmpj947Pt5JKsGVNlf7qRkKpXptmUa03sLPUsCwTjKx0xgYIt30T4YLQKqdM
VNAjd+McXBWjQAVzvQrw5LjbrEvI/nmU7Pedfw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O0ZNqL/UKP82D4/Xmt1WR8Rknfsk+l0wFaq01Qo1Qa7BJuS4IsrkV8RAOp3i4qtiWvOKL/B08XYG
CJXvbFguQPKAZBN/xFUKhDPmxBRZNqtjJfS4IMrq5CBmp9ue6SEMCeJoFbRiqQ3iT9nDtENsb1Sl
1i0ki3aW7xPBgURIkBQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VRxrxSeeLTidTIuLNKQufFOocP+TKsQWZYkUG7bpZtRcWH/9FuJ4VwolbWtONsJSbqrFxsDvjvkh
hf4IASyHbwdXytTTHOEZAw64mQ30FiYPpbDzjGnkD6DTNvHXVvCZby30FTMoq1KeUsCg5I4WODZx
D9eLXSFCBSwRE/LI6yWsZL+TSCkQzNn3MdjVyunsxom1s5kSp4pZ+AgAtY/cHk+qobuFHJUBMC0S
+fJzj49HCo8pD3o4t8Ll4t3uME9OxUdoVVg38zv0hsT2cpZ3eDmaWNgszDL6EzSgxgI+d3ky77ke
XGft3AOiWWKZGiS+7Cwq3JETr/4KlefHXaeqpA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
j3gH9C1D2cmGQMucvePkbHFnyOZgk7tSkPPIUgU05tL9FBDQsc2zDmNs/VqNNS3rjInS664cVS/b
MApXSRmwbMqlScgsWlwiEWj73h5cDgOX6s/TCX2A+gcwej1GbzTYgtjl7nYHiWaC+eERbgAAZZAW
IyjrtcG0IOf+SegjlAIvtJsB1Aa59QLl62pe4o039BB42Soxsm/bl3mx+NSnP4cEfVeIxaIg2QT4
zJr1S2wCkTyUQFUkBCVqBHBmI+sTi09QkbiqCxO4GKt4p8avwYTkvUYqaN+zEkXd0YuSahawXQgS
gT6okIJsDHb1Kvkk/1yZP5PgZtryw1cj4xO9MAw0ZTtmJYtEJXbHwaHymDutbYTzDUjGAdCKpIyu
LMvNuMbYLCB7oKbrF4iuYugUqYoPxbICTFQ5LlNQ/1UcSxd4UPQTRSzHgEo1/3OEV6i4KlLHLEud
rwO8Pk9znIKLINInfKLik5f7b4zPvdw2FQsnLgOTUpUWGOQsAUGTzJMbKOWwrwkMUeT6scyLSSBd
ojvxoANwn4xKxDpmeQee/eCFtemiZAUjjKorwvCF7rK3McmnOQDsL0HAER2gCc8vp4Zv9HOKtWkz
Mm3CuCbs8S5zHG6uCPwjQuSw7yXFuMEcautaquFUCdbvGTauSQ8vlG8f1dL5U8pPGYtGhVHK7LIe
9osNbOn8C1gdjmG7QRLbbtgCpq2FvMWk88gAb+3c+qPHGpx4jFlul3mRb5bgi4EfCgnB6/VzvUOy
RHFrIdRHY3oeOD8i66Iia/kuH0JNQbTtBfgj0uA2odzk7MoYLb4Q8TuW6N3FFKHy2emfwA5EAoHC
2h1VWYlkFypT3fkusWHuAqqPJ51/7DrD6/hVmfLzzwFoG5auGE/CJqVBo0Pfm9uIjzM028t/ea+2
dwPpO9IgV64HVr3f6PJsn1NxPOokPQTQLNxm0/foekRm40pOC3/OYkXn6h9fBIBgeFyuddWpRr1v
y0PlutbFZGdG1VkLOlhwKDtD+8jkpvqx1lgWhJsgQHiGEbR44qS1yEv0oilzOzZYp4GA9nXRymjB
qpPJp/7A1nPBDvr7IlgzTSKy//hBqeKi/g+VfQO9Nnq919qNaxSIcReB/5xUc2xV3N/0sukxB+sk
2t7bRhIOhlmXyT9fG/EIKlrTFefcrOkOFZK6EQNxIxNTZTroWcOY3tv+1Shdv7GD/HrsVS2F0B/Z
c6naH4ww7JDHUeMIy0E7mYZA605SciIhEWgHWUO+SIF4MGUWmlCUZnJ7YK9os7I4l7qPv+wUcCKl
BPKs2o7gpu+4lHl0W9M+qkeXxBYq1q6LSd3wLvt56/3GGlYrRM3DtfQMcw8F0skDvuOyFOa5jcTx
gjLd22mqZGUvOjMWIgbzVO43x0JNuhd3+tTheTiKi0PCqh7aCj2jVwLkd06TIzYzAYMPdNVChE9b
zpJI0ZQ3Wfsz4Z0SsEo+v+ZK1e0aSPQO9iZIkZRIchI769YLGcgh350b8+RAa1PwbpCdqn9Vh4Cn
EtlresgauvzuJGmzQMyd5XUhWDk4sH9En1Zuk30xQ89DdGDeu1fDjKswNT140WBh3hreBjflEzT2
NrOXJ/f+WdDmJJvJD7QJ6lYg3qCPEQ2rvNZfPDjTtKV9SXqDrE27grtSNs/N+9zGYi5r7+WMfwuV
0axX5GFEJszBCf9d04nEUh/gi7QdQCMybgABH9r9NDp1Y+iEwARcTFoqNAw6KWqCpzy86SUUZp/v
ZnqZY2WoK9K1x0ZKJRQsguoP4rLlYc4Byces1QZW31waFNJhweNTtjQ0ZmcGtjq/UaYykJCZyS0P
OYlPSbs/XeU6mcCoDON32FARCCqo0NOidPQ9N3BsFiijIES0+ufDD3ekycueHsxcJ1XDC99bPcbF
XgptpO4xoKyj1s4pi3rrdso5BqD1Yav4ZnmRq1507uVnj8bfmUZkVMGzQUJz57nuNRKxLV9HKP7D
Bq0UQ3foNSVp4JtS5CosEo8A+JqYRUOEguWADTh/0eQ8rpXsqKRauaPrbustY+WUUJHnPIE0DM0G
gto65QxwWWw2cUQnoHp6YDPw4plVG07Y9xANwiCf5B7JAIxPBL+mLfvkkMpG++J7vMFDZZFU5296
CLGBWq94VHcYWMphGPXqDKexvIrv0MW9l9U194BFa7SiBbi4RfvCWgqPNqH530nt0A4Ve896Q/8w
VuxwDhNLcok851t8C44ENKFFBgPHIRlSFRRssTILfvUbecMk3AS6B49pKmfi44pMsVemBpbBvewq
9qpyaRlxV3fnbOs7Xvh1+T7Rj8h56A2DlYPAqk3sAlRtOMsdjEEG847ES457UKIijyMk7gKSAgM+
a/3cJmE1mavAdCc+0mkWyVVs6MrxCHkeq0Qs82z0VwNXHNbTwyW4zgNbhONhJ0/OJq6myDZ0Vh03
L7snbEnWGa80tzgETVi8AdS3tWhm46tyESgFnWtBeaMGkeaUZIowu1Kdisoj8L/2SJjyawWYh9cj
lgviS5Qc3kmCy5ROm/jUesc8EYSSc3WbJ/X9tBO7mvgg8grc4yDlMZPbvtnDZJFyNrqRnxbXJlpl
Yei/VrN7g8CVxPy1xXhTL7s1f/bDCRpB/xaVUKWvzoM0UP7qT+8MRKSuTKS1VprWlkHP8/bat9pV
/pmL+lligrEljdyKy8kwildzrf+DkgbZu9hLktnLqMk1yQS8cZ++xIAaqMhRn9/mq39kUKfFwrgg
rYfQEhMv4pAsaHZJW3QKmCEfyhLspAynsQC4vrdS/Rm0xmfIGJQtCUgWGY8Ql+4grFZesMI25nrG
UBgUqqXXZMp6SV9OVjpLzzybxhBMCoLbEMGZHb071ba5ZcuXs4Lkf2BuL6fv+AdsmvPSPY6VIwCX
sfsJWoumhR9A6ZYg3qfyTCNAmgGvTFfXXTrHgk6GZjBtZV6JS1jRD1hfIiEn1G8f0k0kYgVUQ2Jx
iZzd1FADOAcDonITdfa1wkLOUuEkkC9n5GLImf9gL5xrqN9bl1t3Y5QJcs2prg83qr+hjMLOkp1t
vzQUxQmGR8cyKHncTIWlvEHPTpBUATx743eN879mu0yNlbRp/RdEhdSLzB7SGeNiPZnSsX8M1XKk
OSLqarrTnO0HOA6Pj12oXfrQw6t+bYL/WcvDXAgrrXBWV+yZK2VnRrqsRp+ivVy6RtzhIOysPtS4
jQ6UI5oeERzvbaW7e+oQikFWQh6f2Yi+91yOmeNGKtE+H5YsCGVDcIWhFP9xfwPDNE2u3MwcqPoj
BuIYFfjU6ysmRvC7ks8r2N3rL6SJBAp1A51Hsk3Uj5Ur+2OlKS5Bd6gTXYTpQW4Qr5kVrjBUkupT
NRWVE52rdNZK7fvGHBW4ylsTifko8ZiJnQpV6sdrPwWxN6VO/bVWPOUuIj7WXaYpcYQy3r7znNSb
j9whABBHRB70LeB2dlrnWXILbu+VOa6GFQEPV9JGzo/Iiq3egQgKOW5ayQzd76qkc1XAv4MqWVI1
+UQ6zYuzAPzo0IyoXO76ewf1GmtpuK2HKZdGx1/qvccqshA3njK70OBuj2RI+VUXyBu7WDFMWtph
JS9STtfJwSVVNaAtoa+9w53pI4sC0TPWPCXhzq6EJR+b02ErYJPdsX/R1eHLbx0+OzsSd2q4swh+
/UATxkhuOhE/PdR5diQ0smr5rirlJp+W8VAMAERvELjheVV/V5b5fDZBtGawSaT+k53p5SLvCfmR
an2JPbj+m4CuGgX4gM5hgHa9M2T7HrzIZrn1TxwQaZfsXfsj4rrGJhTc5qNBCUGL/Yq4EKB34Q8h
jm2Gfu/TXjutcJTjux3K5O4k3YcuCVne6AsUU/8Qzp6iEcLqSUGHRJ6x+DEnLs2/oprwkAszDYuS
xm696pXweXDKgmD8P0cxv3LAAVLnrR6r3RPdlZ/M92a2FVmjALqk6HAeleRUz3MOp0iucj+y/gHN
whL56eop/yZwYAt/PYTWZ0dbmlSpQmdn3OFFY4zZRiEiF7jXawWeao3Mzx86Huf7OpZMTo/2WkzQ
hrfUV1c/BuEmVtj1bIY4OIKnQnN0FYgiZM61irkmzLJQ5sdowytex6Tw3HO4OAAnACN+i9w3WJt6
mdZpT1uoN8XwcVYNGtxMKXeIkvN1sFj7U6SbyQ9vGcChCeYwKL9uNumDmhOKXxLZ02v4VYzO6mVK
fvF82nmwcObijMMC7l8tXKDPJSvmDb+jqnQEdBX/ijeoCvAqc8OdPq1I99BPifBRNof7j+fWbQ3C
MkmRVl/9Mzj9QCcHyeHyQ4bHFPIeasQB6PRxjkZcImAl9TFPKANKxa30V/iUfhBNR7905w6PNlJS
WOwOF3tIHngzlwH4OO4ziPk1eKj0XoZdJwdCxcIld/60hPjBFq28ZCFWlsJy19Z2ljjxuAPQJqtc
RS4lH8T3slsp2F8x/Jr7rDa9zc2Qq41ptK/XwLQPI6fS6LFY6XQLLmc47kPXQxiOYSLK88yivFSf
IRHfkKqyHkaP8IvP6oS2/T4E8aBx5jz5LYnUh6VTbPfyE3ym3rpwUA+1IaPcQMCX+Qp7KzC6AT10
p46SuAbmsIDswrhuAOzndKY0ywWe4UiZoE8Ey3+Mf/efUWisSsCJqsy0k4arSo+inC+tCa4omDJw
BzouNIApHac7WAvtEf269vKPsM0iwHtCobPtZIB9ztEGuxQ+NcV2TArMksB8zr1Fr+AeeatXDanl
2SZ7WSs5a9AX/abFZCVtyhTlwqHNSSuErUk7r56gNQmXAHJ4QWrfnXHhpBHRrfO/83LacAIGtUIp
6JHLFSPuVsZymavumCqzvunVDWHz9t/IfAj3tBBOwvVLq9zDpLwviYAGN5EHVFP3S4JO+sZnna69
My+0q+om/uJ876J0VCjlnVF3sxPK3DRMbhYFjFqch6k4bCVQpeMkvayHzqhRocBSDMO5L/cEwgcn
YD8XpUwH5JmnOla/64hwy1LA3gI0G4u6aERerc8I2sRhQg6YYxLxfwVVdDFLtClQS7JT4OMJdUnI
yWrwt794ViMQxt4LlBBno0ai8SuBIRG5SCN4fYl9pO7pg7U4YiPYbxWA8G10f3CHwg8Vh0rMiUhM
EYEJUhDQ0RjHr9QENs4y8OLZAGrezysWkxgYnYDB6Hiw2RpS+B6WIHx6aK4u8KHiP8hwA6ceCwtE
+53l70wBT3g6+V0HUpaB3j0doJ7w7V33oh9hGRk7PpkkYIpn/IvgTb/vse54uukM3AP5OjQ5Gdt/
SV+WF4YNms1/hT/XdHQbkmPe2v/Qw4XZsEpPbWmJBc3CWYcthBE5eIvH7TwIvMbAMBo6kaSP8MW+
S4xepZo8GQtF2aKzGMF0e1gS48RJ0p/Q4FeS7WPEPU1UpXwOqh57yXeao+ztnOGWVg10MzjE22qo
nRVK/DKtMxeLvjncz3YZLWyIrVX88whNcbrfZhL88sEiYdaIFAGdRHGWWVl5v0/41IKLEaT02XCM
ZxDzWBQBa4+jiYusy3giuFYwF1361w9unSOeN7I20P0R/sqTDuq91syMsgqnNhWV8a9h0FqxoR2g
DfjwHaAK7v377yT2Clw6prdJqI7TwIey2wu2n3pKOyhOw5CLcJ0vg3ugJKBBedxCeRS2hz6kGKMu
/lAzX8rbq4ept10H5E6G3zluOLKrSVAcu+p9V26afo4veV1EDLee0APus093zFydPTob68fU5R48
UG1MAdpLzWZFjm7kxUnDsTilZQUuHJ6bi9MXyWvFJeYV4+dfFqmG++X+xNkEoM+INmwiCM5ahMlW
lXldRBbAmdtYDv/wAf6nGwttLJMUBV7qB2Ojxv+/3pACg08212iirmqy/ipbN8cxcfAkjwvFINoi
ijw8jB4bgZ9TXc+625C5MQNTu8J8ZW+1xIw4hJjTK5u6qny0/lUiaZLNDtehn7RpQagczR74tjfW
Pc7z5yGeWfVttGR0yiyh8K1SbTBst3ntuC/wmhQnpD1baNSVocOBLxb0qB+SEfusgPWX843vYJWo
iN93LAAjTv9ZGYlYASeU03JRiEHKyV6BYd5Wz7WrAS613TFfKVDSTlu+HTHy6W5sn9xMt42W6ey3
7WfolNbv5q57iEcjPMQE6x2SIna+W8fFkaTpzJtp0ipShT5N7wtNoWHyYK1SCQyBd2y9u3bNd2JK
jLVUTGTe/JbcqbjjWIj8xiQ7TUITPzl3nkP/IkhjRkWtJUR+LqOoKTIXK0YJ3BzZShwi6/659U/n
BpecITJ1jSACTvKDdJnToCpS465xFCBKtNqxqxvOJk3KNDv99ez7SIQAAO10ydGOARnygloGjwXF
hi6WhOtbxbTCiPfkbFXPNcgoZxDVb33EkwuRCGM9ndUzCi8O8IMROlTAto/Ni2ivNS+bNHBM/nTm
z7OjsZl+c6xDeoYYrDfMG6OhmGiweJnzpzCJ1KV5ja9+f9iv09snhyAUF81Pmq9MIgvotFw+hdz2
qwH0KPTT+lWv6PCji075TqlJGE+LwyOVxvHb92SSNjyL5zbSb7wV2n30aQpaRR4s+PiAWXypwIag
7b+sCCFaYrmdnhXe+on6FiyfJOh/qCuG78BLYtPgjilEtQBTX2ABmbqrUqn8hNfZJ3fAjRBMz76I
maQXkX936s9OVTOqidXn26I7Rr/5r2T7E/rmjuW68eZbLnQEWeLxWqyrrmIDuq3mDqmDxr/BSj5A
wValXA6d8JGEqVp+dUK8ycineeMcWEy6dhlPiihOjGvoZnunoyeH5lIDIoPA9/Hxu/KIfeWqRP+Z
ckBrKBcbjE6NNc0L75Bjk5D+ccTmNaJHSEkrhx5dDcFCfIwTDOPWz/BM0SXzrdWJNHNkznu7PT5I
I99aisy57dGDsDKH5zvcGVBgpBUY8JDMqgRyEpHwFH1SFCg2/Ws+zBfOeqwSsRHHX6jacU9g3QDZ
Bv85CiqhRZxukMXbK8fv5f1+iR7qmoxkm50s2ZmzsJ3m0Eih2MDgdp0w6W8jkTRMOILvV8mhF62/
KFw89Kbgi0nBDNGg5gXTdRu9gqpILuCssyY9QW4V4W1w1i2kKE2OW8lCaGykNaWkJcle9wINO3rE
dVVwQmM4jvC9RHNkfr6HA1rnDT21NyaagwL1Fa9lr4+Pj2/bD4kuQz+JFdMpXmI6C4td1PWSZ39R
I5L/PzP3SvnINMJolJN4eTNhM9I0T+glpT558xD8anJ3Bf7tSUglCgx0LxNWDr3msS7c206puxaD
aLDzuqLxQhgb4v6iKRwxUHkeuYI5v64Idi0W4a9lCKkjWWBslzE/4ZKCeYlUGjS9OqPq70gpkvge
ojcojhFlTEKUx2hjkjhM1UOnKoQCRo3un5eqN9hzTe8B6Zc193WALg4+i2POTBgXtYdn3WhR6kcn
qEVSDr5V1qTsJvp38u5JlqtGAgeotw4uXVky479iYuVHwmPwSEisIT/e+I3CgjTJbVlVlYQcmo4a
by3xEj0FH4zJjsvaWFsI9p0XHv4WKsZOHujgTmd/6sm5AewLOLeSxK6+KzGdPsbUn6X0b2RSEPqd
eWhxf00grBgYsT3kiio3u0kwn60z740aKRe0jo6GurfwsKMz3HA7p3+REzO+MPicZkNeV1e65ADw
io/vZ/NysqhdB2/S2o344hmg3kgGLMe06L1EjfmXqU1y8XYXuU5T5TeM8PfTMw3AaniHJ89U/N7u
/nD6yS92aabyqSY953Kf0MDhgydjeBVcRzzTOhSnH4fTUonx87fEPxiJ9sc0i3SwGEd6Y/dm7Dhv
qrz/WKvW4afKHXOss1rzDqR50k4dgZSjddj1hPpCTM5JwlTGRbrkTiowROd6Kws8q2RXYdbj/siG
D2DuObN+nVs0zW1eJz7MvuX0L67Ic7/uj5Bx5oE2qEMlnkq2uyn/MyIMDJodGa5CQdQQapB8wHyE
aXK46KtvoRGWqKjfs/dgd8a1GnsSuFqkx0tHw8SDOPDQug89iyCqfgtk7dGLIz4NTHr9GxuIB5Cw
E4ndEuqguTx0GUz8rOzI
`protect end_protected

