

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kIka9mpyIubhf4qBEBTWska8iHrcwPvUc3LcKgedWTdZkIPt7vIgBgM2KxGsncuzwrBngAYEBOpT
Yx77dXnbeA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CSBztcRtXBBOozyNVzGxbXoojp2/jM+V7FCgAJzmDxmf+ufv0IZWYU2auz6/7y3UMC1sto+efY36
QkeRz48Zci2luoPcnouEYaP+ZDsQVDUdSgrqKrw3gQJeyFZG3BrUDsmtEMqe8yOqQaaiX63z/ZTs
H9ae6469M9xvgappEok=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eDIT38GMyTLbqQATmvqfMGn6RQHaiiClKg3VSBSPk5lQEHFzT2WQa8vjuelAOuhwLZ39bHNGtac4
rfv9Mb7RVEA7of/3oXv+XzDWm+MRhImKBOzTz0lBYzt7TaxvC+jKcxawC6tFh9N961ITpMeMk0ar
afTGY5qmsZNYudXYkTrtqTOz37A8Xl2PB+iZp3PIv7/wi1iMKgQVaBGP8clYESZcJRKdcqRQyGIO
T883JztBKa2yBJc/LOg+Wh1B2Dskb8h/cNqqLrAUEqugv3Q+ZwXMzLkOB73Zv+9C65ih7mGL3fFb
0FNymyETHPxnIOYvaytGtdvOuppRkkqCovOW/g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BoiVrQrmul8h3Oxra+sFllH3TaTbbcW+J2lZ/qO+K7lHM+An6iMsQ3dVJRysGLRDmNhFGk/iAGzT
kvL6q5azf8tLprZFA14sB0I33ZFuwJhjJSISCPl/fldjlfFlvSUlncrtpHTDUyZXf7mOJoVVpTZO
J9HSO25jgG1htFNGBwU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XviGemZDYO9m7KSPR4B6Gjei2d0jUXKAIaO/c3aAFaB1xle6Ypm/1wGYPE0kGIHvgD2cLnjZs9sn
i4TxhKl7oELTwdGfDz1QsxiJJkgNx4ybUFxHol+GGyGq0IIlYp2Eo8RS2b9DAGHiJougWI0QTQeY
d5oadIETetIZ4RM6pwh25Azu5eIvBT0vZCMhTMvBDVqy3OHCmrzdaOQD4KxfYTZACT+w+HueLfy9
RRTEh+an9axvVAiU9s2JKGTWpmMl5fWUjvM6BWE4tgPZWdLsqfzqC40Z4iufJbvjYKV/aI4YMvQo
/rcBZeHW4/wGDhAtxFSzn/1XEt7L2HtDX9O8Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11632)
`protect data_block
uhmVvxTMBFFTYtCLEh2+IeMWwBVjL5063aAvYDnxQCLXxBKpwHm9kmzhOEUdPOb1gvC+OnobW29P
IFDGiAW+Wa/kQNmzXI6e2hOktWZiH3Mzz6OPbcGCRhDSFVq4SfXicjSZZK81PDITlwuHee3hz0mk
CHaH5cJ1pcluy5aMxj1MpKcpDvUlV6DFvSV6xfsAwfo7h7fHfdy/81cj3dX7+fxbKScrN6UqEkT5
NV2u0y3+VufhfadW69vQpW1WHcvP3LvwhQV/wk0bX31wSTuhnaWmiSPxGzECzxH6c0YMTOGb+aE9
ukZvE7LaY0ZmaQDSqGsZw77xHps3Xa9dXp7CWFZ+tNJIBmc5Kw7Rx0SBKSxGur8ZbhFlZAy2vQC7
kE8FmjjzX2rf2Qe/ckHcSziczGxPqRFsqD97H5jQAOO0fri38OGDMviM1+PGysYosLlY6eAMwGP9
6Xder0PXdoxOFBz1QLwVCd9E3476OKljscwNBpsx5MgB5lorzIv8iZJ7EXQzcqijJ62BjskQvw5Z
sDoTIc84ZKNyvc7W0z8M7ZUPba7F6P0OlLEMVW8Znu3fcI96Zg8QTe+NWI90b2U+GLEy+2n+LA6n
hqO9cSIP987jBnNLyIRxzWg9umLKoiLOaWF8+TNcH8JbX7MKoRf5hKwm3fZJFIYjnLbvT8bZhDv7
6YkvyMycWItPA+1esbEgy/JaJkS8e3r3FjUoWCagN8VuisYFRD2j0ic6mrLhIcNWChpyDeh3KFdf
jnB2AHKRZyB96LxTZTfBSNuHaMPY8ciDZzZ/kai6tNbED1/sksXr31EFeQ8jeSDlVGxR/S/0Jj9b
lQ+e38DwiGfOzsloZNAQ1DIfCyiFtkJeQOJGGk06xqsdfu1GNriI3fhFPBSr/svY73kh617HxeM5
xo149+a3jQupHv6MiF7Ka25QWia/CnfEbFBvJ9b+s6LdIAfHAteEbQa87fsULOdae43m6K6z6Xgq
6O6u9yMnxczPBFX4PlxIxEctWlVGGVS3y1vAzWOQqYynpgs8QxxUSuV1IWsyRKoP59vpks94tcby
B+G4eYhuW9rPEF1k0WcUggOmM0d1wtaN6ROissHxvmL8Cw14rslMDBwHliZQ5BkuR7REcsnWuYem
6nnzKYiXRIt5RmjV6/4T70jEL3DtOaIrL0X0iUTU71AXlRARfMkRlP+oQ7uPFMyH8WbRxj7IYDao
THjSVbnOlXyWjrGqruE5JSC1RPRZ86u+N1RUcKbD8qta0dM1O/bEGksGETacIVQTCxDGl6i5mubp
WJzp493sMf/wwEMiAedSsK6mhct4z+79sAIxFEV+bPDOTclvyh3ibcXgJuutLfbOi+C4EUt3inF4
TcE7d9Nw4wjIKiTc+MXumeQO+aCqaOlBdp+d85Fah6FwPeDqLfpkVav83JWUebtTU+BWe1RtgJyp
4sKkEk0JzMyvIS4txTkfvyiC0IxobUnKUinXh0c8CpRjqMvh/wvlRsbtNLEZva+sJ0/4Pe6F1it6
GZWP+/5CtiA+3+2TxnF3KLa6Tvf9u92nJ9hMRYa7z3S0v71dUjt1z44hMOrBa2xwvfii+DUwmBEY
or9iosBC1fFTzEtM9QBV5+KtbGcmG+7ngvoVgw3IvaiUeZAwHTVU5vaxFa2SOS8Wl6tauOV2Z7LX
4DudUWke5LrEE/ZEh6TKsaMjlmGUWPCCQXSbhhUZXDwi9tpRnhtKZPLzHA92B7ecus79mvGB/Mi7
x+cQszDoiEnWFdIV8Yxsjincy8/eT/qvdYEO4Mno0+mU0rBliKTrhzbLq68rZciTuJ5uWdDGZyAr
duDmHr/H1P2LKjGaHoLWIbhhkIZbJdG58aP4RZKfpx83YiuzGW4SeveJ7SyKnSb4AsJCNbXz1yWa
f7vV9DK2hR0+QZWf1m2iXb+LiFq03j0EbmkPdi/LrJdSp/44DP3ubHV4Zy/ZlUGyVg7ThCw5UcMA
o83Iv3ROBLUGIm9/UMUEkz/o+hy3HPEVz+2bZ/I+/GdBGLP4iaEBdvFa8yM1Z83kBYnuiygCXg8I
jhkWcpqnzi1AE+P0GN3ago9mPUkPYo5m1kXZjNswGDdCd389pBMBYDBYektqrGP00WdHAnBUsYfl
XScBzP7g/EmpUF+yPvivI3gsqlJoKT6kvRLhmmGWPkYl1S/zqz7QP8s3bn8ChTaT6jeOPiweE/Co
+sNgfExGLWAGC0QbiZoq6fxs8AvE/+PPVnYmEqed3Vi0IZ5efqL4Dx8/GG2yufQroFp47b6bm4Ew
/QNNqRfWflA9J1ZMowllyKLXwNuvt6jkUQlehw1OgMowba4qq4ecTk+WdKQSehfS72UFqOqPchKB
mgN1KQChSTGjqENX3E7ZC8+Wr3bbPMkc4xx6XAMinxMw4Snu6WaApc23EuXl/yMM+alYvUSJ0EZC
ZlFaw0XFTFVbBmwFJGDpmnTVQCpmm7l6JN7AKWx1LSdBo5Myy1VsV0BffcD6/ZgMaOHQmBt4/fDu
DQ0TWuTfGiux2lZXOuDec9lg2yYNlsCcJGr3iAza9REvKyqI6VljZphp2GK4UIFP+Jsbb5M0F9Yg
LaKe+WDlyb49Vf5mJ68M+FHsd/VL9Qgxen+tpl32TZMzPhA/cRqTnTHIr4/aE07Q6uhYKC4LGZcr
DpaT4mj+pHymT6mrrXDprGbI+P4S+/4TtEGZtZ9zAa9K2i8WkNFGX0BdpssQ5xQflF6AfodnsRc2
JaFcxBzDI5rIm/bpVIuwvTnRyU3VGQeMCDzEuYNwfC5bec2mSYhD8qjXAvS3+TzfQAda+6tyqYoQ
p/d1a2LcGKDyTfLZkb3YOokYnfRdOhqsh3AQRf2kLs3oS0xCBRZRwV4pV17UqGBIcR/ebf1NXWMg
3vxv15X261SXAQa/5qweZG5TjnyX3nuUexBRc55onvw5vHhBDAwSiT99DnZM2Ankwq7mcSZvdJpQ
zRX1MU3aeKHEUQn73g3hJCrq7D26itT7gJjnbMDu9lY3toQ9Hv5Ybmb+eUQgrWQLuK1mBLu0KeCk
wgAtXXLDawNZmGcTXSYUszoPiwxMUryFfeBWfeFmK774rrB5qirAZJO4AGX4XQenGA0Krfqo6jM1
L8iqvlPAxJEPy8ICJ35vUsDymoMYWdRaTKbDSfoLyBuYFrsWD8gq4K6BrlBkXuxICoS6sXya5gCc
Qn4dhVPxszev+6nqMFZ7XZmXIFTzA+j6U1zfvPe42zbUCpSPCdanHRC3pgz1AFmdjBfUbJ9fH+7l
B8Ilo7ELetBH586kSoc6zqjV8eimVafNLbTasFh0zIWD/GK8dQznfF+0y+WoHticcKalT/coAq3Y
Faoi5iHPatJs8I1e86RQdYKGH11Oknz3UpaEahHahlh4859wOdEg2BnOFoYM6V8J2T2qt4aqfiUu
4a+rlDQbTwBALk8AWLLGoyy8M60WuYWx7dz7L17i//lrncgFvvW+t719rRBUQv7lLYkBnmlAISsn
liPUSUiXBl7x9vnAp2qTymWifMIelWn2N/X+7JUJ/6hC0rG53uZqc0Hxdxh6RSlJW/fTzqY8EVyH
4XVQxwl9O0TIKzhUUtvZb/dbgd3FoW5XDyMvYIUAcDbRsK3BAZJ4Fzne5UnIbb9lKipQ5YgR20x5
4jppmAt1fxmrLTAntsYs+S3w6vMt6RRxJthV+IiXxiCMMu4sa76oHUMZQV/LZDzsc97l1Ef0POVg
6VjucDz8iqNUTy+SQaNSfGr+9izHth6R35Ym+dWmdxZLcFUmDYoht9sPyBJf09P7MoXXbXIVJ+kc
tZ0fj8cMiF+5FFkrO8TV+v9wfr8bCoEk1+p8VHhsM90C4bi5PwLVCDYW6df5k/mRno1CvGjSWXFq
TBAaWwKjs9jaQmWSRxx1AcXPWem0MUgX3ZAmPcgXQxcKRswQgfc758gq6/glUk7Zz1A9a0MElH/f
tzTAMT77p4+iI9Ww4kQaD0zB3N+k0qJcrR6Gjo25LZEVrQlvEOLxYcXwzGfkGR3T8zOkiS/Ikxr4
pV81hGBkw3FQPpMGCWRFaaYA+WRIK8jocLkim4bgnYlPWTMGkXcAyN82xRSDjRylaKs6o80pJfDg
NBCybxY4GQQRRN+ZgESYbh5+QG2TWJnOlHrqg0jetbK7D/LMvbnvM/xS/WrFkiEKrCb2F0o/AahU
qnTERVikaSJ16lsFNkhHexppuUimhhQT8z7wm4sk1ipGDK4tQRBjrEdnzCUTbM7RqdCgyBTnnBvx
vTyKu86wRe9qMdFXFLCYwmB2ICkYNnV+bM+wEwk7WXduyfrS3lnc3olkuC2JJE91cqRCyB9v8607
cAgAMWYx5Y/bebQKXesh8r4p02umEZhZwoslQyiDh7/DOLwYw6AqcXQ9UKop3Sxk0Y+NB6JI9kpi
wgYBLCHtW3TXZYxobM+sx/EvMXcggPhc+PmpCWbtL9LLc1eRnE2yh+Pb4WCOxw3tBw5gU3NyKwy1
a2yROpv1IHfirUlVTGOt5Hsnolxp74C2aNNhfwuTKw02Vbwt8028+ezwdfQJsf+szUo43dlxl1xF
CAqkTJPIlieR7q/J0Dv3XtQynNopX2OZvxpDAYEzpry3O80++QZpExcJTOaIcTCnVDIlZYk3n7bF
OaX3Xjwh90XQmZByRvjosWPZwXMR0QQSnkKBSKaDeu51QfpORMUULq22dRu47q/rV/DKPe7MY7n6
u349vImtFSlWYgU/qPcjieGMbGimU71fq5k0/D2jwB7Xm7AWWUnNlrYxX+X00xcMI85MllG93i0l
P9qGTUvf1M6Nxv/EIQxl4hT91Ai36aN7tkLKfrbn+BxjTomJUne9RchFKDH1a8beRT7blkiUAmDJ
ff2sevAJGb5Aj7RnjedNsWuWv5aaqHs0W3vT8gXC6ncN5+wBlbViyjt01vTT3fXrMs/t+5NqklGL
UvKyA6DByQxsSESWh5MpDJbY6asRcVy4cwJQsUpT2bNjqRDWMkwI4FsvnYf6cqzHuWWR5ceNpmmS
88oQayAZ6G2KkE/ZgXTlDBdDXNOR1Wt5UGp2qYF1UBaZhdP2qnT7iv+r8mVqxXUs1gCvyScIcRs7
xHiTWgr0Ukpz/UiZMqwIpLiR8fYtfoCecFniIFCTyijQ41ux2WDWHhJb1GnFZFWFgPZOfV/XuzY6
rj3/Cih86lWkmHQZfp6dgD6PsKNzbFGDwCpVpjcNyWvef8vb3ziTyGcFmNUGJ3+gJWRGiqil/oHK
L1eKFPlAed2VX5n3GnREY2dVSNg6hmbOkYXb5AGI242MYxpVnJnbiL39gTpo+2Sfhp1fioFPgTP5
ZDOTQNQp3oUY+hLEGRnC87/eNabbBEbivmO+/cnJkb6FBWD8KhOuFcDhiIF1g0cDWuZOX6jPwkgo
xdFw99HvxVHpbtMUbnrhzxXd4FEiN9PjHgVCOvOeJlJw0ICf1fYsb4bKankvj9Y1t4SXNTG4HXez
TFlYvMEteU2MCfyYUY9kEnJs2gcypi+9Bdaek87tSLDcrvrGmyMI26ebarkgKqVMM7Y81X6mhVDG
rl+W9xv6q6JVyx05iJrIJDix4R9PQZ2356axigzdqF3uWr0XT/pZXTKmbJtL9+aN31NqWYCmg5z5
73D7hslHRigPJpXqRD4VA4Z/2AWx6rkpTHTk3lmI6pne2FmBx4WPZQOe4Pdyxuf0l+2uc6GOo86j
KGPn/wEV0bDStYD/SeqNZn7UwRAW1QA9WsiPWzBUjDNZ6raXt+ft6+s9NIXe2i4OPKXfndXmBdpm
NO/gCZdmalcaiwaIVddy0r/nXy3mZKMMoBDBseFFMorFjocyErbTITOTLoC12qRqxVqQEPZUPole
/gu9A4OygJUeSN1MB6sM3jDoQ1VgdbddWfqeYXzwcgIKaoUqlhgAyHkaxxRSODW8AFt0f+5N//cn
RqXR+XG2lP66M0wMyyIY453GKB8g1/C+HUzwnCu5FDUEOcfxcEO6BBc6eDyOxCRqhKiYd6OSTTmf
fKqJ43R5FEZaOQFKsTr8IWBd15WmGsdZndYXV8dYCXxIrc4A4LEWgD9FHGANtrFtNOQkucOO2HFI
/E2/Q8iEXvwQ0EJjSoynSFs6/YUm2ZRX2kKd/THruq3TlzGbKvalrBA0nHLF/x5Y0XCf0JeC5wY6
JNHk7s0nKNtc9+LU7wBerkKyMqZ27CQmrjq4JDFUT+F+vKO3fNLmMUeOQBTbp0nf1L0lIKXTj1HL
s843P+LP5uQqC9n2kWsQd1T4eZLD7VVId5YbzTQ2YEhWfE2LBn6yFVyktRIkVp/RPPFrfPX+1PuH
m6bXwWfGqb4tNFIA6x0hdihDyRMOQEHuqo34anVSBDrDI/flozI3Gi5++D8B4orM+7zDgkP5P/0L
yDv8mrKMirc7u9drXdolsmyRkX5GXjVhM79un+g4sYGD7ZmZ+gVpEHDuhUZdbdgXdtwispr/sgNi
O7DD77RZA746Cf9tj5+3bCrFN/BOcE1queCAHG0YsLBxCl/3+EadGiiZl6h1CI+pUAFaGdOuXo4e
YEKTdjxJPnUtX06ILChiVmnEwuZ5E2pDXmh7P1faw30MhsnUxw+qjQSppm8yDdX4XZoUo+6+ySAv
MLNOLgEYmtt1ZOJ6UbnMYW2tSdy38/kjsGP/HJr504PjC4ZzekZ8zQ0fQlwE9d6MPZub86DT5N5v
SgtNE52737Yvb45ryAl0BaRQmxPyfEZTJrF4PF0nq6O3nYfJUhk1ZKcP7VU5/O+X54mJ1PQxWpMY
2euNubCEO+VgPCT3ISn9y+RZN4NCzlVn0K4xkYUobDTC9Hc7RhC44U5gnwkr/nav8tUP6DfWuMse
9bLcU7ZoJlQsXLaJe7CSZCfy5fcnVUPINUWfSJdefvs2l+vPOsRVQfCWneBOtNkv8UQQRejseo6E
3Se+NWV4ZIGDHv5d0UMZzkYzdKgLnUvdMkIUZLTRaczo3KF3D6j1SPz9JJE9LO+yVc4xiGskhJpW
KnvFodAQH7rWOh8uC6JKsBL72SkDyC2wzrxa0S/sHJAyEiM8hGh+t0tpnGrclSiVxtZsMn+6afB1
WKVY34CsEJx+IwWdFMQLQhnhj+JD3TOxmeEjB8i+n2lJ8E5PF22LonxFAkPoaq87elS429tell2t
/nxe6nB+X77AK3jtonm+LIhdWl/moR1Ib5kZBtj4up/c6zv2KadZAn9CUKk0gb/bgYFLm85kb0sI
Two4fpTKm/n1FpYGp6oJcymEFHJTQiMHJrfDWtwLLSRXpqStAkAoFeZuvZfcDfq83lrUtDg1+Wvc
Y+vHb8i7CMHIOxfwOqtfuFJTWuqqFmMvx0m7CdyTZAnemRyH8vDuauuE4cEUYLguroqacUB6qPGc
AkySuNltw1ASUICiouBmEIzR4gGDihJKhwoBYoCLLkChwEAURlrt45rx3HvX1pCBTQTNCMtG6yDi
Ga4FUY4PCAIY/hlIDuDNQBAKnZ+Z0JjIdmBRSeCjEOLaVHno0k/i8hlqqakIP37/ueFY9taLsT9z
1I7vdr/fvNeiLA9S5GmMGcneAkR0fiNX8sL8JcEL/UvOA+DlFAGvm0ZAdChUQTj40pqwA377KdtG
Q4RYsDzGk/6dCWknX7F/ukizPLUQqhPQHVr3JPd9L0/00cHnM6afegbwxyGgNuSqBFs1MNRldz91
poYlvxdVyBtJ3Rzc+K1XNFYiuoyUw99pBb2nQRZ7B+1CeoFgpWi3uk52xZAlDcm1B3NfoAT10t46
qGb+neamuh9cPhF/PaTeb/o7FJnsu51mvlGP839B7PHGA0ewJ9R3Oy9c1WYR1YyNT/nBoVxfS1GK
OID/SqQeTD6c5ZMUMUQhQLy3Sx8XLvVm5RFfFilVfp8WKRy+B/C5RE5bMomy5zgyqRcUP/EFHaQy
nA1FdeLjQ1VkDFC8DBaEHJ9XeeTpl78OOiYflUVh6uZLBOauOKkJS4t+91N6E/HIxh70JPJsHbZy
II+fW5+NAgld9r7A9efrmVWR0R3IMLKkZjVSVcHWIrbuJrpACMqm2+zxI5Bp4b2/FIEzPj0qVX9s
iI3uW/s00au9zsGkyl5vT2bZ4L8053aL6MU/c3enIYIoYXgIXVoU/ljMqfJMVDTtIVASvhMHGCvs
yYQVHjia8fsEywUwnKX4zDS5uti2Ph0P1XnfiNHmrp8TZaAQv+uGspGVTiRDXSg2X6hnGTM3GuHD
wp4ALhhO6AX3WVzl41Nfa6y2x0uEmh6WDJ3ehFAElGoa0132ogvfGfKmROiM2zhticep6Btr8mSL
RiJUYtI/M1tswWdJRJwOHkkxH5GHpfbWQeWM4TtFmNuKiD28xqJDZZ4A98hfMii95+7p5iUy7yyi
B2PcU7aPG4L1PdBousNw8CSpjeLAfA2BlJ42wNzddRPUN35FEBvyDRQErqgyIyXi83J74sfoBhji
llE64JZd+FIdsNP7ALufmhmIBov81JhNQhIB02eFNmh9ggpr7TNy4+XWVtzZ1Q41dPuaZni4yloF
Yy4bxuAOyEXuq4HpQVyRxdmDsUCTf8YBzuCh75Mv4R7yuEzSCIGIsx2C31dQMi3tUArEod4snHNw
j8bn1oR33YTFInOsPDPD1NAPj5/fXrcq+bhBTQD0d2SDosUfDGYEG+KgTuSghs4LHvxFq47z78dt
VkTFSCtWJZP581Giqj2N6c3ySGLedJf3egDzy/SW+gVCQomYD9HxOQWGQlpJ5C4GUYCemib606VN
WMHr9m2ZuJaFWihEasmDB756VrgAu/+ic7hAOv0JeTUnsEVYJgb2nlijLUYKQ9btrYtqQc2DSJZI
kEVt2xpqgjtbOZf0haw10NaFCD/pGlQmNtAD0Kc7AVXh/PziaHQbfMM6GfCPBbOzp92iGBRlW3VY
8bC+Qxh0Itug6u6GqhP/fa2nA3y7kfGmJBpQtfb0hOEGdCkLG07NLZSyDp1Hi+rRdD1LZd6d/Uzr
yiIXWr67tgn9SJT3ipbiFECp9wQafNlyE7V0nfCLakh3lXEWN3wLhWyjOR6TsSEYoRU59JXo+ERv
ckN72PrOXKkVQWPXL7ikcN0+We99X+iYdWmJ7xjmrJIT4++vZVGxq6GAkckQiD9jdqaU2lRP1wpk
oRiXeBZu/UR6IicgfCtvDm5dLB+0Cmc85cZE6C5HvqN0kJL/ZuG2wFP+yYeT0VcG5Wabbl6tz0HB
ZDsrp+KqkNggeRU6C3vGaT2R+U27mNY5ZNpM9fezVabXMqyEAnGfMRJLY3UWWhBP3GeZ/8tr47Da
uwMg6m8lCwEzQUIwoH/cERjXy+1wzks6g1vROnyABD7JHeqML/TAaKV9osEWYgf81dq+nED2dFbJ
3pfs9yzf3VCNUSQJgsbCe9aDUp+PHsBqhNSoG68xwfDTT7qQFp/rB/pjnWhsSB/EG/oDQzFwwJDn
54uwo0+nvTcvLHZzIcrLIt+NypraGwel8z4GuVl7WBMr4F4/xHWy6XrJrpJpypOUGCTxTu3yJH68
a8tIFSdUQhWE1XR0p4jqXL2AXqDwNGa37Z6/9Tld8mU1ZehCqV7M+DbWJ5/XLTSLgTrSw/aH6Vr0
j3v4mfrgtzve8nq3yRQeei+6BDq7UrvCWjI6DZVGVncyqvPaFpr8WeRVwI81sCScOgJgADW9kj/f
v59L5p+S31RLZis+d5d85sGg+naA5JI703pNy7ixeA3ModWWfUHXG7xh9m8wKm+nfY1cL+ahiyLg
iXV4dGSnV8KcERvYxGguyEDfMk7V+ynAszUKHhFWhMnFKSEJgnF+oc7hsK13pEGgv5l+cvO08CvE
Oo5dRrAkv1aVzkc2fcSDOpzrtzw/9BJde8kpMJbGbZYA5XT08cwfVpls4Qo/b9rZZ20iD9aFtZS1
OT8hkdvvy4l5553YHLeFpXCJNHZhiLP9bke7kCX4pIU9+tTjkd2lK99HUVDpIbpka32TYceGIsn/
zZIfPjdDa+i7m+fqXvW3VpnTGqdcMS9pjEL7v1UzAI/v6tWj1d56fvQkwrhXmN1qtgJyZmwPqBG0
zaCbPlGjxm46qIfCFig2b0csAW3QSx6c9yMhknY2mYBsukJuldJrge9MWyB/ElavYhOb1+IQJKvt
Ae2kKXibwXRQAfQa13czSl9W/ztjNGR8OfRBWRP+7e0TeiFTNTZAbhkbH687LV9k7VAGkLtgzLZP
J5fYqPf9ySqD8Cu3rJlQ5ihMEKfMi00WuBypqn/+5BPz0b6XV9junfQzoHr8g8VxAfyXZrQElDrL
jVqtE7cfXeSI0uGDQbC2gmW72yXHDgAbu/nVxySDTGOb+++Hk8e3gejlUaTcrUDYS+enNuBNN3kQ
bSLR7XtT8G33vxxPAD88GI7MNcxgHOcQ5tol/1IVF88zZgfYej6Y7T2HH/JDVUkQy9HmX0PgUWLH
fOxgtivTzUp56dH+MzOcITcNz/a5Q5/ugHfW6492NUYo4/+dg3uiluQwg/1jiBF6g9InU3VqttfS
+hevkClcVWvlT8peJbZzfDECp0FBCsAufmWJ+NRU0bvO3d/urOxlPLwtV8Y7YBLyjikAO9X0gdB7
O8N7KRlKTLhmTeELq1tzOw6m8E0S8fbMl4QIok+pMx/mrEar4srsQb9cXpK+Ml1Iq2p3mYrqqESY
lN1g5YFa5fmhX5nNGftIOgu8GCstJn5YvTeiNSAMkW3daDCtVabKkyITDzzfHeCeS8xMvyncn2Qz
zgi4gWQ1vyBVONZpb0ZnEuWfrYvdzaFL4PHgK85Q7e5bsoATk8pV5cs1BOBV0pXAZtYvslU8AhC0
ot/1ZAbw+kY+y4Y9f/W+oqR9dL71/zHk7OT6t9DM2Wdoy5fM5eVb5SwvqJyG4/QiqZkNnzar1zve
rX9II0gxdn3oQjcpyVLlepVLwFmQWkd8DD/SbHkF2QJjytpcg1lsTxr9StGjeviWZaMEBp1CE3ml
G5AIzJ1E80UqgpN34aEt5uu7mXXe5E+5SLiY3rUoCO6PfQKmBTJSYDxvc2Td7YAWeVzcV5EURFP+
+vfCIsGQM/83HmzxXaQMEuwQB/B6EUF23NfWlQd04o8HEeg/vC3nJFbMYpohJNlGSS71L9dzMCKI
3JnOzYcJLim91OP+5VCSWFczyXS8ymJtaTk2t/yQC9V1O8rWaYTfFOwWkR1lMwWKxmjwR0pr3ECq
wKPjM3Uu15/AC0/3gK/FFb7xIkpLtypBLfCj6qiHv2/6XCmFOjDyESqZUcYNLhrLPvHIOw5QenNM
GM8qRe9Mo+T4qLFvH6lu8BGAOrDC3uZXhNSPijNQTQvX36uRjL+Ni20K1hxnT/62Mhy6YHoAlbc/
CkLF7kKKHNX6AXbOi5PQyoXHe82ViyMYoL+OkpFSxLGts/vc/DXRrnC6scuZhju+1+CqxgpFilsm
mBUjCp3mh+n2epHE4YkRs23wrYDYga6fu0KNgXwl+HikaOZ5gPRcoIT/AGFft3I6P2aUH2t43M1f
GYL9Q48aeFwXXL1GsAlI4noshmEyUz4ACfJSgMw4s4ZYsqZiwbwyKMHcQ6iY2dEedYgB75g16zOb
ogzGGCIXibey4mZkohmFAQJLkW2m+S6lqEuXv7vPJXHStQ87yCkDJXqjjbsC80b5JYk4UVWY18MB
6O1XDE7EyIVOsnZbZHVQgVGyoEi4jAB7CNN+WrMhzknIac+ng7FrJgJFeaSyJOdb5H2kAcUMe3Ff
lzaEHFOv73W1nd7C6W3cnY7XDZ9kbxfvDXtEb2EDPw1NWr4Bj90EL5az5ZQE2j3KzfRcwtKjhQQI
1SinpY90uRii4tyFTh5Ij38IFW2wTrxbjGnmR+aqMobl8EgxAklDa08w5mEH9k9IUGDGIPKU5Kpi
DMTXnj/FmmdhQ6b4aOdG40eTGTXYC8f4NyDr+sNGhsEfItt1GUVJ0g/zalvU8WwaX8wxTU0Wmk3b
qI4nLBhYyyctWMfMzVwqkOC6G14JqyIcXFPcqZec9kvVhpgUfLj0h1073cDlIIiCcSfvNlpqyeLP
PHC7NGVZZD/KrVLtV2UmrGPF0zlHBYRn+njZRkROGb6V6MWLYjZRLgQiI6Ss8iUd9v2rZ/MijdyR
iOjUrNqWRj1BpOpida63xtN7ZDKNAfJeU+utd3p6nEt0o3cY9ANh/t7wi3Z42IeihzXjaaudQfCf
ozbAmxZ6oIivNpERJc4gM/C3gzNkigGAB4gxxvYtRCzlEMedfA8qr8/0f874izXDbIbi4EmBwWK7
0XAqf3LYPiG7pOOR0p6+YNAmBQFrJraB65yg+ioe4yuPW+sdhtQVsI84HYKhc0dEI1qLKf9VzkaV
YGZSGJPqfZHbuBQrUJwAPyK/ckJcMBajYo2X6oCIsdfMMdT4Gh2f/mRx+8jWLkESKmaTSWuh1jjf
lcBOO19FlvU+w+KEsMeYu8n2K5vmE/fAWFhcAMDaqM5NwpfUCYRhk2EcNRpCP1bzRAeQo2X+oeSM
lghE8j9DQJPaGLAmk1dOAdNdoQZpygBmZhk9AY9ngWMX0ntOA59ifNV4xE5XZVgsG7Mn5oHYg4hW
+sW9oE/Q8k3DyxTngfrKjTS0DNgdRznfxR/l38XQCoRAPrQDMCO6vroiNWSIttnEGiprwuDPRU0A
M1ueSmzBvv7GTghIxc+zGdp8sKAtetSoOEa0UtWtFEeGYMMZ/v6WqNttZD0Lp8Ijw6et76VJ1WAU
/9963vZL96X9/W/V4tNxgW+GURHNOpRhIYLgyFYeyeYh5sC+7BUz50hqmk9FZ62Mcnx61UrkaB2J
KbaM5NjO/rqTRkCN/Yo+VqmlIE87TjYQTilp64TVBq44Mi7Znuo0Kf5+eBnD1rvRHD192TaiJJ9e
2ACpQ6nAWVMbp98X+VVxzqQnwr5yqqbaD9bTZTCcekGVwYN7RToiVDLPzr65YPg/xohFsqbiVXkS
33UJwkQvoHXNXn+7tuyaKZ1WyGw+bhUq0QtGpQKNUVybdj4HGlSjlJzak9sQaszm27t74vOnnVo1
JIWG5MUoFhz+l90MPrN9iQExxJDCti4HWBswXmuAXIM/NgX4q5IYVEg0CCl1bFtnZRxF0u/J/1Kn
wuNHqaxzCO79C315jG3R50nQXyXYE4mxzY2HYR4Im4rAP0wLITDGid2J7CMPp7kTJjrueiTTICSH
XyK9bIKkTAzp5EqeOx/UqmFpQ0zxKzV9O77cTYjyrNBFMYVvpbuJX99SM2cNxcNT+DAJ57Ap5/7s
Z4zsWgoQTzCheKKN2NacCZQGZ7kc3/JJ9CLU5lEWnPLFLeVzQaYagf97zBvhg0r7EhyfXx+hv3Mp
tbeF3WCG7lBeVp5LkXFLV9Y9qjrPhck++505MBKdB4EUDJ2uRiyaa2seCRqtMGXi7fbAUw9YgHMx
U3qOOge0q5ZCAuJWuowv5IaS00VcqYA2VnZ82zGnSaNxQFE9ODC0PuCAdGHxWE6s/Y814qq3+xPk
EgJguRdoHNl1Y9SywyAg2uGp+PdHRbI6r768xmvddknx7SNYc6CsBI4c5AMXso4H4L0E0M4hoYFK
EvAd7LqP1Q4O1+9fvcz2LI8DkZcLcUGz+JaD/KtfHl63Ql+AjMuffPKDZMbgNAzohE81JUHSO1yV
5nof5EyA+JfCe5O23n8/nz09/Mycx6ulve64Nt7WAISw7KT5Yr2Rn3S8HtB/IW5c98nBORdw6I3n
WMkkg3xGHMRiIlp9y2i6CsadKTNRbxiTfq8VenYyCVo3TfLvWOtdHqfyS2Hb6EPmJ9YL7t7pfY5u
mLeZyv3Ah28sYdv9fMNdC5vx22bgTWIv/+HizpiYS+/JL9+51684ViTQQuzVHnD9PKjieN2HHuVk
oii7aLMpD0LFKVcRjY/YMIgjro6163JE0oWIAOT9S5iB47ChU1CIU9EwgHTgol/hOvyl+UUuqXHT
ZNmPFY33KprjnBbOsXiCMwfakapQ9jgdMyr8STeJMtb0oW3jvGqZzJ/s6B8GjOeET6qL/2rg57KT
aG6FqrcgtSgDDbiYcmK8jttckby3I30RcldMKj6SY+HzW1S7ejXpzxqWnSO84lYLM3kSqp3TIras
NT6bN789r6F2LBRtpcEBksVVw0VlOdfbnE93sADMH49+1bBgY1FRcBRZZ/3A0H+8sn8BSNJnzT+H
4Juge33KmowSW86rPlHhpUS8Mt44pmEmt1XQYXcevU4egtPBXoATsqidCXVDoEbAFUgt8NOs1P4/
w7cmblB8nRarAD+djOkzFM/xI86ByV3ylQhArVmpOfAkPKtYjwDwAfXn1REqIdif7XvltA5rtCSX
3jH4vUTdSDb/MzFzWF+GTRZ0p/4zTEkP032MII0Qe6aQfpyFNl3IGvnaR3U5eCgM+I4MpL6Fb9nk
Zik/1HZaabdTHkeRm+6i/iQwWV+0fyxRXHyRwYYU7BQreyvOob1XHF9lPT0dGCmKdMWDRZpoPh2K
hKDkIhpKZuRWkQ67KyTmWpO+c0tEXQ9+IP4krJEmN//r6GZcDYkXoHp2J9Cc5MMw6wf7eUHBcy7m
wSEI7oQxrkDBqgTWNAVXhE1TJ0+cqW9sYOXPwip1MQWsmElBSXB7E7ElxzuDUy/Ao8d7QZQCW+8T
26VXDp49F4doZ5WN6jFbYX0f1RY487d40/RoSiYs+JVnvOqbumKLtTHAgob+eT+bjZ4Gn6bokcQz
Wi33q8DXdgdQdWRhYhXwGbyXDz4Fm8Yr0xsulgS9K5dZWWgBJo9mhbjTNX/uFPKkEuc5r1TKLEMh
Le/uFd26ZR33nrQBTOYkZX/RDt0KicBtpdG+syP7sFJdyr0FdvGf5LUlxI7Ccvkdb49INTBk7qNT
+Nuv/tQlQsEqfL+5vyvsIv5U33GQCKxt6eFSU7Sb+DMBQKdhvZkgqAtSr/n/CdC3d94nGtQAiJdO
Q2a5VpGIY4Umq2/kxspMsfiKJapmP2zhTEUlFSPz5BrlA00UAuWvZ+JZZ1XlOVmPAmopoqKxPztt
FgUAmTXXIBv6nW6ucrIneWE8IyOS07w/uqst7j62b1BkRAIkFdEctmzMI8psgnGlA1gx9qqtbzOE
2P2CWhi+U+hpSez/Jik44mSlrjj0yG2bXw6IdOdn+RaQ/u4hUjdGQ64s2PrUOe0DLISsLs8YhDIh
uZE84ipCRObnCrgCu4TUgIyalklgSuJ28EQ2PIqMpUdubi+OFCLA4DvQniMvPe/WKQRheGOiQtyT
mGI+DGMnPpv2A6Wp+u5dxPOcbiPnib7zc5mkKt7JOucbmgLEx8Ks7MIjjQw+b5ykFdqjl0JKtJtB
l4VRWtDEU+/ja2mpzOzpJYchi9++9OLFm4lv/fjJD0rzTXr2+5AkDB/dVH8t5r3OMvU9bfpCs9TU
AiSu8J58zsRnTK7irZIjx9eirg/oY7asuvEf4Xll9SgmS6s9TLHCBDAvDSpZw5yL8ErBSft7q8qq
a0W8gfuxpuHXcbWAmgiGF+KqhpZZgSoteI4gIz0nCd7B3CGML7yI6hcxVWdI0hD6lykfyMLT8cUo
q3KEAA==
`protect end_protected

