    parameter   NumValidBlock = 8192,
                Recursion = 4   
