    parameter   NumValidBlock = 16384,
                Recursion = 4   
