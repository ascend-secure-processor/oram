

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qzm8npojBy5X6iP7jyevIJP3CQn+/y5ibELWBAPHJDDWM+rA571xoKuK8oM/80ooBxMbkVzM1bM7
Do0ukVUmoQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d1em3+E4PJs5ThHs4+oMmnJxLj3tD5+Ra/5RsbjWP/I4Q7yCQkHNK50b8ad5w6/29ukBqogecpb1
C/z00aZKahRNc1nGB6amPP/+zQH2BikQn0wIa9ajIzTq8fofwJOer4JISGU96P7ksvAxy7uVrQdf
UgHjeDR54WtHfXmCcmo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VeWCfNtT1SfugmTw9QuiIMpE/0/Ol0qTe9d1O75IjHhhcPsTobfUrB7T7Y773kY9iDle3arydGPJ
s2ynUVb6OPvlbQlxcl/OB0ax/USEoVY7kQM7/E86kxioyoq5/eyFJxWImSW8X4KXWa5kVBCX1Fe0
SM4S6xnc+JF6QTSmVsIsCI60YwIujmumqwvRSSYb2nCdkbilvK1EW0JRRhBM1EFc+LOhgJ6RM5qE
zl+1hVWMtY+G6WCMj2j6wRKkPgZwZqF3r4hK1qrBIsP18ic/yryunLNLNIfx3LrCXpWH1S60LpSI
GowjMnkJyTNrbzPOPchZUxfEc8UJVfoQD1iJgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KeiCZKgVR7Gyj3FuM1ZQpqudc531MqeOtYGyMzjuYc1CCFBWg4ar8o7sj24KUAdwFxGCjtA8kZeu
AC/QleKkLVBkvy/nYQ6h+tCtkYhw4dFqO7jQH+zmN64hdbxtLKMMvWGNcBk4RNNDw3tCOy/fvcSg
VpR4dfNmwqhOxECAL+I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MBqlz4UTPdTtYsudqWtZ2XIC87j7URCcdqGp8uSc8nsS+26esIXxxekhuvPNueflHk2SPMoZSSPj
kPwzacuJ5NrIgyKnvvuOXmf99uupWSGpW2uEnGxbNEh6mnnkQlEf+84Rr9yTclKiwo3DsGY8uNcB
55Ek5dQOyZjFRdkaUPI1mFy7jxoScAOFocTGRSDc9zrkQk1/KyW0yChIJygbi6ZJ7IbTEcDbxox5
TXK+7NyNj5qTou2wY+Qnm0NvhC2SIC48v1rlOFlPNy4/afwGzguKo7KQfcSBfV8S/P+ecGTmu4Ze
c+Qcb9SWdwb+VBsde+7H2KvtGT/Zu+NTN+/VJQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10272)
`protect data_block
kQmiTzRsQYGyN7ZQYbRaAYldO7T80IMrQYr4bo/rZGPyR/1vNP/AFJ9s3umPXnqkZSCnuGDCzSbr
qrU+TM7PeoCm4poXyZhLImOIgHgZaPdMkTXgqQ8wJJ/FPIM2pYgv+AuRuFj+8kri2UloZCUuwxeb
/Cn3NnMMvhUCMUB2tAQqP+vRAoLajfKe33lZTixLgdLD1vn9X3/ppSbZPrAS3zp1mLI7aYY0d/JJ
LNOy82f94zq5kmPB5cb6FhXNmRAMy0a0IUAohbrY+TPWtkmZo5XapEpuqKpdbUfjwF+l2XDaV5kF
sNr2FR5FzLGo137Kfwhrlv4IDQ7c6BFgQpHyBfGi7/S4ftKdQXIHKc20eKUxMxFt/xfDC2JY1BKh
xUS4ECXO5OdqZl3Kfx+VR5IGEFfsHTgioUdbuMPwzvrU8VvtPikEmEHC8Rcu1jv/0/jj02nmKHAG
nIfVZuCdEbLUzbfVKpJHHax4zOknsoz1hPf0NiOmCf/pk4NycD6B24jv1moppGIg8XlkErmUnlS8
sss3usiRPLKNBa8TUMGHoZSeRYGWc61yJFKeRw8gfVN1IaI5RJZrgGN/ZN20lQ6BCJnKExnUMv7w
+FsKC+6JiJj9pMlrlSrMKiXW2maTKlJA2wPGHmAdjyBr7SVuAkxhSxX7deNYF5WQkxxQS/cPsB33
OrVX7LutGRE3sSLnwWXHIcyy45/pc3u6LHgWds7ksAp6xsuDV+V4uRfB0YWzyMdahiCvzwjvyFcu
ywHfdtL09/r/Eg36ATDXV3exs4epIF2R440M7UYQP3Hot9xpmWEzO468w6qsRzHpDdDOJWZFPvTu
GZV9192Wafo+yQdVrg7gL8rKx+sDtm5rLjrawkgyo59BZIu7jkxX8OVFTQVuqJWyXAf76noUgFAm
Ew46rNntrGh2FGxoE148mCgTa3TkM1AKpjEqhzfNypjXLd0T8Kc4k0Qp+KrtZMM9K8T/YWmgWUQt
9D8vuDL81DlcxwLw29lt0r4TkuzjVUZ2f/OhgwSpKCe+7cqnSfxaWVrOpa0laFFCHZrwoqKA71bB
VUk2kB2Sn4RjLSzobpuR6vKLiIklnXTCVFEUlqn3qFaXclO8CyF3TA0nxeHfPS4stPxvYDr3tctU
QHNXbitFqV5moj9eTWl6GRbnN/O23JVRXnOXZ9kV0Z99X6RU0BFFmz8e9UCA7/AIsuvFBEo4WYX7
CyTqpeiJhnJxSLsJB8YxG/Aahsf0p5GFt4xxvQh5UI2SfG3qTdAe5bFgTPngGtaLIm//4HvKVesr
qr0eYNu1ekchVLALmaHU5Dcin36ue9ocjBlqTBOW971azuGOy/KuKnnRJJ3WaWoQ5cQ/x/D39S5H
Q74KZORbTTx8gSq7h65NSH0VQnQtAJLskOkFHHm4fF0RMZQl7f82ClUCggWWs/hgKjgSgwt7X0OP
xyoxG2JC7MfAVVhzeTt222ntBThXMzD7RnTa+xTgpTBUe+MSGw1PyyItezMjSLTYEFUJTqUdUVUD
/sg4ES0009yzQrWNXeAtVb5mqDcKQJd5DHMJ2/tjpdQbgoVdMtz5kszrhc+8EsFok7DYGp7HgqoC
FAQHt7Js10ZiR8XutnxAMc1GTkCo9u2LtolOdKZ3mNldvUseuEHy11dstcFH6q0oApt6+LCwqXaq
EXj1cccqoGKz+lpRKOvKcnFuVle4Fu961s2HXwUy8yeKPgGSfaIpf5VfJ9zSWfjipSH3OK2x6wNx
FgkaWpiy1EV4vUKc3Z/wpB/jzdVK9M2FDWNe8FYqpzwSD0Z/ZIqPJXbEzd1uk289/oINFRTdInwO
Zxizu4brNsatxtk5WXBMaMEBipp/eIH9RMsbXS5cIPSyr8L7Lo/vRNWN1PNND20o6K4d0VRFCcA4
Vb51MdKPVscmnkZkk1SsXKXGKFh3gFtqPHz2ADKjfGyrkAL86B+/6b7J2BviWBVpF1nnjpM0pNHl
YWKaUnqSOrVVfThy3HQ3Zf2xvg9FQ/EpxBslaLVCsFYot0IhOQyXXe8oGxsEOf7YaYBkpdtrM9S0
RfJPEkgOjDZKsUmw5BirZLxmwV0cS6LMuojO3UWYS7BDwS7KTU/+pptJgwo+nEIjT3SJLtKt+JbK
5tg9hqoQcdc5XJnrqmrE1UrJfN0TaLi3dfGJOzQI7dHg7X+XdVnFmzn5jKtVMCQ2DTppwU1aLNeh
eH8uPssRfv4m1hmRtfGi0XkfRsFDqnGoth3dtOBRDZqT/SG2vN1i8U/ckZWQSa7sPxnurpzU5r8r
BFqkDLIChAzN5s8zilVG7XVbV3xmUDVmP9TRyMtzCEvuVrOLof5yHt8565jT8K66igEsGaD5RRn2
76eZSoW2U4MrTSMdMMdWyhQMe1qieE5L0TZw/UFw3BbWqvIcu9FU4CKWNFv1wK/wt3l6x0aQALas
YblPRzruK8e6+HMg26lJLJjigULdPZPaxCSNN5dn0dnt+ae5034Oo3b/LnbxsmScbO06j5T1/DBM
BZwtoPjrbhrn0lrOJ6gfrd7LvLNdzZaUY3PwpDUd9tWuuXpxdqNsorOTSNL6gDLBMrN2kF/fsrFU
UsaaiWoRNKTgqpYrXZyZp2W8Afi0b1ivtyIaJR103/QtCoinusjoc89shQiKM3Iw8ky9wU0u13XO
gxWSgnnSGZF9O9vfFIJm93voudWLlr23JhTMG5TP2Uj01SGtAOrsECHgcTVI4ic0wu4E1+rS/vKX
OZ7usVpZW03fMVWKd0qFybI5MAcXvgJ6Ts/a3cMXALk4LDp1X3+wfgQGNBdG8n/s4ozCqPueSa4s
YxJUI3yM/ojacNPy8XDREeFq1fdvo0BK0KoiM4DnfwSYjzJ4IFIdtF9+visrCisThe2Ou682BG/J
PjkjGjKI+uBjL2gWMjE/tvaV/tBfU8u4EVDcDAlmwQT67lk9kUJ3tibDnlm4F9K8pURwKPe4jbEK
TZK7ryjIc8zYoIeNCxwIEXokz2Ywo47ii53yPbl/ipGVkJgP/iJwgQqirvlwUpQkGe1yJWsnzO0o
U5QKmy0HrUmOo4Emepzxk9XslbW7GlIYNKQEZZ86IK+kyUw5gUBXAh0gkoIRj+83Yg3A6RILqaSo
KQ7J3REOQegbbOH4ac4wUYe0h2thHegTt/yxKMOtsGhWumUBs0Qu9kZBe68g25NranDAAXerQs/f
SkV37OIaOn2BeoX0mlPFwps9X1D5ZvSzv9RLXdvvnlyhryFQvWvEDV2EFxZYMbOj2X6Kj7m6eRKH
9rNPvCMXBjgA63KB6BEMt50oYVdDbvPPA4fxb1jNOARWO2wHV79QLSR1U5yiS00xMt9rakqCQFXv
ThPDZjgzf7gul2T/eG8rzuuPOAWM9twHU7v/GRdRwHcCOirduDED5+fGzDWbMOak+ON8nzTIeJDW
vcKRNKyCokeCe0H1BiU0qMiuiCMGGhRDBvpd03OIPfb0TvS1uH94cVHq9jCauvrArjYidaIRFGZ+
Xe64ueZsY+sF+PfIBWDyWlZHFDRz+3rcQ8+QkJs8abyKE8WRXJh0B1YFESOHLM7qIKXZVn7pYl4R
aOYzo8y0nA+mkxIWuBWAp7ewGoZMVSxOpQPqRmq75qSrVigrJTeyY3bz2nzn2hE2EXSO0ARQp3Ca
UXIkfnWfWT/xBv6LQ1h69gYf4KyYR+ATWx9vGIgkQWeiT4nh9xNxu24NDc+YVa7RsaLGOGxSjyAI
UaVH4v+N1xDTl60yBLgIA6PzDer4twpTPgEm4X8vLz4LJK+JiSMJ/7fu8Z1q1EvKZxb+CgWWwSM7
lCPH2cFj1Ggga9lKGDMi6jQ2g0USiNpLgt7hIekSnsiwoYa/s4Cdqk+zYlYW85jwKwAtH1lZe7Mg
HsM+gLdBT9wqD0sOYQhAlRvBC7R/vIq9kO0Ufj05fZp5VT7G24WFj5MnIQKJ6S0oQoYOACaLKAtY
C/RO9HoQSgVvqqrZIW1BQRdF25VRwKyxgzISsTj2aCUcEyRooce+ydJyUinfG0+rJFJtF7KcHndY
w5qOrqxHlHiIWfUHIlFaoJWDP2sGalculA+lfcmBXCbUX391TVE65LUOcY5IlriYE7dkw2kaHAQk
BhH/8+TWibvdZ2c0Qt5k5EbGLbcjw8dgYVVyetQbn8h4yhHdG2iwdTQzJZjmAq1sZwmyHvYu9VHX
wTUWHjWzsCCfxNIlTmY7nFiIRALhDyWdTiagWM01WT7DGhoC+4Dek6XOkHt7p+O0QbzIuzzPIaNv
ie9ePoTlg93bp1XtVTrh7+RsgkxNrepT9VDFQ1HR0rsTs6VlBNG5ylRtIkumxOAIVuNU4zSxKqFT
ZCVXOSOg2TcPAwqWnsd2YuZVgrunrLTVoHcehM/w3YEIf59DoiDyIx2v/3lU5Ei44ju5S/q+oULf
Wsgm9j6WSMeIeoph3akjFdqYpNlfrfDseotFLy//wrg5CImKqFFzIsdhXTkjjGxFH3le2dRmLR++
PzEPBkcthvQvY0veaWgEvfkQS7JpXdfyrFJ7oyhx9WQ48rxuA3oJVnSzddcbTCAIoSnT8QRN2YOZ
/+CvzkGLTss+1Z90J5V8WxaQmMEJp24uyCgaQSgbaUMTAuUkGzIiVzhmvVvowv1RNNp4zu+8Q+o9
dRJb9iVnIpOMbXVXFjgLMyvLCc/XrEL1yEaQ52/aZB4rMmisW9Kq0td+S5CGuqZflNI7Tj04f1Qb
Le5QexMtGLs+iYw0sjEm6/hLC8i8Z0BXq2VdWe3gdeVDB1xYu0LuVNnaYHSKkzo7DDkFu8jEsbId
j8upvhapXrIdYWDYcw6dWS9XiSNp9cO7sCOrQBuCuYG0cM/LdxZvKQhKc+rwSNlCT/pBcJ8YViKO
UV07U0tpO6Mpc2PWlkVHkobs/4SK+wrzQxmfkLq8i7Mwnq+XksbxiwtvlHDbOhL1m/ThqkGQVB/t
Uc0H3froqo6QxBBCMtG/etR8IlUvaR58rwEIY2YB7/akOQ+lxXJf9eIbtLlxOYHMya6W6NhHHQVM
pqNVSuMSkT8Ihg2gNbE5p9v5GG3dh9l7Hez7xbahnwkq+hdLzvvR0M/JxER78UNOrHV1wB941mGX
po2apuwEFxywClGh1QUPOL2gEqGwsyv8JILq0p6f1VNYJ9/s03OFifi7gnz2NqxSrBr7hXNREixf
ZmdvssdRKY841a7qQ2BzES+YgCPCP8RvRykwXaCCsMEVOL0uJ30mT4mmjbe5qaU/etW3k2ZtpQ2D
Z4KxDS0EOSR2c+SdZ86TNcflbLle3mmFvgeTKEfHC/Vy7UCD6h8DoWApjUYYMPWeOJ8mX1Ig/7EO
4r9WEjO9FdxbabCoPfuJu7ZYtj6VfzdIv2yszc7LIJaLPoNs4hhWIZtCi4TctWhS1s/SSq9BSTlb
Fd4DE/3T8sdU4DhdCSoFQ1Md8YZh4RmyZJLvsczsygkv+Q/WwsiiQKXDGex6a2JYVcu0qqpr7qT3
D8CRIvUdfJGXriRZAS3ymzbXdDUKU86FCirbcnXL8QeFwDqrR2/FygdY7m9Lq0+WRyd6Y/ai0smh
hEn9NL69Oh7/twvfbZOE2d5GPvrnjbqYtMoaADq2+937yPClOU5fF596h8WOKFyLgcPuEE9LjRN+
cwBIgq2Uhg/bGrVpKfBDIr6gTREwTBul20OR5Fa8qWRDGfBOlJKCMjJZF2OQfNvBXgePz/sDX4fh
9up6DiaEXd2i+WaII/2xWV5B+Fa3ZW8v6mLSy68ARgGknMCSyzuuCwTkLEWcAQyV7aA4eZzLbVgn
CIKw3FjNW2/6RavO7RrRKtYAlUZikYsTE/++yCvfwpEMF6IIgqlOntGL5u4h95Dn/EBjXXaRs9zS
v88PJQwnzegDwjhBCE67C8nxoOhLGPI3+FUs7wyvpLuclVfQWzeEQCLFjtlkjCQbUXzKOTkQ63ME
cSNr1AjPh11lux+o5gSo6/FkvKMSy1vENflkOVkFfY+17efL/xCk5jc9a2jll6a84UK27bKVEI4R
ImybKe3ivNiYhhhLCxG/fSY7NBMePUfPB2hAT2eK/GSPg9CPVANYcf2gYuKogAxGcxiTEF414RE5
smsD96gTvtNdZW4pyyI87rnKlqFSbSCuIpAeaSD+9t0Aki/dskGyUecdwY0snb4cy7EJVXEFeDMp
/piF3x2XBTM/DCnkbbrL8VfpubvahXE18dcskkmg4GSiWErmGNVJJcvDhI3uV+HZV04w9Kvl1oBc
kFEyv55VzwUgeXirloo7cN/eMLDhEzyu5epVUTD6Awr3vISlSl7/MCeUkrQpLEG+tDvSV8w4sYVL
zlqgACXNlx2Wb5JfvfRcmfi0ItvTzBjkzq4sVIHHGse2M7cNNNspbyk30MtGlPXHf/dvxJfknLN1
nUcar9E2CYtDTHSZOGu40GkXLTizAOf/Bzvfq9t0Gb+zdCKmR3rwPB3G1B+MKZBQ4KI2JgIxZSsD
ehPX+j+J9A9d4dMjHgxkDg845xkLYhbZE3H2tk4FsbZa0J7IrmGXd6RbOoEiws4obH8ogpw0yLnK
D1Jc5DL6m7qPk+DWCkUNjuOcGTwrDM1Hs5HAGwRQVARrvlX1D7g6V8qo+MyekkmwGzmaUKycIEAf
fKG4m7xw2vHI2tL5vNIZEDXa+khyGaACixD/fNG4at4VlX25TR8jPAQmyqRDrYlNye350F+o9XAe
gKSA3tKCZvPt4BGN+QFGM2kl6/bRdzLVwtFbrUl9JoLMu2ER7JK9r2+03rpab4QMmhVdGnD+c384
kUqqzrd6FL3aKjXOAZh4g69IB8WwiafjWcpkBf77NHeVUdpGeMnNgAEmuM6pJrjHWrqOlVXT1x6V
lw/pvrwyN6J49lO3jvzjOP1fqwZAQKgzdu6P/8kEUbVHc6OiqA/eQ6b6FzTzdLWW00cI37m1cFtJ
VFnl6CjEvlZFf++Rjg4vSyZBij1hXsaHu88YDR9vTjoRL7CsRn4mpXN+ovLtGDkYpxYv5fPAlJtg
v4hNR2e0JoAmhiMbsZWwwCsEYJncGDwBxXQJ38QD6YZpDfzaI1beafTKPq/f7rGy9mxMIerZEv3r
vt0QG9yvRIictYlHsvB0qLg/GjGkjXRJ6wkZGxu4GVxkddnUbhElV1lLKTQgTTkfY6122rVskf8p
RMKdRLkKCqQhPoGcJcoSWH0rzChMOF3UjWYENPBCLnpurk32AMV9HGKSXjks+JH7HbNUOOaDpCx1
X0OItQ8qD/MhHgtoinR19JD4cWZt05c9daVIjgmd7pJmhUx/XjE17XsqwL+svcg3UlJgnXdpAvEn
BCPKWEwXR88sRh3O2HkepPMAluXxL2w/xxh2INq1rpEjCEj2/ohe5lKJCI/dsMfkX8ceKgCJl6te
+67I6V4V3sAJrYvs6AynhFkhz/dsEaKou1LTvU3/ndU04lCY0+tfHoLO+pmJ5lJ9fcMbPT2u6d7E
/aPD+9L7qgWBj3FId1CW9GPzaxXdx4ZY/Eh/7rgUDydjVN+LLBdJ+rm2mXrbuU4r499PTP+6Jb/R
QQnEUsW/v9dvRpDH7DxWkzenZn3HKITuBW28gNMLMI3P4NgMo0dNNV6Pgb83OX2uEWG2jQqo4Dwz
VhqvvMuRcBug5O1xyml4WB8b6DSgUyK6wy9M+n+zLnu81JTOzknX1xYyuFnq4rIpQV45DVmlWigh
MPteo7/KXFOTGV5kSF9Ku4XgG8165swZVZZHr/YJpDFdj/95vxXs8fQ0n8patKtbmvsssu/eRJom
Vy5eHwRoAX6dlYIps9LynIBCPyO3n7jk0cSPp8PUbItxqMjma+W4V4p5HvxM5LwRNFkyGbb4z2tm
Tc/mP+ve06ykDo7Kh2KcZG2ZiKLvR+FQUaOH08aGs9GVxIikrYydysPZKhXUUie4fREqrlYwAZCX
FWMgbT1Wvatr92XGbpD+IC6ARRvmJSo6/rRuHF05+G3qB9lfAcGKxrrKodXd1si4KH3SVjAZ6NwD
BGfooKrbZzL8zfP6K2uwXuLkd5wVV4gut3rufFg+899pPj6PSqCdxa/gzBzrt/JOISIJTvzQy3UP
D1KzmKgx8MX4ceaegGfiq2bpBKqqlNox2Fn4PK1Z1Ea3/Qwn/cicQdRpcIEGpMtEHUF1/odVhXIS
LjZqp+k8dcER4zCxPoxaYKy4o9/DCtv57NY9OXm5xm8QyqOwqSmWF3PXhYnHNXK9HGcQZnZfoMBR
yDlWKVCIG2KW9jxqul7MEVGDh5LYyXRDlS5bFLaQ48WxuJgoHA0Q+s29Udrh40gZchG4XW4tXPt/
+3QeFlUVCdga4a+c0ZxWIj3HhTKRwEJP/CVt0JXbIbMp5Hfne4cmzDcRtvHvM9q/pLT1wyR4qD2A
xJwfbT5MV6YbOyEUT79T9KQBiTnU579L7XXwFx4fEs23tJrqszquXrnNZUyEtsJSD9vxKKOm3T0P
F+Vhe/eBohQG3t97gzxRThH1AbKkEMLDoPzxoIPnPEjShH8wXobAxjiBB9fSG6pIp1W66815dluS
4zsVl+YlrAsEO5bSvipARKXJsRxMQxPCdxJRWzbrFpxPwBDXad2l/N4QB7buOMBfZ1IhN1uLgo8O
ZbLRnSeuotBZW/pl5C+mVV07F4NT7MyVAihx7RFEalX3uclyKNlKgMvTeTx8fvrd61gtxYcW4m5Y
BSLeilfW1Q4Jry3gdii7Rla6amGx2pcGnUl3O22niVr9sm3PzP32Ny57oYFcW9iKvo4wggkXRX1Q
2XP13XzRkPbbJpY5jmg1Hg09zm8lLapiVr5xHd7/nfddTK2OUnhrI08tnAAocUeyDtdSI0xiXbWr
08SRwpEm7IL6y41pfxMH44Yk1ymDqqTsdkHWDNZSpNiEGx3hE7x3rZWuBxC66+hSCNuUuT0jdUoT
B5HnnolqURNTeS5YONCiELOYem79dmpnmlTdOyF0Up3oelAFmCxfyex+V4cHk9647DdHo6Sw3gXt
AWpwJBgt+VgUKIkQHt0v8lxLpDCr284FYIL4OntDsMte0UgeoBb1r3haQqwKoWMMV0cgbjlpQbat
9ar5Mmpbw1h2/ZhKs5zShuBKxWgOor6BMQtamLZKjCDv1Ok7tylAvqJO3lXrSk58jPmA2+gGOKqZ
QeEV7H6nD0UbBhsZ5aILnSP7aFzcIYeKuZCYP+2TTAthN65+KndmqsYDMQLrX6TNyom5fla7PFmQ
8nD4K0AovCl5A+gb77S60zuvR6NwSzIaKTUcuTz2U+4SdclqNC8gQum/x9BYFlinuWIx/RcbMb49
UZj6KIkGc1eJ3iXSe4kYrt8LGj19aoZ9QaKW3ntnVXr5jcXv9tEuJB43lUsLiacWFhpUnA0vy1B5
diuLLs9hcHE7KtSFSaD3aGcBN6b1T1vRPYb7SRyqAvET0q16HbOxIJtUfKyATRpaFtJ6UKn/LYvB
wtouKfoX60LClBZHK4sP+gOHCse4SyxQM6aOPgfh9nDq1aJNEUrOIh1CTqR4omhHQIUAXzon0HhL
dKjTc63h0vMHaSIADLfAH0O2v2FOt+qsqropE7oQw/hvWFn0J0vOXf2AQsWPBE5HGzdhjGG409tW
2MtFwqZCWpnZPfVQ4CT6DNA1jFidlCrUjxaGHFa6vOH/EMIW2hMyz3W/kS0+Qw6HyN139Nfg2uJZ
eLxSC3mz6Yb9ljOb785ZZ6YAFN+pxc0RLlZC7x2OwWqDYX0SQtQO+HAR/CPQB9rbT62Dr6ZYaksd
NjP0eymEVa5BNuuNz9s5ir+gqU6KfsTy3iBOng1bEAx+YLW9WSN/R6BN1fw1L9PP9qZfS7gwLJ7+
fWtcGu6av92YDJN7uC5FPf+aTFFI65Un12rQj9FgLFb2kBOLsrCstnPX9HoBbJxaypHdMXOssyVx
VV6GzwrIi8c0J+U2yEUvYFcBruZZxPSnYIrK4oqjc252lBZ+u0FlOOyc1M0ADf1oU5zbYsHcXQxo
Z8gpwH4CJ8BAH0dy3mkijMKtaBPE7jK2yDDK7gmZJpklHA6ViNbhCSRw8pa/awVPoe2TpzowY7gJ
fuzxBJQrIyc7JI8yYoz5kUwIwkaL5Xq0YtWrnoeBzW7hWf14ZW8NuPrdvDkww8VGvLv5OkPUg5Np
+D7VbzDRIBug5l3SDKYUx9s8WmDUauuNBUEUH1VLOGS/NTZNZ8bLYan113AGKJ4WGIVh9+jsz5aO
TsvCNaK/at0zpMd+DXLrLjFMUelgcNYPqxLv755DhlqXp3I3rnBGNn+PQNcnsNpRyTWwQIioN1aA
aI7Knkv/KSdQ42Nvd0sPw+zuS4vSUuW0hM6KTXescjX1t5u2iS//Rhb7h6tL2Dyh0uYKxAdi+Zmc
QeN6+SFLEE/OAIzPnFziBgKrXZC7edkXVHumbZBfFR3+4t/+LO48U9DjN9vnbtLoM9HndHn2B9qd
UoHhuE5uQDdD+D9kPMTOrp5BGD1mrq2NNokcEP5GwdgQVAfTl4nID2pJRjxql9IXbLCGCuOkOtzU
8Q1t0PeeJDf8x9G8RKQfTJ2S8BGvVfrI0qW55DSH/FnqoPUqCoAjhyZHNxtDfqog/i3+7oreMwKB
/cmWdlcbLPDB+IlK7grvrz5LHL1BxoXDs+9vR2kPF68BCmOUpG+VmYMyi5JRtGsO9YRC9YUPJY9c
POfu/kUh2W5J6s0Of+w/zjGlkRFulXBNOm2pANqaI8koMkr0fn1+qPHl6bVi6fSqzn5kwKU0ksmL
HfgQ3k8KJuDQ7EteR1xvMOwm031D9rE7vTZ6P8a9UWnR3xYpL8V5ckKC91F0GmGGMW36LUsDEEUw
sieNHeVeqlAyEaOUEiG9ERO1EElkjX9y78zc0GidnPa4w2OVCcCtj+D5gtRXq9FeWPJZMFXllUGA
CW/UqUFcK9KtZKBuD09B9nxYKx03lWaou9oQNmqnFvZH0NwQg3kGkad28kUIMKJZ/UWmHh9yAqhV
9ACv5y49okvl0VhVq6vdbPbBS89aMj3j/OTp9Q64/tK7sAbwQSfxdykwuTEge8TtIH9FEQEEsso8
4Na2gwwjRAWl1TZqSybj1l0urHhx9T1l4IYzrAm5etWu/kSioJEiGdNh2AZZdw8CHi5BORJL/T6z
KlnL7YJVCPaEl4l5pWnS/DvdVP0g0HC35KWclBGP6y7l0GLyW+bVTXwru2XaBGkkq7tzK27XMTwf
fLGz9qDxvXIamEZkfeITJZG2QZX2OjHHzq44STX9oY7sygUcbsMlWGoJoy5ogcf4Dl2uFh9x/UjG
F9ciixzt9IcBN8mb+HdLGuz0rxDsP1PJWrRzIfT37ZRinqyi8TPmNflUoNYAm2eIeLhLM83jcl0Z
e3dnBo3C3qnzdpEEjxJN+oh3PV0cCUpS2OSKakdXqC4OMqIkWkBVwOLDQLg+Q96ftulteQj+C8XM
NZb7itO4gbEmrVVdhRjaw5vZspv+6UCn8K3TPX3CEczl9EbIczHvUs56vZXKXAFX99cpcV71SAge
q2t2Z2/rAj59bjN/3d7JjpAYA28+eGiL+CqUHl5Nd5sgb7930/3mm9qZI5szA5tD7dm+wPDEyIgO
6SmKJ2CIOmYeMfArSdL+qQRATpZCNoLyGCQnKebYFZzU7AwJif4HOyD+6PFdSFcZBQt9fNwy2X5V
Q7BXsHNZSeHOx9DQCljQBSBiZIb3GniUbUkrRIEoEOPzbqNsahtNGH4BKmKUCy8pZx4hjzWdmL2I
UrM+nK/YtzePUZIbQiMHLZweYlBQS9UYNBSmXeHi1yRgzLDKYaRn1VDnykG8BTiOFfzPBfdmLLR+
Ad4T1LM0dvMWZVXJf9bNzkrediY3pp1IDGnLDD6FaO1Wv8dBkZV69umD8A2y8jWgBmWQ6E+7NDts
Smmn8dTK2VoVlXg2/vxXPoo1iQc7bRvZIqt+dmiBA0zNmGj9gL618e3rBUhqwy/7wUG/4AqhTF1W
yUnKDXlOkVXsf2GBv8mRf6n9YDwJyFOUMKGyTVAAKC76wt1HKeRUolqDcSg024osx7/VLVMoe4Cm
+AN9PGp4kM0OIPp3n3xzVZ76J8w5FwUdBiWi0GLeMU0mz0+TImzsdNIETxs9rnwJXnmPeiaDr1Xo
VcOALfWskE8PuDO78XyZrIKhn1XJGw3xVEwMILdUi6hZ2v87jFm4I+jUHpvML8R2F6sXzvUpx737
X/Q2nwxH1ZItb0/wkauqSPsNQa/xFWezvmxCS+W2cSXCIQBXWba9jUiI6J9Rw78wyhDFZUQQ4NN9
ELQdkq8pKF1FDMs8Y9OiGHQVwjXFuDd9lCZJ5pIM+16pOdJZOHyz/roYUv5IzY7ieRg7Adxntz4E
plLdrZZHgqrRBrC9hbN+MPPxScOgFLb9tVoHglLxZqKTfAj4HOJ8nRVWOFUYFqOIheD/Ytj4fUGH
tiL4LSgl1QslXsiEvx5yaKNeY/gNx7EgyKX5F6mU3fb+bmCSDxPHHLZVyMAoBSODZLJi4RXhUpy5
zz/AaIg6SPLp366TZgloZ/0hXNYoKPiGXMGwyk8JHTprl/WyNlZNMIw5atg2pwrqjjT3ETnzZ9LA
muPCKLr+GQE384vklQiBWLO6XuuN/8YaQZ2A+Mx/k6Vb71pjpwf6sHuUuBPLDGTN6iOmYI6I13BR
V9arwvF+Ru7x9ZqjPZJbtgzlO8hODWAEDv1ZbrzieYRkIIUj6oMiSPfTKzJuw3HLaw3Bc+PvidJI
IG1cuB4KaD+x4HAxfRkmuFB9ivlL/qRp058EtNtcQR7/pK7/CNIEWobA0TEGADsfGXZsLM9bWu4q
UGaWTcpk0hyTTIulzL6dIThzL17gEzPjDzgvaHYIu2kkqqD94fPArX2iJjR/ZHlfBUBi1nqK3KnX
PMd2C1ZLChgIdIzDKUrZ28hYTrtmG+wsczyU5c99nH+BqH2z/oY5skzxeIHNJ33bqsKxS1+Yp3D/
cCnRXwvxBeurS5PYM6w3x8uAYnRCv7ZzRYtAZ88Cc7ott238VTYIibzD6vD8mZwQIjF6Nq0xT/LY
SmZvYUhGelHLfZilcYYtr11LazeW4B4VBobmmTYmg9ub/C1gU21f1HE0b43XaZO86oL5EtqpOQjm
IxMw0TatNaLZiaJyMqMHGQ6qwK3n+69arr2e+3aN4YKzDpgpb5lmCpJ6QwJWliUEzTgB40ZrYKF4
uq1xGGVxeZKQgbgmInG74MW/nIQ3ewGC7KMRvaX8o9folaX9aPmo6IoS0jNHJjDyNPM/Ukkiomke
3WJhg+EKwqFuaw2MIuLWU2wMRRE+tfnHXQt/dEF/XGmb9qtsJkq/X/HvuHEvUs2I333KWoZl0SuD
tJ+1O9cjAbLl6HVV93Knpk7J1N8RXwUkRMniEk1MqqgRzYeHPcrfeLJ0U624YkDipW3qW/pUmO5e
CpygE72QmPZHU31iGPiH8I5LtmRov+az9ZacIOD2OxUut2qaS66R/ErbYTpLssbGzYp98vcoGMOE
bkutajsit3db5auXPzJW8nYPGVlxH/LoVJnUhdyOTlsRh/ujB50oTliIJw9/sWLKOqQ5golX39sy
5G1xBN3pdT6KajVQBxiYh8Ox8rHv/+s+0QLotuQMZkscdiOh1dj0FA/I+imuiN/fxo0+qnrPkrOv
0UxcC/QSyp+zjBGi2jFpqIHuLDAlw2OEJpBI1bAPmIU5QkozM4qtijLeTVztlllR0jCGS0Y4o/uv
1qAKK7o5imtdp5HI
`protect end_protected

