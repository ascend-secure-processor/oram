
	parameter					IVEntropyWidth =	64,
	           					AESWidth      =	128,
                                AESDelay      = 12

