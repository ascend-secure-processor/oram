

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
o1XvyBeyYUoQDOkuIN0oDJjvwiHFFX+bswujaMpyJzOQlV1nkjT27C72UqkZJvl9s7KOg9k9Oa0C
5fzbVCEAJw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WUHHSycD4lfGHQmYkeW5jAIpY/pS+Oa+1kdJ72e4/EI4GNhwFYqpLLMifP0/wWKx3SScVLyx9Fkd
Y9T2Z9ax6OOU+SBjgs6QfK3u35fGaAtNoauEUEQ/gwBrfb5ao/iOnNytNj9TSyr0Emjp/2XPlMs0
6KFASJInKpTKA4bSH5c=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
6I8npnGm7xIt06lnFk3e1mR5MbLVIm52LTiNl/E/ygvPk3huZV66seOo2ogAo9G49iIqP0UhwWSl
q412vt9tWcyqlhMGIbafpkYonbtRtwBu/kAnMjkHr2on9m/5eYlHkT4bAlnJq0vt0ASXOMZyLvsG
G0/iPf8cHHMioupJAawSi9BGa0JWcJIUamOxGWqLup+1FsG07TTBZGHQ0iPIA/2Rep83EZ9B9o1r
gXQ21F2AMMycqVgABeZDtY7HpNHGYD7WUoCNomjeNMWtbxR8gBdx0SkglWprD12Tpt1Qd5SR5NBJ
P2QB4qnzk05IOXLWvowwsUNBbahAe3L8RoTf6w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o+Z9UY3360k0KddMZqfJI0r/8nF1YwH2Dz4FkvMmCdoJGy4I0qdgEw0SaWcYSokohm+06YcH34JZ
QtWktTnNUbv2dk7q4KDyoYKNLC+LuRoHzm32TI+7Qs23AaK35wiEDBTyLWWzB131xMCgD43HTyA5
zwngqF9Nu6KkAGintoc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pjc8e2FySm9yNf/MAbDZld9020UDzpMgj6rZa+T3xWltY7MDrzySC2rP2GckhPTpRhn51Stm1PNd
0M5CGBu1A+H9NUOzITEPvLpCl8JAy/Jxd66lyywunXEbLC0WaCSL7Z7o10ZYth2wO4ZcaFAmCru/
xMBUgMaTTDp4mkVL8o9V2P5vVTUas+PdS5cwSKGzmlpzXq0A/f5geODz41VcS4gSWSu/CkiAQMtm
Y9mSGWhhtYd26rbMVTKO6LdKE2rBX8lBW5UVdSCOyZGbZR+0MkaaN/PBXaUL8kxdJqayjKW4Ko08
VM5Oc/WpltIAF8obG84Hfut3h30TZJh+B7R8hg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
MzasatMf96NHk8eu2EBJHz/zqtmQPXKsc1gd05fxAqQiyYgzO+uttsf/xlTY97vLwYFMBBPcX3CC
oXDQK+7VFe3eJGKsuDwHb5CWgfmxTJWNbnsSdd86DLcEHpPz7Y/1r4Cg3t8vH13DZvXK3R6Z3Lb3
WO3bKoywcQpf0BlQmzv5jmzVf6nWXO03/p9m4zcOGabyzk1iP4qRIocf+yp5EsYdGfzDQubYs78f
pxfWmaoQg7ZOCcHSZSKVIZ02D7RIwUEVBT0xQTAIujsnbaC2SCm1uMroZYR9UZVXi+MpZolcb2/Z
C17U/f2H44o7hQVWP19HnlIYikHDbJP8/XRF6tWZZJdKUK1DWHi25zI/MHrH2/NuAjeYakE+DC8B
wLWTy2wfumu96O+H8anGts5wxRjcnGjMsXivws7lcFm4TxDu22jmT7pVbTvn6X8eVtEWrgasHQ2f
zk8mZOL6pjb6g3x8uovvThaNZjkEcpFuj5dAZ4DINpVOZmSDd//rMsJT1eMwFaO/7pQfpQzvjmjT
KcwP24v7l2q/tp++diWlW64TYSHv5dCUy8N1iksXaht8s0NrBdwG9AqGlfKoIsWGWierztlpxvmp
myO18lN1co99CflsGl1cByd64DPt5NzV5mgKXwbNZyJHxxlO6qlnvr1h0XU+ggdjONf+xxCDpQNh
/pRhIiZBBv5dMDNpSsTVv4ZR9IH4vLm9/Eg7BXTlpBTssIWeHYswYnzRF3KMmgeyUc8+D9rlgU7i
i8hc5JXFCbT6CKE5V6uwlXAoG66lWFmygRyIA34BhlZqKBbKqwQdJSWNLRNP0X2JFqbQUIT9Keb/
BdRkZhgGUDX8eZgGYC/dMxwDvXyvTupV8NU5T9epyYQLkdZrgCTuGgMZ8oR47WUmxs3jAcGr88Fm
w7bb0nyR859EX5XoqAWzZETf+eYLwEpr1TuUcOEL122D2tSf542u4N1TPYqQwZgdeOlMLptBpVlt
1pam2S3N0xyULH0lr8UrT2k4B6XY/xK+yqvu4BLETXf9wK8K/XSbMuxK5wdCYNN3TAu2EiRqArNA
hxbxJ0495tRYxp+sHMSuhvBdwScY/YWB8css7an/xrHJG9nNbiopM0eTZR9Nvptl5Z/vf8YVwigA
TE9KLb7g2sQiDQpvk+4cECubQ8SDaO0xstq4wI3KX9yRGc01WG5HD+nOf2XZTckdMnyIE0GEKAam
oev4kQM/c2mnyNBqzzGlU74LERBWuSBOCHdXt5l50KrMfsD9LwjBaYmqN/HIwBL+aQc/XT7iYa2N
vvnMhY9TBejbAxkePOtthU7Ivt+R/mHI7Tai2nW40OmfdtRy91QOUTLspDZrXEaFPfLZImGUOTkm
eb4llKzACohtPTHRXKFsBb5liKSeFH2Q4DI0qN4IRO4D1tv3yVVA+6PPDlQ2Tlp8qCSBkNPX/Qr2
cZyl96b/a9EJlj2W/DSItGuvThgAx3qHx67XniyHwg8MCR2sC4J0HhU/Hmk7z7wpKlo1OdxvE6T4
7UHzdPQHpPd4JEp57hcV4ofvJ2Y+MUoUh4dlhPXjGsc3ahch2K0xNDiE9dir/5Pil8seduOOCfh6
Ekw/UBsn5iIq3uj0WumIXry/uzzrLtiSTkwG03LQIMTwh7r21qJOzFsQXUMblywuwSoPsIu8KcjM
nBGceDWxmsROtQbWulg7qVXzmhrXqtek/jV0661XjrG2R+iVykqTGI3YcKXLBVkh3WVrfSvkKoOe
sUxhBfXr7eXGlQKsoc1VU/zGJqeqIqOnEYVx1fNh1vIyH7TQtYMZBjlsq62JNUNrwejocBYGuXQa
a6yAnRvSKT2dGPxDkmrx7/Nk52Lyqu/3sE/T4ez8cX94QtkHUAMs/fSBncNQz1dlDNYMTb2SSVIy
nWcYouw4v3KjsFP7Xd2ty107ra+tKfMT/nsAtbGXC0LowrGjNp7gPMGh2BHxBG7P9jbjjTSR0dsk
oJ09TAMilGpDih+I8+1hydRVEYXe4xZWSmh/Oc8Ix3LLDtUrCwmAkz6kOknxJRwZpeaGhpqni9iX
MLHUGBn19v8xjfgOuhwX8treS9/8WRQWjHtr/KWY+2qN2AeHYD5PHmll4kMU8s0TFV8S44PvrQqa
DYEm+jxSUOnW1lpCebgKCBFPzEK8YTzAoz9YDfzGKBC8aDHxDiroxLR4ie98KwLfBhHpaGoFQtZD
YV94jV8US1HQiKrH2Db5skO3SjRpr0ZYNUDZ72AsZrXzDDIURfObsMdWHkZ+8LVJ0aevz060IX0K
5GKQOfNkLjIyD/oMNU6+jjGFs6ZO4/F7rffRyZJ1yYL/8U8XWI2uEqfmOLlj3fp4Ut30uLFWJTh6
SN8KOUCraX7PL2gbF9TGAU4I1MjOWWh6jN/QhDaXmRiUdCkZamlFxvAEYRLLNitFDHZR1mLX1wI6
FLOtdt7Nz5dP0AzQVUkrMU5UPKcvQutBp2fp0mOIAhLwdgrxwhvP9OJsIQ0kLIi+7HwjO6gjCdBu
UKGs3zIJMSxUc1gM0QSDPobxeJb0KF3Y44zSAre0S/dKnheYn5Lp0/DOM+16y1YZ4+atOVYtNpKQ
aS/iW1ZjyMeZKems43QOedRQouvp2EayAo9oDFIl9dT/IfzZZ2kx76Qsj1jNGZGmdaprlESydy1R
gTgm54WrlJpzZhVA6W8DRSgK37Kks0Et5MQeaJSYiByqhJhuLjRxmI0j7vjhSHZ6GjS3hWxtzRjy
aBevIxdk72aUVjStRpZBnjGvjAAxxMQHQ6H5oLZicNnDuLoyl+COl2ILO0R3hobSg+bPdTmDbn44
aT+4COChBLHScf9JPbLq/dYgdngkE8ti3kKvGDe8wNOMzs0X9oMShbiUE4NdtQaqLsyzC1Vx7n0C
gbvw+VAEoJAvp0Dy5cBQwwsunXoX+CgL8cv5OL4SGAHiXC8IZpf6/sBWPvRU7sL/OGbazUXvYQwL
eHuU2AKByjO++K6Lc5Br6DWaFWc+0IZ8EX0zstG+N+SDr9M2QYgR0UQU0S0src2+P5fiWXL779eS
uqt8JDRcGGsTrFiRBjYcqk5ESNT3a/cyj6de26HWw2GsRZg5gUsTekkbt+vEmK1MNBVNIaez8wVX
kKZZRWMzzHNDQ7PTkYaqJplsHCuWz/ifsDz+zks+QKdg/Xntj0c5bFFBHQiHBgX2b00r+7L8oB0M
W0w4NoEe5GbPkntbeKnJlTwCc3jzjRxiddyPwK6kKHPAYVmJTrlOnbxnFWlR6zfN9c3j0/qrU78q
0e1QMnr0QzyVwedixskjFd1RbJuQqrpDfqgQ67dfxXFAtz+ML7+Juzk9kR+Anq38GTa2camPvQ4h
FnmuWJIRu/rPyDA8EjUifQlOCkvZQ2pEt+UaLC7oo6mLJaU0+Q85fP0idO2PqzGSdzD8tMnWRvru
tkIyrTEdXvxByWqLvHIIS2/uQcP7NQNSaYRtmnB7LdPs8OwEkM8D73X2GIrU22E4JsCiHRVIFSS9
PUXLDHRJLgMMeIIIf70HpKEV5chqsnZzcQ5alJrKNyoFY85V+UTIkHJegR/AvLPTx+cX0GtM7oen
DRB/M1OZka17K+kj6pTJVaph4N+5lkPCp8Tp7YHnvsZf8jL028kOTjinYC+Sr42OfEcO7W2Zu99o
wzzUmmPX68k1R/d4imZnIAUezLSrpUtWCZH7/JdzGIBSF25PRyFQfffFeBY/F23S7t5raRSpWiwr
QeHLGuFdXx8XDX5LN6u+LwlEO01Jk4NbjkaLpgrVGn6yHcm+znK+ZFvwU1jIRJY9qBKx/nOM72Zo
BdNNX7OCnN/4R1+Q7swJxfTKSKfGX//HAWnCOwxhOjquekc39fYwio/JyHlMtvI8j/tyDMsc1Bu/
fvKhYeatwhVUc7RdvVdAw9xI9KdNqHcTowwuG+dvY9DTjAuVDiH0he4MKU+hP3LdD705LcJgLrWn
Uw9g/QLWfyFu7nfThY1wpTSLz1vw0yK38TSIDM7usDD6Fu9R2LCnMud/WPa+PiQU5yUmtOJSr6Az
p11dAGZ35x0+H8YCn8BIxRId7BKiJfKebIoWOTKOumS27XFaDIOF9DmrHa4R34mLoS89fZyg65tA
7mMKKCTCWh5l/76QxACn3JeIiQRskedCsk6irT+6cpqV05sRKdIJXCHtFgeXlXUNYDfNL6+CyT4d
rBrAa4yTHIYf7KwCDwfVwefcyjrxx3eS6vF6cAPfL7+YEil912i2mYydg7T8B8a1WN2brOccX6sz
Kc+oGvS/35qaJ85jo4ivrIFTp9V71caQP9U5221YEbjERsTfMvEe6A4XJ7lXr87tfN9QysaSQvrp
Mzphfm2Fp+04qdvAS9cgQXUNZ3Dbsu/abgYfsoe4GArQBtJahMn9/nWgDjzhHhMAu8QlzcdOp5Ub
8hloAwUhJoVk7e1btDVfUNSOzulJKCVKC7Efva4l1c/tvpOTxMULIfRbw6W5UzE5K+opw0dVtIWv
H5AD14ckZxtNEHKDxfM82qcpYS3wOIX+voukgTMUVi9hxyIfgWXnCj9PEEVoNE3DhJtQhLnxLODN
n91IirMNX9NRQhfI5DF8HsNQ2MAqzWMAUHAxJa/t+V5L59q4UayrQTNIw0aSdO4BER6cEthecYC0
f3qDarY5PMCTJKIgKRAJn11Z5K9xVDnKvyMUQS1vx+iSt/2u0ksFp4+a55EDbZm/XsNZvNOxFPnR
kbjl3dXDFUjn7ML6nvbLzdfUiUXKQbWIeDecIQygBMUPhIhIq0oUIrE6SxBesNIbb5kK8c1Lz3DN
mgF3j89C+nhoBLXNYR/1cWsknrgzTMzEzv5yg2h9WRC7DK26cxFLi3W5WDqD1ABBZrJfRu7zLRPn
IzsnBOUAkXJijbGl/DXOvDkJnHpa+fiJU66mXR8iNLyxRmD1BTY2/7jICvqj6MaxPuEqlDGp/38M
xfNG55Eua3l0Wfa1G2uvVBYYcGTJU1lWjDIL/qas+5LJ+QdUwUJ/zhWom2TaevxHSV/lvVxwxzlr
IHMPGJTEvxLM51FjcYwVCMD7Hf8O6+lhX3c96ufnQX/SFKIlDAxn14wdt4wU5D7Oqrb9jfsRJm7d
GQCIgIIUCPyzyrK+MU9qw0Rm4Ex5BpHqmPRwHIALgWUbJdPnzFD9iv81DJCyx0wpyGECwNLOGAAr
9CO4qHI5Xe97YHSlhOcIpMRTwlkXZuUztFz18tGswwJXpw2YDEOBKYwNNFbpmcdrJV9vqVcNnMEe
IuXFCXjeEHzBfJDH9L2kANYBq/+s6a0QlMzRhiyQKk+SuQ5cqLPQAFBk/gKrEq/fvRdm9ySu6RLh
pnTAe01p+NrWMevdGUlCmeU3zxCfi4FB+iU=
`protect end_protected

