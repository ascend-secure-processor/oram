    parameter   LeafWidth = 32,         // in bits       // TODO is this just ORAML? A: Padded to power of 2; TODO lets make it a localparam then
                PLBCapacity = 1024     // in bits
