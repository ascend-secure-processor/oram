

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fURN3Zq45stNmPJ5IrSg558z4RMDyVlVmhpcHoBFEqHebUEHfGFMPVaL60i5dxPJaEkm/pacXdgn
/hPz47mUqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NE+vLUxN+6YACOi/HGEvILmbo7vO6LThzmb8yL+KwJNikvJgR6XvgJsw61mSrG/vhcyQQh1n2teU
93IgiadOAfQelF9ge9UOfqKOPnXd41WY7MXMbH4k2zZVVZuNKhzrGRptmilMY2MERM+LXqERkX/m
yUhz+h560RT2vxGT1Hc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fNXUhAfXYy6/HaF3bzi0ZtYepC0Jn1NjDNdoFSni1DXhmqvDRWVvpIk2shxxj/yZec19Z1twrJOl
1MaJOuHzSoQMRd1SMK8+WFx0CSOBnlOtTCqmJBbh8Gwf2fctcbnELLGfu4wyLZ1XrA/vEc5V6ZrQ
Xft6CUGWvRanStEUMjaF7W6t7XBaVk+okk+YcalulOhZdpqZ7pdoiYYjWjwBg0E5IfrgwpGOuAdo
ucI4FlE1Li7gbgq0oG7uYUz2YkY2UI71y93kkUGHNDe6tu/27aXvHpMiPaldWy4JaJVMFk0Hn5I9
P7hQexG+6liDXwBJ1RuRw+0knBBvf4Mjcm5EuA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TPKU51+omWWDLZMw5KpovA7iViHZJ047vxTifLnOlKJPQyQv3x/JRWRaTxKZ3f1ymLUZt8tK+GHy
9Vx8yo9MIupwv8aPEN73CF38TT+HDQSG4raldbWXu8L8hswlBW4E2iWRPFMetnqFQ3+Gzf2pt6J3
AADDbPYlqt3DmQ7lADE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j6/Kob+LYYqLPMWBLANmTaGld6jHrTdK78QmaYExMgV2m4rlm3L3YTkjjinSyYSOk1JhfEAdrm2J
WMN7JsxVanPhc6aNqRd3/KjTbvcl1AGY7AK0pnEF6RzvKVfZHz6/cKThd+09PDUGpbegNjB6rQPv
1QeY6nuyrvHfsAJ7YslWGQ0wWsreunRUwcnoeJND0Hr6+w+qgc85Cugsx4eJ6R5LptuoyI0rXWBo
M7ts/hzSAo/XRuOlPjohOqi4DFpQi/MHkb7cSrgoxAwCaGmFO2DcGiXE5xMHsoOu32ZkMksDKLsG
DMnnXK5ErFhL91RYcpM8ywjQxj1ZPe4du8bWnA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
5RoGP19S9JBABgs+Z1LTC2cFtAc9xQUXUKvRCP+rM+zyT/O6f8MBbduNZ0/TvC5pOdmeb3qvyYa/
kKJNUM/1hwInyBTPcW9Uj6q4eTW0EJZhC/OMpV+quVFCTUjnCOB0czkNZjllNa2ZFc337hVbuLub
o4P375H7yqzLMejw2+K/JPPEpVWPL7JI88iBnzc1uIfr0S4c3y8ZpOhq78q40FRZrPCaC+9zalEm
Dob7O1MC3yQUlcDMIPXBojqQrZvZqZRpV0Pztb4HYNozBjj3+mYKs/5g/LAYXXnicZ6lPj1uhNJG
gvEp5FEBLAENAyhJfzXaTiWzDlBfMKn9o4g/j2mD1ZrYILbF0qh+VA7f+0w3hOhB/Jwb9j2TTbAx
/zHOBp3B5oXnetjSe3RKFky8BjTeBh17e1qP5lpsx0PvhliR3CFiKYw9nWolvSwNAMZqlvnBhcrf
BfCzt49PfcKsf8Al4CBSNrqSPdHEJ/n3baDaNrrLVVtmxwMPQa0i3GazYtuvkXKZRjpom6pwHfOu
nhm92pKL4h+7LgWm37lEleohBBZoyAQ+cwc+j8JvT/dNgzBylucpjhTQKFBaouDgnUUF59LEKeqR
NcFp5dD4y9ojVWYN4/u7+4IEakTfs6d0atkSMt/fB/AYFlXUu83M4LyA1+uW+Snnl1rIrf9OBqd2
fCpjSFrgtFh5ye8FMUxfq5RHxX017buwm2R4MQLAaLKLygl7BQX1uMLy+XLMkBskByfRXL/KJY/w
UyxFO1yNXCsxoiAjwRg8ZCjXkjKJJpMRY2CxpnqKHJHh9GjmdkpT3F/NS3GZoPo6hKUmLvXX5nZG
2fl7qLPHM2Hqb2iSf5Bug4d5DRtbFqnuwoUvTMCcJRPoIFOONmUmxfoaAkjDJDeDyhBHcvdKpUx/
ADZjnUcnvv7JHKSx4FPcwgAHI0qbwzgXCoh3/Vl0beQBVRK6YU3xxQc9xbDNyFZP9fTEA+7SHgao
wAkXzO+EL3Sea1HfAJZT0zbR66pUJMYtLXIr0Bjv7+XASp4qLh8GagwOyPOPk3ZokkQ6zCKE/0KZ
E+E/9T5LI+KWKidCxpAQ4KKYEvekZVkfws3n/mWZgTnMMTBVe0iJY/eK0M6OOMRdf93c2QzJpKJu
eM9eIhzuWL0gOEbEyP4U10nbbdt6Q8dH7Dqo7YwEJL+APaXZUdi3R8QsQlE8A8sA7tggROnKheep
OyJnD0n+rAqSu0Hq99AWju9AqJygDM7YdyGTroc90CUTLpOYQNhWbX/Ovq182vxDcl1dwCFwJYWt
XA+Dpl/fUN7hbhfxfl+MfMvps86mM/LBjZfkZeY+/5M+SyUl2nwBZ9xyP7Te5Arii7z0Ct9A48Z/
1/6Z8PdJF7Ie8jycQb8ILfxYlBTREcQVB+ULkMWDlW4F1tYNys2wEErE8IejRdZ+pQ/VpViMep0O
LJoZXrNTBLDqGlsKOTlClrU83o0blv06T6QzPyw5Yd2jFKcYbjjOTkjbB86nmxlnjxnjNTDMyCzb
i+8D2tfOx7cs4TrPNRxdwgFSXBxzTMXi/LIqxflr/ar86nlzFkgSTwFBSPeTFeYRJqyiDbdCMF4j
yrusnwafZYCo/fApNByq6pc3u06r2E8ht9k5l6K8xAg70dgGPHearqNbMMrG5hPSraj3skNDMIhl
GBA7bKtTcHuxRRmuwMdddqZ7P17MS6mu+1paRV3SO5XgRD8ES1o+QO/s8vDdHw743s9Pm1d9Ao4K
1JXxcQ326LUfCHdG2m9L2Qt1GvtcljMHRXCQuyenKkbJHwAbRhr6pJ5z1dp0GksTN7DUH71d9xj8
+5qGojDC25a9SFxMva7VOxXOJvezzKXKjMOy+mVSlk8NIBhKqYfyM1411sy3g1vxlyzi3WEolGl3
0NILfriYdz6TL8x+fn8/1LvsHlvMtVvjyTePBbDYObjaN5NnYNZoOZ95TmPy6bJHFFNlKOZYYKm7
Zj5z6bgpR6B2PAliN2jSZhPy6tTN6i1paYy6m53xr0oTh/0N+4MJalBl4m+Kv4EuYGqH0DQHwylU
4QohAhq8eX5rUfsbE1wR29Mma7REV7U39UMSwr7Q+dUVxWJjXa4lqIyNR7bZRFmMwt8ReF317Dvf
Dq1o+8dKyBMLc0EramjYv/0VdchSvsA4O7JJzFC4Gf4vglv7OZz9d66qnHjQYZIGOiB1HbSS0COC
P+LLp9ElFHoEojxLCmZNL0o4Q65nF6Wmet/af+0k8QbiEvr5/otNmW6eOHylcxYcBpHjTTuNqiJq
QSLDuKxHD502yioXmvFWirdyna5aJ1LbyaOUhJVT9/gOJ6ij+k92LnR6EdVwmrpxC9/fCqV9O6hN
l0BsFI/AKLnwewb4B3kWx9onYvv/dD7p6SIPgyRjudVO+gsYAqVgFm38U+zCIHpQDsO0z4OZaEKt
0fxfgvKG33nhVdNOL7nuUjNmV22ILhNserCIl185VM1HJbNWdp/XEnmPjtU4Tm4x5+7hs7LOqdp6
ljr4UUkbR7vtoCVvvZEkaQP98fVo711NMwQL723XG6o+3n4r6imVdJoR5TwD2UNV/FvQJMS0NUr8
OS7wIQtGW4KGBtnoC2/dz+qH+BXtwaV464TXTJuU3xiE7haTDaR1ZRWXCJl0F5KxhoBNb6OHQCU/
yWwTag6yTsJahV4RZdWBWf1aLlBG71GueDLb4P7tOAElLbKo0u3D3Z8uanpjarpGI+kfn0w8ows5
0xoXLgKnkGb3Hvl9nzuNZCwv8kJZIMZC8I7+fMW9Q01Bhob/ULT2d6miF8GsgxL5/nO4I0/IEAr0
5Qoz264fn3OknqcR3VX5pfrC0ylS/LfANFAF+54C5mTLoPovXVD7IQL/3Vy0gCO7LjqvpD2YNtEA
2IttzOMUfpPM20HJulEjWWkHDCszsjhs5r+1HOap4WZrlYdDLXfEl06swGxVyOK39sK88HimHHau
88hMI1gC+zHARvGpV3A4Aa3BvNMRWNN363lfVN0c2Mxu9hNdumREuigQJlzxkmKe0/eR/XfqbC8C
s74LzGYKmyFm4aEjGkvcp/073WgTjE+bj9NHsiftwXqoaggHfSp9aVYy8cY4lkrqFjNv01UROUms
DjUG9BY6NMMawspJ8tkNVr1dtZqeqtRNIAXhZIInLR41vw6TEjlGMC8+ZFG3YkU67EXa0Rfg2Q3e
FhCsZ4Y2BwyhoQS2wK/SRlxD6XbLuo2Yr/fAlvewi3r9zYZXWiAKdBpH9h97PP05WL8+5OU4Vi+2
yjtWLSUcICZQ+ghxHT5qqnD1kd1wWFAatejDKIE9SnUKHHQfp21YguPJewBybvp4nyvd09cKsESz
K5MXflKTbEjSyNMxn+bUtWou+MvF9IPsczwqJUhKvTAb2rClJiQtKC42+cxLUETiEuJ8f4RLQo0b
ILrUxKcT464Fy2CQqlvgpEr02rZR3y33SrI7JFgBTtFeYn8dQYEpyCEymUMGOT/gekYDYwYn/yA9
jDzKauldydxI2hTjbB4b/1FRw9j/gwcGEsjo8CkqJudXgoFnkEkaE9vdj7/baGVXz5SzdoJgaYDh
kD4J9IyJnG2pkMoeAzpCKmAunEQrIxDv8k5GxuRHsAgShxJPa9HmDZwMUbCbYWMa4fg9z6RjgzRI
onXLz+IQoc85wd31R99rz55/GL3xzw377zj5Y21VvnQeMrxgVhPgJ2aoOJg4BqHcYlAPqGHzz8RN
lSFVb/ZNm9rBN7mk+IVt4OpETDfznBB4pjA+UtMveAOGfLSKUw4lqT15eEQxc/IbS68gzx681Wef
/CDLTs6QHTEdSlC8zGEM4GRmAHILFpSmIbKQmyi7xX9M+cqD6fwf/SaYuIWNYGfPXdHxURiM8pNd
wMvLzWHxIuf9gw9e339QbATGRg2RFuVfO0/Ewy/BP7RBF7oxi/bmo7Mc76Loi5tvM9brpkvQOtmy
tc+i3YUopbIpdGNFsf/KTlbiEOivFAwsDdi9/NJR6i/SLXDDTo/kFYehlQs49WMXeLe0WEM7cqpX
qMrlbBzbYXggmBphOr5Lec7mrmxpQ4zoZQsh6pFOvFJebjh/A8AaB7omB8BhGaLAOAJpQe3ONchI
VbSy6NFF2oyPVdGBIwttScx8p46gw/yWwWrbyPwiXL1igJkBPaOceV2Hc1Y7SDY+mDnOozTxIitE
nCNv8EVPpS+tpvSl03evZohGm4VNDOENGaW4MyhhZvGClDPL80ZchEUMET08I0M0RZrgIe+Mnn+5
daqhfGaQlKYSrOYjHeILvavil2Z2Ppbj59kIvwwAs6OknqmPIpSumXa+xZWQBvptRTfllAx/IpJ7
dVALUzmihrA3HtQcZ+EdwfT2iNy7k8S02IZHTlBbfsIYsth/cXyeZ7h6jVNQWdlcvnU1FDPUT31S
GrmrQG84Wzx0UmFACaXIvu3UH0dBxh0eEjqPTLTvKwKAm0GW8ujFf8Imapsa/RnYsRxK4Wg2Ltft
Te0mbzMxzt7q2NJFdrNKqJosfsFTbnfJB4tTjvnuUXsETZnFTCLsOCz2/A2kcLUbeI2829XkK77P
7BdUoRsGaloG/hUDZrKzCbJJagtlA0VG52Snw5fvfjpfDmIG/dcbiyCRQZfheovhPE4Q7hopyVF9
Yh1m63KonxWkUZm5vixRnQ7RS2TFPm2PYf2/9qXxYGDzcMBjhVj9aPaYlpfTN06fRZ63u/fEwMcQ
tqXxli1G5A08uuPoNn/jfMKgXz0bylc7lVI/w/Pc9AM+96ef45/wnUjlGY2RJUZlxjOGptDlKsZW
hukuJFtM7OQ6RAhOPY6T7qqr/2HBVR4v898vZaarrKJiG2fhqjD/XRTyh5WGYBAYaWyqTmOGiCPd
Tj77dejd6P2oISLkWuFEsXnrct2xUrOw1dDgLcJ/XnRDZu+bZrLY+Da0IIsmNFRUjb6+SM6YCwhg
lqB0WbL5OmO+LOtEOC/14LIowDCmVCPlckAeyVORWL6vcxG7/xoRlZNBEZHbHaf9UopAymkfbtqx
htykhKcOoQvcv0iqqMONA8fS4Ck3F9CwHlrZqZxaGb7K9OEkQ7pTMAWV74lLgJ0YP0wlcezm5fw6
CnqvZjN+TtwIbAux8W9aUhpUkMv1BsBQjAOr085htYMROEzlKRs8aNypdT4Tjqy8zSCAwaXSnsXh
S8MU1+kbGCH+7l6NCHTtX5oWdI0o6Pv12weR0wcG+5Ff8E9jTBAue8JzZwMZI/fHzWiLJdHKDpDS
r55tZB+mrNLdyYqcww2t33jAfPcMJE0uf7Yqa27c4LW1fUrWdzJiVrRAHr8jXYgdSUERIyRrZy8T
9VMwGUqRW1z6yB8cTacP7OtB+LXNc7L7x35T64ovaKDQ9w0B/OjQC8H8RfMNcLWuaXa6nMKaSaqv
WYoq1QAqnDEHn4SrIEKX0RITozZMWDLgfQQnC4et6bs6P9/BV9EInVuc6tNc0irI/9fLihXYC2h/
HDpb4MmxMqcTw8n5esPhueUn5SQatNbpaoAEYKjo4WKpS+q4zlfE3rLILgD8s9WjzQu0V5DO92e/
QfGCBtEKwHCgeQ0xwXEoo+Ly7XIlBpZVQGSzuvbe0fyqWVqqGppt3+imtptP3/hUy/FaOzwih1Kc
BOYoTORKb1avjCWzSpGn3iBCylJQneXgmXYxRsLc15O6o5m7eQtRJq4ccEZLSMyd8tNKzSYPw/7m
PPTGU6OE2yc3H3wCjxB2IsSc7buFcVDkY9vjqQMDEta9dNZV2Qo4idmqEejLWMWMC88yQMKATX67
qxD7St5Yp8NpcHVtGCvCz75E4pFGOGXRgOHZj6kk5KCU+IcUE3RHOyK3Bz5Zgwo4jzcvHmw/2s9U
wTmK9alzYRtfFrsgIS6x3m0EdbXdW3+I8L88cQ+JSRVI1JD9xpqMaaA/F2KRRg0pCrOc/izDjTz3
NJl4ubm9R42kd+tGtTFJBEEIPXc1yab4+CT7LwZpO76IQqCHYYdeUU8toZW+A7zU6A+zi921lJSU
XsmEBnNKv1HbhavTRCHqMiMeX07ncdm0ABfYmNnaT6GldMiwHu2Wi+kgn5eIMfVBrwFw089SqNLx
Kh6UIluK8nkCZO8O4KCx33TIy70tkF+904rAf/yPyg/E6dD24m6F44mDzN5veG2tgutrCjUsa/M9
N55b+6U5/oXqd3QzlEIB+gXEhRduUJfbGC4ddmlMK4ovjHDnqoaSV9Yv0x+UWl6hqP70jdAPX2xs
CQEY0Vk4b1SYkUOmIpGLCCcxywMW1fO2bsyH7luBnzSIlGsC+1z+9LPDXN07PY+sav4FOXHDfr5n
kP50Xz7fJ6cAJCT8+l6sGq3G2t+WIcXy38NPHHMh7OlWEtXJug==
`protect end_protected

