    parameter   LeafWidth = 32,         // in bits       // TODO is this just ORAML? A: Padded to power of 2
                PLBCapacity = 1024     // in bits
