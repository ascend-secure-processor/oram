

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NqcfqrCPxDxtqyqqf/QHxGnHhIUhihWFuY0kmWS9IPfBZdzXhtS9uZPGm+TxEbwpE8udxIw/bdzl
G1esVjxAgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R10MBYKxuoiYqsWoBycNwnxpi2/F3QzEnsu09toaVoJ3D857m+RmX3rDJkr3ew68p8BOLjXDxD9s
EShErHKWRNWRlb074lSKFmAVVCLYXErPI2MUPV1NDcnWHVtNL9/QrawjAKrVx9bn7++a6tkYcX4b
m14SmwGqm65B2+O+Wgk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0jdFYLy2Gpa8kRAt6/Uk3URZQ8d6THO4nWvvx2tS4yO2aUWFCUPcemPDP5ITevq27mscdxdHnZ1x
c+xMJCY5JZ8MAW/dkGlaiEghsnCQkR5dzJIrytoNC7YEi1RJgEQlB38eoAQtpNchwK9k5Ll93oSD
WO8niXDrt5/bqs2qWXvseUpF8G6kMYIyzEdI3VEVe2oF+UmRGB4tPqhpbGazBZi/JZuW5kA3sYt2
BGZh4+UZ5+plnVak7VQlDX4rBX0W+BtQhjZqyI2o/JjubxX5fhAz6VYOacwKTulzxUHmfCfXa/lD
KZJjFbFBLW3kHJKaf8Hay6+2j4jIx1+6E/j/3Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BC09+VWe39OHYM6AXzLVauRINp+xDuHHWG9XTFn4YdP/4pwWrMqMTjg4RZzOr1uWMt1lou184kh7
KSjQFzTzWzcbu0w/AJLXnsZOt90S+A0+htqNBXb1XaJAHcm6lUgLS/YzmpEQaN02uCH0H+QnDB1o
1L+KWQmmi8TEy2ZtXiE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QYtt6SX/XX1ZrSr9b1xC48SVo2QXqOh4Mr/sxLvUM+YipwT8kDJeSzSOAIYJqJMnhv57bocfB4lX
WXiNcXreudr0v1boAvr49k+rurzjOz+yijzrxWCfjEXExHboi6HKXcD6YsbM7IcpoE7uZafSO/fc
JBvSQKLmlSMAYvgdZ6ZjK+kVt1/KbK7r6kUzOGP4tliCxCUnPft4zCFbUITqjGIC9ubteMGuhQJZ
oAQJMxO87Lz7BTqaOhg20QI+T2MhFhf3T918+9jJ6Odu901Z+pd9rfy5P8C3ZoO7pNhMYb/gCj6z
y6m6UQDeae6SUu9JTuA3dynOYWXiyyI5zL9cvg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3632)
`protect data_block
JGGzKCTqy0e+GdsQZvSg4zZCr4D+eU8cpNiV/wdsyxSYjmlgBf2riTBqpjmYrFjxHZ/bKppXf/kw
NaCgFG72PLQYqXCupdu6/cmi6+SYTFjCh8VedXS/RYSr5oXh+igk/cfXu9C7zhQUTEeQadCGsu7H
UfS9WExScla3fJ98bLEadrTXZjgB0BJwsU6PjjCDD/rmSz3MiP+c8dbhxA/X3CoDHE1npeipBcsX
L43vKa1fvS+dzBgEzpBZM+oCuBjV9o3DnMHtsAM43Xzi67iHoV6HNFNmHvNFtZilyJjMQSXXPSTP
NtAk6dlymCBN3kMH2Tki21VwKJj+MSzwLzBkVqljZ6cYcvr4wexy7MoC51E2S62X9tDLGwVjmBa8
84TnX4GcnItvfOkIXO2PyIum6SV5wUapx0nU73QL+FMRkeCtFiJkc46HzxkixDHfJT//teJsUeis
ux7vZkwChVPXpPTWB+zGssd/CZNDwnvGmqXXaaSnN23Wfw0LSO94dAx1zxYPMEmmexFMFNs+tCh1
1BVZUAWggo7o0eqvLY+i86k60KEfkATwpLgBuw4a/euJqdbbR7iyN/kNmoveiHTx3hGHHo9e6j51
RqJmZOowidjaGKHfftGFqmXs75Q7uIvJfFnVCZ+0b/jRvF2Sz/YG/nn0PAoCqbt7uvwDjrXZjcux
Oy8SRKYcEnLsgBxP3Kg5contBn85NckGxauxtIAlNlWwbJno1bMCoCBSS54V9YSLWKTuYw+3kS6P
L99ntTnrD5/bprk9hKBHIpQk6T0BovsAqC3ZCuZLWlWy+w44W3gQ+TfA8xrfPjMFlOCL2v4a2RcC
ddTIWfAv6d+RjMYsE/S+zrAxdejCGQOj/Q4H2e5DIFqIwu2F8mirTtIjl9KZ0EMFg0XhdXJCEWbO
K8mtyp8Upjn90nYg7rbyI+hYeAYT7Et1/M2wxsM0V0C/3vqWflTCfwUjIgVh91CnRzWzzq/e5T2Q
iwNVvLeoCO1rpFluqkBMbNhTVG3fm+RQ3oyL9gSgy/UX35B2Dqj7CUU1KKxoqoY4I3lmJiiGFhuQ
G6MkXzTFXWqEVjy+50OOXOJqGLgitEas74xiwclt12VVQd8QeGm6Zo9xA2PUlJpTBfD7THEWF83P
rT8C1qZhVM982x8kEJcdesNehUfaOgVBo3K1tNZtKQz6ocZ97OsT5nydleqF6148W5D9tUw5jzhV
K1LVbLOdlR/0WH3IYNF5p3hA3i7PZ/CIuqP+De4M8MSk5vXeeY6u++e/rxqP1aHk7B7vZ+LNhGkL
9hbI/VkZRT9/DKeCu/bhNhdi+y4QZ/hgLeX0IxRvjFJ9n+bkeZ6OOULQDP99jQ6hZtaixmb2OH7p
b1t44NBC/CZepP6IkZmEKUaw6AdbKeCdkcXHHkpx2FHkTHixyRgGlxmN5mDCho0kRrPe2WQovxlm
rZdZfBBJsYBgxbEY+Zv9+Rv+kpeNiEcP6OW++OwE8xOqbEAEsqNLQgPdzXJxQXvnLYn5aMgqYVUZ
E/Urd5Ofvr8Sj+l4ypu8tb+VTdkeMfu3h8qSfsAJSXomnheUS3TtCr9Nyn2vpKLOOWH88ntaG0VI
0o+YNsuFHdnMxMkXu8el49ZEGwfyuKcDFxjUG6oHK5OfYwCRxPmtSMEY5p4+FcgQgn6ODwYWdceC
o/4jmDHvNJc+4vX9gIUI8NDGfAq31ddUfXL2T8Oegkqee/K7KX6FkbukIfjJ97Za1j3J5ax9Q8Lf
fIDgR9CMksrBumymZiTJCfobYQ+QYuIJOqvS9EaZOrR7DRhDeSr4x+WE7s3X8e/kdAPlqCYqW9sB
MOffB+sEQ3FAPEXd8qalszBkq1hCa6VcRr5aAbFxeijTwKsVENy3MpxEvDdGShLnzUbpksA2LvhU
wHTpHIuiFW0Xio9Qe9Tq32FteXTDn8xNJQroEh1NjFwkUhdEfn0M6TnkBx2m3iPp3cTRlPJhp1Nv
OfDNPpEpPfPLx002pQRrN054ZNXNbSbYWcbe8JenmHP9iQ8Wo2tPDWjfELXS+TAKgAJFRMs93War
kGAQehHZ4Y+Ujg7KPQsQx9AucAsQyG1FX3zvVhfva7TwP5cB5BmkfnBUM8A5LIxz5SrS7YR/SROx
K7vDPwS47HR/ZN1s2vzL1/bvhtWYGPkIakRKD7GAaZxdV3b7GU/uS+WjNrfo4UBlChBFgVNbELrO
s/JTUiupN/FMBn5w2PaSw62y7WaewxuCuz49cxyEnVt8aZBxAn+YjtflRIfkfkJul0IGnsCdVEvN
esJr4v/jV4ihxKVwPSU9iWUzCdhFjRfo2ZT1+srexH1nBN7cZrckS5A4eV+IlYVuwvHKR3lA4sTw
opgDeRoM1cB5R11TqywiGBvi70f6aqhNKLW5AIRpv7fF50+pWkWT96ntJUXmkJP9V8yq2tHzZTg8
PddZh1lw9eCZlhu1bR57gXYdZDd6LtlG1PF8gu4Yqyt+T93ZUdkulsK+NSPudpbYdhKFpqasfdQC
n+1gPlrGZR1kSQKPo3fLRGkFL8eg6+xnIrD5cDLRRk25AxxaTPXAxYhq6U7nHUykMTZoQZLFcDnw
djOGWjuIih0FMxhK/AxvIbX7MNei8isnaHA0ug+RPhA7fCA+Kgl3/YMZv8aL89HJnWVJ70ce7qCq
ZHJzdXE6H5RGfFd116ODHGPVOlD3NPG5WjtkKvFVr5fUYSmjk6Vt5cJkOJDc1ip53Mri1TvFu6oK
c95KTi7LvwhIOrXvsQJm5WxGfpJK3q3jCwpPhLoh9k6GNHQ78R0WYveDTWVUF+uT/lzBz2MBYwQe
TIdIT5cibrGNxiqlTazYFhV69nqQOoZcwBhDtngjtUpUPf1goDa5qMQbNdmfXWZe4KV5Dzf+Xr5P
DRelxC6jxXnGp7OTSoL28A1L6EkG/KYeXRzSrZ/OJUYxRW0uMOqjMmRcvZ41PJVQBeKwfgqsZm8H
0k9Cha/VVxkFguj6+zpfbd8x+BRY80Rlmr3d7aEzzWfgFmcUU8lvp1UWLHp1BrkKhXfFdOyR7m9s
KbUELeUXAvv5nVtE+/3gBzR8v/Ym+rWIeTvfc1O9Jt/4O5VG+x2y1BtQRfQ0YED9yOrGmAsmnx6u
kyuftmjbbYuYOgZpkYt3M8jwlITdx78PBaAwcMceQ9ZDaP4kakhgt5ZDWpFmmt31LzwdCBjUL2yj
orkoeYbtIuwmGlNRFE2KapfbyjpTT1eeGykis7sz2vJYF31o+f5ayHW6S+TMp3vGLuldIrcYIH8Z
D9pxf4y5flTlpev3fG73So4J4UnU5bbaIwxH0ottJpkoeEyV85bDgJuatzdhSDXWUbMQkWbPsPUo
VtRBm6jCyUzLStqihGQq4Zwiga2iCgZhbZ7oWGJ7bx8qjJt2f7WVZefj9mb1jcr15nIQOVpYqOS0
EC5wH7uwMeM9V+5r/ik78vOTMZFzzj+ygj42Wh0T3aXyG1PPPGsh+mDBE/sFqVMmUF73cK2lNlm0
vpCAj9GUuMPgFaxn13GJLvYZoGpyPAWQzabvotgPxF3h7gH+7RI5TUZmF5yZhDHT/O4Jps744kfk
fnpYdA/sqzIymTQeasquvUHCbjvXTCOfnHSm6w5pBry1RLiYIyrxm1XaEQTnYKNWvYkjGdWqkIZE
xprSF91Y97yvYSdvnEgAZax8n0AYbs5js1CXogf4FkfBZXbyrfBTVmF9Wrj9S6SthDAy0M/8D2Ti
Mw23G6U6jXBSvvRLdrPbAon5V8uNwI1kvCGe1fcVefwSKy1Ye92J/C3wXUoQfL5lVSethD+AVz/W
7Pw3+clvs533m6Lwj1rprNmDhMhki5yYu/nqR0Gvl2/7PmO0BGY+6NlKaoY0hAYW4nG8cUBWd6/P
LEk9MUg8BMFfJGWMCwt2zH6F5nKVyc3a3kVnmft1+3MrYnGFf5lEQ67fY6OoNTOFmc1q7+OyZP12
uI4nWfe/Z4cGUD9nR0rZ6Udqqc5qzEWDJTXQrMXgB067Hr6kFHrB7sWlPYrCqGp+6YQfbjNHP4F+
LI/Ja9SfbZ9Vz/m8I5FLSvvUu3Aqa1VPuIMd1YPY+LLm5lhH1PDfoxHkxiDLrRBrpGOxFwxnrfGz
2sYXqBnuJQopYBduizfnFY46pq/Z3HQ4nfRP2KLXls9zTY2XVIRnRyu9lXipsodvES/B+AGsI8qq
DR7MIKQHc1dS0lJmZNTGVTYUMNs2H5o+E02YtF22E3Bw+xMzj9iL8TZOQlK21UgpOBsVamKFBscB
xkSeH5gLi2FjT/PNPzd3TLE7Y+6fh6yBcRcK7xkoIAVMrYI6pFcOdeIB0NS0oFSjguhobwcGYwMg
pzQX6w/3Xh639eEVj90F9lhhR7FHzEFDNx9PlK71dXbRtBXr2KfsM2nchQqIjbZK0iNI6HgQK0GA
J+/OPs8pPv2DF2/JrJhHYlCShjDCzYuPs1vy6rz0uPi7Fu+3TXzIhX53VC2T6hrx0lGlc7QHIgQI
gfjiJBvQmImgIPruaeXT6nngaWuvOEfcPfBWXgM4MfqGb7UnTgM7j7IcxWsxlmEOHzLTr+Xls/qi
er1qrd0zAi1HIpSYZojbPDsnFqElGGc+y0pCIQMb/1Q3LWELOzo8NzW5jGpR6NIu2BIo1BvYAoa5
Q0yh16Oxbmcie4He1p+EkReIzAHcshXT0MCl8mxuYdvsnLg/fB5g1SRtg16xUTgTusmUm4E3TCOr
wTHrcfxC7WhBJH2aEc6SP/B1gWWdSIWbxDvLonXDIYcDFdAHUNZwziNGPt9U1LD2/+z51d98kpi9
31mrER8Sn/nzAv2zpmB2ea9kd30+sC1YUxZkAgJKYyc4ctxt/6iNdO0=
`protect end_protected

