

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MhHHu/EwrU6V1lFw9QOiyIulzumAAzXIhBEyPusapwCVDrVVOPo1pCJqx7P8oZW4O+/9kKanbF7o
pu86MhqXxg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j810kuRYS2eKWBbLN47fZFXdxIM19y2PUGjMq2wzKbYb7CapIwrWDWR+iDuU6oiT1U+ELD9i3W01
JtcmM32IYDIU6IyZgVzSr28yKufPZngx4thn2cePJARB5Bj/C6sm73DclsHgqJoL5FcfnpPqhgiL
bKn3Gxa4Bw2CMfVGYXk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xL3TKtD3A5K8c95YU6m7lojPbkMQQAfSOzzkWsPu09jxl6J1Koc6TMu8QY6+zWCm4ZLoPq2c3dVF
v0OpuzOhshUr9LvpvqSTwBWqEbL3lnkPHXgU77mQr1uGbQAhdJC2CRXbV6gbaEB5RfZa22fXJhK5
qOpAp2/v9d+FHIxEI9OldFekV4D1DEJ+I29aLFQrybivNmun5VjnGW2IJfV44v6WqqliMg/yWfck
ioFoJlGPSiLTNUpMwQZIPW2X6xjsxT4Inpfdv/QQHMG8KnsAsMpY24bIGbDNuZhzv/Dxv/QGmBV/
SkOlU2YllWxMVulnGrfltdJm1CwTYGvvnHpzdA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UfemKMsL6yhRONjbIIgpWfUKOUQyJxe1FC4jxHkffUTEwSdyTzwMtudNsb9dU4N10IX2FdHZrMFK
MG1AUarO3PM9+F/NE78E+a5TIIe48pTBhhY141u0QRGkTJ2VEGhTToqJNi15z/ATq+VA8RpLMFGO
MDIJ9X+C7WqtMTh+/dg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M6NevUSft05kaB6hd6t4wiJslySTu5tKPW783+U8fNluG0fgWtTAAtA97WCk3Y6ZGl0UpojzPieN
1YEMhEe2I/Vwtv3k784i19VJccv6ALKJvjXDc1XxoCLELmLpLA9SUNn+qViQsrLMxUo1wee8OGmi
yNEWJEar6ZkpCYRpWqiU53OJ9SSo/LKmYq8lgyGOjvhqIlPhVYnzC+hRqIxZNAu8b9V+LKYY/PQM
P3NruyV+Nh154nETQjuOGymsT6WSTfOSR0bni0DnLU8wGKzBGZoWb9TGCfEJ2aWSgplUeyMAww7Y
CAxGDCQWvSvMizOcpCx77I/+BgwU8dhB3Ovhuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4192)
`protect data_block
L/PoFUIrbWMWn05ha9PdcJ8Ec+WdxCK19X9xlANx7vv+2c6xNMztxukOZKMoNikBFUzS29QgWz0W
/NZyOdkaiVrHeD4uqIi14ST0EbdVyHtP39uS92F/QAKYFJX+wQW2KJo8/IOLVXXqNwWBZHHyXGrR
s2ZeqEBKmoBCzlpN3I0C5uUNtwo8wXGD1wTS7jqTcvgFwZKwAWHBQtwCHe77qMXqguUp2+2GpE6J
fCiquVK3er6kdC767H46AYmhXrSAYlZwvhmLo11tw7RX8f+KVqESGiX1cviqhe1j5vHUzvWMCURa
LhfHuOkZQ9LWpcOOuhZGDJhZAyJuJs4tLou7JTeA67ObON+MOFosV58GrrQ+8ppEHFkfRuoNJHN0
UBfa6Jsk/sDPL7ZY4j0q/E8NObbHfUccn8dSBrLmnODmjWzr0vJ4uYa0yavSNrbEPh/1CjaFf92y
3Q4fYJ2QB2xt8R7dDGUsa8LK99PgUg6wogIZnuENdjGSxmyps4dghNntrLf0VHrEuJ7TI2LG+oci
cY6Hge/BsYmT2mUMMBEB4xVMzsjoeN2ensSF78TuYuvWSHihkqcFXsQPphQVAeKOXAH8r0UiXD6G
3SDKeakkLll9ImFmAYGRI7OxCJa32k+/sH35XS/zgN5ot5fOWlChZ0tM9iFXu4fjK9ugIM/V05vu
GXdRbyPX5HV+qU/b2bhO1p8IKLF/CK0fVtKNBaHbkM2JcNMkGJ3zxGsjjHUELTTKw7QP0p0WDke6
YCxyp3OUnkZpzj3Qf5KgGFD1mLNFvdX56Ph2Sa53chFvwgrTXwBJTjKX0IH0o6pbtomvPDW5qnvY
fYnRnLKF/ZeEZ/0/GsBshoVXyYDpD0p+BOqfzndsVg2WD3AFO+Y0E5CRqFhMH356fOq0E/BWorqs
CO882We/li6IsyzRrPVhOSoO+6g2Jczpqz7nchGJB4N5dIuVQIOLvYBmMQmWqgwN/up/XJkItYIN
UwRp9VrnM9yuzeGaHMerkBt3DXaPJ5FnCQ+yKaUVIV90xZT9wUB+DFXR3HkMS4fJCOwzUIk/nQiV
hXlIIAFQ/eEyfoMqe4RBWBrX2ma6syEdLGPIpmvCJb1FhgfDbvKSr2x9TVHID7AJHuEIg84u0Jeh
qsSggmlgr57WY+O+StEj3FptUcTx065O4U+dktpoWgnUvKdB3DFA8Sod6TbDkTFQ9RMKoMbJqdXw
QvzEsR0JG5pQQ/5Cv2Z82LrYgQDM7wfgnolybvMKFEVBzl/KgmbmTFWKJP+4KMiHEGI7VXWO9egY
vCAFjYJfWXRNsNRsXN1TbyRRU0pCsU9RGHLwSBNFt3vhrBS+cHIz0Xljv1ujNvCzV1TGHC8TY11P
dUO755CWsDJ7Z//mKs4XZBIELkUBLaQ/7eHG9vZYTjraOBe7kNv9Tz0L5ZYwddrcA4RP59Z+3jvM
122uac14BMHDUO92hhoAhvptegK0nDoyA2UpRBMQvn2mggMOzEd8zb44UqpmsweG5fHOInFKWy9J
KF9jxnmNRdTOZPp5rcjj3eU1m9ThRY2pphsXqCVYxoZTxKFuFWv3iogGRWJU+auGAHDEBQBVCjKe
3Jjbjr4Gi3GINtCIx1KA7f5zeAT98FosXxUnoR2/KQc+PRbuFaeYF0nRAvjqMcGhfUUmyS3f7upd
llqF3GkB/QDLyDMQ+PwPhck2VbI8Hpv+JgRyy2fiSO6oH5flNmyR7hQxlf9EqNsg/f8+KZyGzHdC
5T2f2vmx28T9GHIs1GgUJXGVSN3sOFgXRYcxOiqwL8xsgRUbTvP7P39ag5aG8M7JDYRLpz8+opqQ
sxgbXC2t70EO1NBFqPLcGbTckjounom9uLrQ0TAzhnXrbJUOzsidgKRJYaX1P4YutcYHsh9EsItt
VihP7KIpfvkmn7+N72BCDycOPJQDQvnu8j+FNmreFQsLO0Rx1xvPBJ0TzCHDWh2Vy5GSm1fBi51T
ExqxObd4BkZnBXjEKVvzZbDsZ2EovEIcujGCah2xmJyCRkTrI8KsndKVjkDuoMkAmb6Q1/SzDvwd
oirRq0vmUm2VpS43Zcm/i3Can9GSDTTZBn81FTwP8RPhxZKq4NVocwuZvpmDWbkZ67J+Yqzj34sY
d2sxn58dPWN7ID+MGTttXLtu97xZhD/oE75hQIisXtci8f4gyqNdpxiov0HmIsYTDSGDJuGin8aI
mSgizg1VPkPIh7v8WYnsezJrVc+Umh8JjNrOz8EfYJlefJz3DVGIA+p94dtN5T3CAS5/FclSjr4Y
Him60hlnku4pv4pTqSnQpNB7I2q9j+n9npA3PWvOzBciOAUL8FxhK4htgvQzS5VoCvW+JoR6HYxO
pblXyuPRMibJRC2BindT5Izn839TJDybN8OHZ5qLfrHQC2W4+eaU8IynStBzzg75KUfw1kp81eSp
g95w4GF7vcVy9M60ukgnzXvyj3VPgDM+8/FzskPdodSj6ZeX1QyygbKAfTk8hiFwegB+1ApXoDth
k1UGjh5ytKtgFJUkTug/AQKHqNnSBBq3FnY+yN+zSLbyXpkNk06f1bqyo1xj/dqvaGSP0xnUCToM
ERbuJ7+QHXe2KhcTa7IR21sxtdBPgejeij+lUssdAR9A08rwOUnfTCxVWL+8ZBHixIwW8su70s4n
dfxUP7o/d9N0EfCqGgGGqa3h3c+kEUGchnWA6bGrTsPI7JD3Ly2mws91TgsX++ojUrc7PvK6aW8i
BpHZmsty5Fe5BF68Gs1Nw6RV4FaTKUCsO6VR042RoZdjW5dR5aqn92htnKz3dgqSKtnLglsHXifb
fzAuuaXgpDHs5jTgAm8qMj8nJii5xqC5OhRihg87VsqqZhkdfuPoXDahYUasdvWbH+QBw80PWkzK
It14spc+DG/JNaGK+aFY+X4adXyuQ4zpeSvHb1IF9yc7u3Tjd0Dg9Qqd5NndKDx9HbZhdRZQ/AOg
4X+V6XXfIvfKq2rIzHjJg1XYQxKTP8swBSLp0DWZeh5uPy5PhC9ks7SRjaQe1/fZXYm/vvb9kYmF
jWIw+rk3DbfQrTYti6CD7nrGr5jKtIf0kuJ//LvK9md6ZP1LtB+C0vs+MnbzMp2lqDhWUAYzuYWu
TOrRszkp0BCovgj+0I3ZfMEYK0Gr3k/Ty1Xa8X6ZC/qlTDWbOMcG072j+PHJv9TVcgHp9lq1iUX2
xwjPCmbnYZYhhpO0v2t5POa6VJRo4XUlOoh9tV81xpfwAryuaXKWAGY9V0OKupx4otuubjtJ2LH5
oz6c6ofGPayFm27wTjLUVJXaGcMZU2I8BTvysYLPXqP+On2SS5NNLzo6DivcHx40ZKvj7IbAxwHS
lVYmJvHKP5OUDvxsPrkGjQMsDy5KEaTA1WozRK8cjlwSZo1AAc/5WlIvd+hHXk5PkdMXvgs8XWHk
qkmTsWpAibdiN3MzhHfChtuP6fZbftaRJ3QaR/GlwBgBiVziyKRi5Lwab7vF3WsYLsgrZPSVieJc
mvxdA2+BtW+Pyg9N+rHhTH/O4W+iMX0tY2X6F1E8e4F98zitxBESjRO+uS+9+2uBU8AstSpxLIjX
c/Pkcy9CeBGAk+o8CIxLi5y8SAPftLNjEUTnuDMhiyB5JNGEdoxPGFpL78liwtw9TQI8p13o8FSt
pqnRSgUPx6KKIuyyHYY+iIpCUFBl1N9bvNKAtPpI/e2H4jzJGassc8gf4Ef9iqYMUCM/D/r/cNFh
/W8MteKYYhB1j8mkc5tUhHcR9gYG8kJF8TVYWeTIYfxVQspHNg3G6ExBXQG6ko6Ahh4RD7a87V92
tr7VRkcAQNcvW9lqoKW6qTY6D0CrjiGsHHWmH8rl2eywS0ftbkiqZTU/gKouLkNllaWwGFtjEAeh
e2RjN/m9TXbPddZDUzRYepCCnsK+yu49afxICIoDi5fMLAkm72PDjofaWxgQvf27qCQ5gZkJIAl5
dCYwIgUF1aEyq4K9nPaNL7pqyuxKpzyfL6beOSpnEE0jXTHHP2Ts93DibrJjKnvouxv49OR9Ymd9
wGIUeYi49MyquCxbpc2W6/f9iT45z7yTtVfEQW2gPoThd0SMuEqVC4vp9j2jx6GmbkHlDolw/ptw
qq5DB7FtGvgbGdRZq4dWGbOI9XBufwRj7Vt0p170okcrft4vAaOkxo75JIuWODciPp6y7aZNhmXr
hVxTw0Pf+eEaT1nOCS3pHF44hJ85NYXghJvRskCDVQNnNw3IgUDo+otOCYiihqtYabiDwAaIwk4p
RuoIDIdbOUkJIJnwTTGKHqMTyrvlDsjpVPnT9ICCDraoiNkDxFiyjruOzpHznVbsj4gDphG44cfU
LCVtySlAjV4braHY4uwaPzf3AOMnSuRi1rLM55QG/Mf2alNwO9Si/VtGKmK+/S0gHqGSnHicGcmX
CA7mamBsUprsiaEf14/Cd2v2scneql2pWmZ+kkViuizdFeIZBegSdro0oGbUdWBDrqU1WzZ5OHGT
Iwy2HNasVRUAUKwY/06DnwIM/fXo3iLODMEnOdIl4w8EaB4Hy+ii03ufVSOQBCtw+yagtQ5cSjFp
9thvyPFBCv+X5E3gM/aNE1Nbh6+08MmYFvg6YsKdvV6UUc0agRAqGirtQ4eeMrBQZ7bpr1Z6PZip
YFMpdHNLEMgnq8GaI62YEvXpz7U4v+LAvhvqtkZoC2TN/oWgN5si6bHO0ruVFbXPpiJBz3lP8tqQ
6UroELc/hX0Fl7VOB+RenJSnA1CKQQKSr26gEhmiJc1P51FD+qyI26+rSPJBAt8USnd3Q32BlNaf
2KCtAVeEWgAErx9Ai78RLODqrDc9Zpi7EPFiR1XZJLlrEFRsNpGHc3E/OXM2b50/R7GDDouiu7wc
PehkRVMfaKUPtpZwkSighnVHfKny+doALbbl97haOjFUuV9cAhMwt3otWHzrwRfGHCkZB7iOHaqY
UzMLHpFQ6gn5rZVuXjyEkW1yj3ng8kCNkI+c2esMhpMmYDnl44bCbFZO6UzKJMp6/tjPvAhHw5uK
k/lmPGvJGgoubRaSC6Tq61YpZmpfOZZR2+7UKHnqCskSMEHljAhRwXFGRek9zMsa5rghmUNWROIc
zyqktv8Se5Nn6/emlXjTDRiTRTfbeWpcXPolUUk+3pYP5gRg2N5q8Uz3Oyh2OLgVuh7nAT87PXNm
cWYSQ5DXv9/F256bLLj5OA7+gKWHfOm4B8xY+j2y9e5ZO8BCaBir3dX2Nbpx3PQhrNHPM0ycTxbT
u7R02QA3Pv4t0nG7qibNUsNROwPTMvH+w1WtD602kfqqaHj6uBuPg9K87eevKFqfFB5Bqjp/DKGn
+qfd91gjgzCrAuhS7pegyPAdauXJMKkMdjHnKHSvvDhBnwpRShN0cWMosYlDEcDEYiY7imWVKP0H
2N5BSJgjbEMfqSbvDg1I4LN6NGoQB/a8uILBSy+DEueZO6poOmN/pG/XU1Bql3eBjuSa7+Gc3zjQ
QIGCNVdgbngAGtC9jZguQfUE+QR8Zy4RD7jbHAY9x2CR8l4OPFuiIkImlxVfujCcVXYlN4qn+5m3
4KHLnLgnzb2eNjSaMBcwBvJ9hSjdP2feQtMtoWqTwg==
`protect end_protected

