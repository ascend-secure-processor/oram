

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KfLthwf0WHQIA80szzjpIUtLyag/hGKx/V/H10zUrT8gkNcHF8KdUjbIk0G1sK1O94j4FUbNpuz5
XDDU/iNbBQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pTSqL62MyELv3rBj9WrWvWnFClNqkkzlckYP9f/g8B7vFC/32jbFMM1dxZp4gUu9an7LDO2m8aYK
sVYBwc/bGLZtn892gQ+LTWrWq6EzKh9cfrcEwaidFuj6Po/X9vX88bbpD9n2DlWQ0HV46xZp1N5H
Kcc2mMyHTRivjXwnyfk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tailcOcBlzLWArRLM93ZbvLSkJZieQOFSfrYmr5bL6+4uI9nZ9ZXJcdxGh6T829I4EBjNN10SSWZ
K7lPEJ+xNq1EUbGQPVSAi6WqRAd7N2/uFJHP70zY4CNwsauQ1Dd/9ivD3HIyVu6NMuygBS+5qbF1
PShy+sVtuLjI2duGftB3tTk0Fa98frloziZ5XNbDLNZwXrKgmFSG1yUaB8/Cit0cV3lGDjbpA2Y1
C2TfDg7hsKhJ7lTnOWm2jEJrg4WpJvt7Ybg5re8J2C/Rzqzha3JbxJEbPFJW+vVsmnCr75gDhp5i
dLwpof2oYW68+QqgZl9AZcibfpqdtC60d+9pgA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PG+nJv0T2NotLfYOlGEOwRu4Xv3Pr4pLmn5+8T70+nsaOZmCiIPoKe4vEXcZ4iCpVobnTg2neeLl
LEScFQSU53OkPqaAngv06Sux6O+X92HjxqVSYNypouJiVRIGQYgARRnonjrLUH1zCMMRgLRxw5vY
kPXcQCf5HZDtDK84xAI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNsB0d9SJpI6ALOqxLCVJQUftaNbAWn4lgHUYFdyl3RCrNmLmrxSsKeEonRjWp9wdCL4XhTQHsr2
ndGA2oIsN1U8hfgncqyUpbCf6trTIE9TdqYaEZJWKh5d5m8m5/WDegHKhyacw5GTarf1eT9RNQY2
Fh3g1D0P5p8Oi1+MMj4BgslrwZeXyNXcGo14+ZL2ZOlIjVrzfbFBW2U7M4QlEA17SdGQFd66PWqG
ERyb3FnjSpiEXuFfWffZR5wiUlGnXlTRSs+Y95Pp8/ccSn1ZeXVDN+OXQFGeLVcZXVzQMlzxYL9V
B87vBucDsoMM0qwwu0xN7zNV+OpMazFPeHShrQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9904)
`protect data_block
4j582Twxii7Kr+Qj1A+0J6b2w4J5kaMZEKYthazxTZ7GjGKKOMYZYhbwC30244utGbmjZ9H3AAMX
L6KJkGzAaTL7p2ZCPh1a6f/VfRvx7CAessOQGuxAqScVm7QPOxjAhll++G3dsrRTKRIbSKsV05cZ
eM+rfsEJSQwJNS85GFIUU8XEMKk54Tj0/Qob8Z6p4FJ9vW0G+YP+vnTF6Rs51GyOa0INgT/jVZJo
ZO5zn5a9RA16AYNK/MvfiugVCEtgOxC9CmaXMTSunTVeG9nRUU65QgV9gBvTpLFxwnZRD3thCG20
W4Jqv+xxEHQs48y83vubmPqwU13XlUGwiNzGNmpyQF0xW37v+UyI0MbsaKZsk50CmO6sTqoMpUP8
58RnJ+Pt0L+ji/IctIfeI05H+f3xgZTE+WVSU2gytMKuP+f/8gWIJUXLp0ifHddnAkKO31g3gDs2
U3zGv9dr72Zt3RV1FMDMKZ4PHoFfYzRqqT3bkS4C41FDV4/vmeP4g0V7d35X4fRFfa2FzvJoWmr8
kfd8ph3GTT7sJqVYzmD9222JbIxiKhKE21LuVT/DjBnvKYjUNKulvAHW8/3FFzMTcriRayrgPfPc
tzwuG1nIEsCBrSobesJ8MOiclNIzmZcT2+vR1b/VUrDseMoIdS6js4SYHk9kPP59caCPiiwVrKMb
SRyDZjVVbvgQ2KgCUDqzDmmf2Esukz8GVVbovFEW70PWsqbESUQQTc48MHUu6LMN/qiYBQG6cPHl
z0LHRTDMjQJ28iIsuOXSaRtJSQaO9gUf75JBUOI0ZncrUWO28kLF/sjWwR6DW+bZSYU2FMZGw4fk
kL/vGJuh6xofRCLxXDnbTcdPwgEppkIUa+XvQ0vcA9yrFKKzVPXAoHiyCFCjU46bz0IMmQuOk7cy
GBXanC+MyDQGsLIqYSUORg+uGjKLF+CwhP4yEQ1sr/UgwFS3M4r99mOy7bKvbJ5Y8aH/4BTLeppe
qVm0Xb3buwkbwzgzZYNtcVIp1f0rPvci3JOSnBa+Ou9+tJsz5C+SRDowTCSDWKZaxikaa+lHbFOC
lnlgIY3NBtCIgcDHLknDMS+TBY/lUue44Ut+Nj3CSdkHSRcl6Z4OdWmTY+tVKPgQQ9mUdNj5iU2S
csiOXaoWSnpSRC0rc+JmIxI+ugltL1e4Rr5XLQHborp1WwGGEqw30pOCkjn1zG6HmEh/7lUYknfx
xswG7hLPLvgWuZP/VaLxvwvzotmkazA2msK/jt+bSn5JT4DnVURoKefV4L3h4lFgywqDB0EDUlw1
+tZ1xN1yVWleg1pHvk47YEYatpV1C5BHhqmxbAPmj6WdgM8SDB0I+SKRyhswbKoX7BOOsvZa4TCA
vFpXh65VezGZ1kujrF8UT3wBegMIjUNPOeEO3AL2Yjzl4KgUD81hi0DjCuApxt/rgnRdMQ6oOxxP
VtIYvJXziBro3srjBC8eZv7oSP+GtO+1tcJPP9hBqbBuv27MreMHFpjiuJhjawF3VUg1vQ7YINox
WYoA+paEQ2UnBTjW9QA/LC7qYLVIwDE7H9tAezZIx8OHivd/FySRr7xSde60JSewv2OWOpbwRmrS
BhwgX2xNVY6p2DRcKwS3076v1y/p8t9WkkOkQ3vn2IkSHVUaDkaE6+PhkUEQcNqDTvjdJAUpDUJU
emmLNjjSd+TSAHakpt5IIntSMKyjp3Pbvb1odVN/gL+f21M7FfLTbTLsiz9IaT52yjWP/RTTDeg/
iRi3sl2h5qJpPhTzzfP2Uf9cbBJ8ZtG3xo/1TUxCJvogNKpkcHITi/8ZDJh3rfXRAvcl/owk5hOL
RF1EhWnrdxW8K3XGseJQBv38LOsrzNUSiAEXCledq1EmcVT6vpztJYfEEtqv8Q03JWxNNw90cGLx
tA9BuXuLFWWyL71zj1X0oNXItGrwRCQuYw1mYq+X8TZYeDtRjG0p/yHxW0+2V4xwpmrV4kxDfwN4
qn9m1fzl6II7pV0TBYkD9yDCGPq21rsvpQ2ro19DU+ysXBqjm6uiLrDed5gACWEGiza1vAd1Er7m
htuDoLECj8I92rXNVqa++Kum3nTdBJKb3VHYs33TXj7DflXSqu3OYoCbveXeCZUXyyNs55LfsFOA
Dr/65ehGyWHteL51P2uX7A0If7BPW+TbbdwIG1sQaaORMjhrVCalryX0UHuswD+u4CrSMaulFiHe
52wpFZ+NBvDS1vCZwyXmcsG5VjkDq4M4cW2SxJHbFaEhpMlEicOMhZdRut0L/bi5Wvf/2N9TdYn1
EzMoyx5bFSazxXFu4q7z6ZM+s9ygngE1wywT6Rp2MyLz+ZImJeKF275MP4SUosYmh8aJ+YWd+rtX
cMDGH9iGrnhS1uB0TVxNGEIueK42ptugyaIIF8cK6B/G6IboaLF42rPO0D2lUiQovag5bT/+Ws7B
Fe3ldpl/NsJWGfu6W393oNK1A3zBtCoWl/oDY9XhHhtyNbwILDXHYShZqv2n1lvRnRaUei4AIhgA
bnTOyWRkQJvFONJN0AH6IemK8R1U4k+svKNF65XOkaXL43t0RVaHBbNuI5jraaf5qa1lHRMyHlUd
ZIoHov386yqlsz4w1Latl8Bq5R7ditlQdDomO2skKlcv0Ifah1Yy7O00jUOlT4pZKfjL+2ceCMJF
p9Y3cUa5xMPKRv5WakgxoYRpYiFax3DTEF/NDv2wU8AKwiMbsa3LttTWL0W24hB/y0+4pHLP6HG1
pGEH/48MBiLykdTjBI0+lpdtrHvvFVdPHe+ruoMJzNZGByRFyOXc+UfRfjyP1xiLhZ/Ek4RyqJ7c
jeegUWX/JJcwuh4g/9uE3IVoC0IKcphSLiWJ2UV10JbQ8EI6jDUfoJ7oLz6sEwdekqqzIwv2/LQn
jUVYFs8T+ItC5oADfN6P7WPBP2AKTF2I5ZUaFjrLJG/Cj+TTfmzXD2PNRg1SzxHvsw0zskjrGYwO
wGZjAFVFroOr/yMF3NUQQ3eQQtZ00MkbfPcVArMw7qJrpzV5Y5kIyG3HtzEMWwjPDR1Ksa1+Y7CG
lI7zdGVX1uVJoys8PvxdKfB8RkmoxeZNNUM3UbVXFyJvT1pzkb+FxHgHmf7XJyGuLOrph/XeUOfm
nLAnXM5IHtpVbQa3xrXicwAR/snqkjTIm1wu/tha6ul7trnG5hQkxGpBZg+2EAT1hroth3qccHyb
uZaDIc61AxSL+u3TdwgUafDCiM/sfjeV3ATQV63l0rh3+pSppBI7EgRr2oESrFcTWtqrvEclze4A
H/XBwLtZ/bWbJ4G6gfpOadrXxpt6Uiuztp0eER5iWiaTc3uNiiGWs9zRagQEH7UAX+yG6lPoHIrj
gvqJ2GGQSzYLvEB1G/+IG3Be+rsX533iETDlu8ckbnMvFV6cdpC6m6TJ3PoP/7S3aoXSmcUApsMK
RayGOLloW1Jw/sBMxoDwsVwX7dZXSTGQdS/3qkKmpy58wllXuxDgHQo2f8yUgY7+t0OBw3pn23Be
6jFeQBxCGjbRXrzf9HsX+cii3jjpgYJ1bPxmK6T4LH83emQ/apjtK0AE3kZdfe6jRYjDP6ixaXPf
vf75AA1uHNhedlhtb3049ZDFSdXOwFbgwoeZFOHT0aI/ybkLQQ3lntUsdU5x44GqRhHhUI3MMmi7
/lqD4/A4a40wzAoTxhJ/knLdExeFGH+mvTKa7P+sXJWkyZnTE/6r/CnkqnRdTauo3ypBalW9EuIX
XfcvEugjLucvd1xLipbel6EY7zymvu1A8BgBtALg25V25WZjw94J1zRnNRjGizTG5z/LWwc9/zZX
ITcJIlVhc89WFS7bvC2eo2JXS9MmYidMjrNbvQbNmH3IZepc0ZNksdl5w/ydIoeIVzBxRgU4bFg5
dsMJ1XtUGU60UP64nLR6Eq/OXTvDnFviPo8hqnv7g+/hP8J7Gk14obKzMNaFNbkD5Z6u36Ys/aFu
i06PXsMG4Bx6KyALVl1yTXrqa+P+bBdyx5reboGD3eiyK3EWU8d8TTBQ5VBhsdly8j+4EAQn7Xs9
umz7GB5V5SgL+p+hPWV3x55LsL4/bVFPuMUXOByIfVyXMVMZV45yyZHZLiJgcZ+DLh4HX3RFta6a
ENYPw8bUZjKCYnrLpErfn+GRh85Z+0pUzHvh1BjCWIYSbBqxHMb5PDAgw66pIT5INEjLau32ghh3
xooV72jKj7nKXHYQIgRbIbcV+XNZzukfSkjSTOrbRcDLtaCON0/pG0fqaUYXHoJUXfIAnciMeP9U
z7LQmM1RN7l/dMb/jPNWGnWr/nvFRnNZ4oif2I5gyv0Sqqs9Q3VAd8/gplk4c6LBtN+Wn1ltt0/Y
fVfTXIDCZv2VgQo18xQX5YD++7v+5qx6irFK9cxcI6yuj2Y0Q0e/TRM05seUwgQDBAXEWw4DdCpr
eVoXzf1HzUxG2l1y7uPOKmrEW0WCGn0CJykef5UOv1Dkv/EyPE5Y2sAGvVYigEisULeBtXhdqrC/
1EQKUWc2u5vNTp3DxAkKPecgwNxffH6tH+5MVC0LCYSTjEsgPesi1WPQkfKows9cU6XMfoyOAsxa
1pCJ7Nv8toOl7UHU/O9IHCdJnE+htwNaVUYC7vnnk5glmvLOsuYvXwHZ6uyB/lEGnba/ooTqqOd5
4Au9aY5hSrQysFJATpylrWbeecmA8a5K7i+669GTrri3nVjxGmAB/4gjm2P2BLg9FToq8ZzXFXez
ag9QtO4KAtPtQZgFBI271v4SFh50CX+7AdL5Qdg/YcFq64otV4byE+AMZb2dpx/LpbHBMSqjsABs
sjSKfGDhAFukB8x+hlqdhUCu3YqGcbe8BxMw5WCEAoXrjNam37ehp0Had1TH2m3iF0zKDTdatilH
vJ1hESJD/Ybpd263tISfXEFtdC7sN1jy5pmPN/m1iHZVZ42jgQvJIOLZCSQQJ0ci2HDt4KCVZYNE
mPvpAYaizgL0PsAQ3Ac8W/gk59VvZlJ7eIskmYPvOVWXhMEZDIiNAB0KWKA65d4LOt0KG6JyRw4H
F3LwCjbQf0nChobHe4eTG3DL70NRgJqpB9dwAFZ0aQsSgEze4h+6rjw4Z7KlQDHOyRfhJN0KfhNU
dLKuTvwZcBWNMk7OHswOYKmel+denPdKwqeWoC+q2UQQBiLRl5KgPpWdfmxO63a58vTfEF00MXUs
aOU3L0xg1j11RyT9VUDD1Z8Hg6Y/oTYg8NYZWG+Ekj1D8w+munb1WQFScqB4CdiNvshVUcHzKO8/
snjaHCj7B0ZKIdnJxNzvAjfQENSsaleXPJFCn+fmqLVB3eE7j5MEoeoprAmL9GsiGIarbmvERVzM
4UpHNR3PdLTarcayARXZgoHtle2CSlkTTw0b7FP5LfxAZBpOZY2zoNNPcfNUhozUOUQvOhLM82y1
21/gsMzwUhY9CryrN9+Znftem2C+kZulUZMc2ChP1CpnjW4UrPtdDpaePO7D3otyIHRcdtNLC+Tu
j1/kvZL5hh0qEIuxmzRCHwZ5893uV4NRuu+QQDu+rwb/LTkUPhHvdO3vSc6ugQUVfMbXXCZC82xp
Xfg4Zzx53Hg0xF3BTojJyKFgSvkIqIYjv+t4nptg1kHcrmalTDyUwfoWSj6uKm7dhXQlP3MkvcB8
Cfr5FODznODc+aSwJrDYG7ZR/bgIB6caBuRIK2e9MvBPgFtilxMvY3hYqfKx2y5Nf0a2iLeW5Gx/
Y08yNMl0hsV+QhdtaXVpwlS6jfG/CBaL0ebhvq4+EI+HtgxmNCv72bzIyNOHmJA4NeRCCLUWN9KE
+T/d9DkEZD7jm9UvbGo5357pwl+6V2nrebhGUDlmGFbpe7cbupxetDJIaWq2gvWPuPsWU4fV9DRO
+s2D6tKghFZpASbZl4lwbKI0L4/FbsHe7wqe+YNFJWb6sXhtZRHsE8vSOiWUIA5R/CFah43wnCiB
MDZeXfjNGYM3PaiYJ5TJr4/IBc1p92UJlpXtJNopqUXWhY/mijahIxxxvdCeYg8cRQZlznrawVuI
vw5eqYAVheLgRua529qxQhLhIAnedvygEqGmEc21sFlhH4zWO/xNezm9gs7SKJlO4f2sYzLQoVK4
vmHtcERWyP/CVq+pxBPm1CUOLuR7UHsphKccP7WqYYTo6kBEvnfD98jVLYZqcBtYEUdj8hWHNv6G
bRDsELenbsq7/bacOtoiLVHqIPmf64ifAcOZLIM/xYfHXPYuK1t2axy01G6F4VreRgUTKqELZfKY
R2dPL1t7M7FKTKKuI7Zd1uuAbGR4HA5efxXLR7+uamcFfI7QOcGEIuFEqbCMEvy8eY1nQIqkyLlc
AjmovJ1w5UIfEWam57zx0LUhup66Q09wwy3eIq794tqsR9jkYXEhRuRUHWUYkKkGsqdkV1StnqEv
7XQsszTfYEFyRG7ekWEyZyANz5UnWwP1O89pSz8WUWEp+T3e5XNw8Lal9xVDxiNGmZ7sOMPE6v+f
aE/L5SVjN8794Z2EyI9CBgs/6PnfBcOc7YhmCUQ2Gq8nDkvSQZrS1ly9t0az+HgfZ+vxPlWkPeKC
+zE3Rsqqrqn4nMFWPJ3JGKRji2bwkN4gHtPJormIGsECetw6j27HK9kpYwCXz/KlBCR0/be7li+u
N6J/0gNhohqAsOYnGb6F2GrzTSpgmCdugMHBVbPnMAOJNTTkVOlzalGy8iPNwqZw/tOkbV/NTaH/
P35UjZjfQsim5M+VES5nqSn9IIYk0CV6ylFk635EQsQWPSDvSxBDEMX3yrP7U8a9Ieycqj9uq+E5
9d4ZL1wdWOynu67CiSw8/zmVGNonTKM1Jy4hZL1yNbTKN2RhZF9EXzKJi6xut3ymsLx7tbfTvmBO
DJ3CsHayTyuojiC9IFWBqwRV0elG/IAFAmggb/e6wLAPOMmbjUGrRmuJ29kssL8l8WQ9x246Jib8
57kb9mrt0h9roMV3JVIJ5U8Jfq4830YdGh/7OG3Ek+Z9MrJQ/+k9B9ala3JajYC1fJdMsysEHXOA
WMC/gpewBnXkWjEEc/Jee3IXPK59cbjPC/QLw29gOt45RoqiBYThb5Ou37vxqQuQlPELNM1e8ENR
UQUc4v1FHgGFXygNdLC+v6yX8EjOBpHbFY4/hgRUx67dAyqQFbYWgdlQv8xFqb3/b24WqCtHT9cg
KnGM4ly1BZD5NFZcDkjlgiAHWuiWa3Pjel31eGYjKffkwTQ1fZCSvxwTNRtsE/YOipVbWbVUGYz6
Z/bJDRDuDeArnaoqN4xeQpTngvswVzK5DOLKG1crZ3C9+JtxwGfVwExboZZ4zh7jEziKhaXrelC2
pxqHizvIgHCN2sP0nKa+cGUtjRY2NTSOVLjlUXzQt9FL3oo2q8JHbT2PT/T4mOXDUcDc6ORNHHpU
gjdlpflHXoJ6uKwMb6tDYWO/M+p+BoRtZ/8zX1NsX2VMcglZWbKzcU4FG2aWcOF9UPzSC9PD6IdC
GhrDtat4toyzomU7VV7mZwIVuEYjrIRzUypRIEcVrWqOyZ3H+n+xsliWR8zB8Il4nxB9IbqOOLNa
cNtv8iHzXZ4sKk6qhg/QAYu7R1yqpdF2b0BFeTMAzhAZdtMJhw+Rj7LVAoqqBKrj+MxdznxJOC7k
HVG2aMAVUBoDmzCBMBQD0E0GyJY+m+PblI9nfD2KqWjWK+3zk2hBtRagLhmAbAKqakAyjAkEybHE
MX7t2V+Br6ErhRxtTKOSOaDX/Oy1afWqhiRJhSW9rQ84lq1DGA8asVdaYcZYyTbbeKNV20t1qHbO
t3oJdmnmUSV9o0MsmNeVyfO7+piOKGVI1jtM7byiLEBQITQ/7rKnl3pvnz+V0i7M08D8cQtEdxlm
LYNw8LB3xxx0x+9QTuFJj0xhaiOKuKSEtkHa+05jP2FUi+tLxGwwoLN1AE1UTW3oVhrHVBInskMq
ShWK8KV69BQQ7alaupsHkJkjmNGl5bvyZwID5i9Q9oOpUoJVGT+xLbKSw1vOEJvjhfE5cdYadyxH
wO8ENqJ5hQdRgthQP9AFIPhWuqo8uagYcuAuW+xVHZLLhexAXblHJz0V29oD23IItGOzvHkXArQ0
7cFVjkHPBDE/1f/2J0r6v4ePNB7DlGiK5pMqZLLV9/dO0I9DC+oGO1DnOB3sSOe12CKzHzYkX2vk
G5bijhrDJzMz1PRrbcny6BMX/obZpmDKd2HapZAywLMiuCuFle4oxiktXuXPHxQg0zwJVwRowseQ
klDVtvYz8SIlhfgUO3XEemCyegVBoAmMMteIecddleI+eTKs79mRm7jPEpfbl7LU3/dVF/VLF+xk
B3pIa/nEdkjaN5R/X+B+qhk1zNjyjT+NJiIyZRSZ7plMgUFEAnGbReWkCJr85bLSiprM41FehtqQ
IfAoXyiKLe3jAG6Pg4BFyJDARocQoUAy1xhDdGgAOq8TCPakrkQn5stNwNy7oHPDL3hqjpX9EoHF
0NcT9WNxl2RjByyOwSlyZtK7atwNKvu1QCnv+8hZBYB14jAXAAkPeRQJGBPs/z7MlVxMQbtREv/i
qrGfFTg0uPgq1QdBWCmOBOql18EkZw8qh+WY2s2zyEUa5JMi7zBnicxmmlW+7GYLIakjrHcQLOCe
pNzHd5WD4gDd4vUg8TmCpGgtigSqEDuE7Ort51s/57Qkvry7mYXxWgRLBHElgfBzInbc3IdQODG3
BZnDniOQqxtfFW1ZvuknschHVFevjEJQPmwxpTYWSOcZ9bjQxZr0gyw/MULxFZPZzP9fmxNY018X
p44IRoTMYvpeFwCUI928Yk2c0kP0uKRQ/Kb12mBVLH/nUst7t9IJ39ZHKMBP67bKYW/6fRl/LE4P
B7R7s6ltPBSF4EEEWZvfwt6+ZL/GJ1KIlzpgBtUMEYsWY7q8j7hyH6/TrheUzz7cevv5pwjRi7Qq
S4YuhEA+Pnvg2LyuPzdE6ccXc5Hmp+A0x+xebOtxF3XWvGDN3hLvSCOri/lC2NpHcuOvvknn5DJe
pTw2SyLwK6UjMxHztVZ2zr554dk+melgvHaVvsOyAwdR3+uqTyU8XldZlpK9kPM8xUTvzrAo2BGe
JIxNjgp4wcaPPNvbjBGtXCAmkgAWDhgPG1lUZeh6ptyMwBv6nNfIKk77DTkeSj+mRi3zE4Z5Y8G0
4RD/nwan0p++a/FcA+FJwkhsaZt0By0MKX0IxmS2/MA0PBpkYXMFF9QlZJDCDr33fgJ4v59y9JN6
NMdvMUlhNM8X4qHFQ0gkvBkg77CEf54n+0gQBpJ6bI18/gOdTqL3QxluBKMqtVJj5iZUTE6D8Ldq
rsRPRQOv4I0RYjck1rPIk1rq9nWoeA4nbTmvzcyY0pipTW05bvxl5BiDoAGpgmJZPA9hKeQ3nvIW
lwDTfq/bwIVhoQY2Kbsk7anScADqeqrjHCfU7DurwH4mMmkfEFf3Ee+0h8/8e5BJ7uAaW/9huAMC
SqbryCIpbqYR9Zx9pAPs3LXJPlGuGzPGUUXbPwF3qxFQZblD3M2hI3RknAIgVpCzX6DkLxJTPCOG
nXAf2Ccg+z0LuSxCgW/9jUwVyamWkPmmdktpg0lwhTYnuNebUC+dote2KneDqUFkdz+3VrW563Jf
BRjUpUSOP7HjinPd9QzhWWEzvpBy1LkC4eaH905mGBTjaUkObfqf3S3oQzegtMF13+JtyKCsW19R
eUauzaW+J+45bXcZV19Lhz5c1H9PRRPi4KE8O2ybCleIyfzre6NtsfwNB85QAatn0kfu/XwNrRtr
SpPo8afInhZpAp0lBr3Sj9hY/eJ/0Z1MXwajzsdqJt6dCjIB5/v+Xa/HjK7N8t9KiiVf+QZtp7Pz
QLan7cWCaoGuT7+wHbp3upskVAjd5JoYhrq1ZWsWyS9yK0iOyr0CACKKsfU5M+BFBn7xvw9IGiD2
rvePP+TJvHuiTPQ6T1/WZx4pAgyD67ukA0WFl8MEPsasTI0ErSwbWvW953j34EcmHh3gGbKlo4Sh
QJNRGFPgiWlx3x+Wpp8/1pMJdduiPIaZyoFBScJBQ17jtA8VScTmmvF1Ze/fmR5rHYetdS/KP+RV
DKwoukGX48LqiNTImU9cPGl34nmGi/dccTCWIZnNAlvv2DQtbsSvjKKQ5lU0CBo0FUMZdeJlcJLO
AQMOMqOC8zFb5tKlANjBmHKXBwWdJ9RVu0vvvyUhDadZP29clsS6WXAQEHiUSHF4GIooRE+0+KOU
jsr0ZCN6SjuHN6JWbN+RAN2QjKR5L1arDdhBrnRjjYtCyzeRYS9Q/TIylbh+0iP5stZPFpbowYTx
i+cOmcM1PlHOO7uH5nFqPg/Mquq2uTkkUjxNAE6XxyNI31dSpUckemr9e4glJiZbuOIyRoExK+2Q
blZzJEOcYoHDBfTEbzmYu3tblxmTnBq9deaqdSvRhDn6WdTJv5Vpwq5Bz5aMvKRbqmEsUN7Eba/2
OvPNB60O88ITzjte6ZzY2wVgdg460SBzKkN9QJ/FJPi0KDCvfmWGXtK0QIERODSyoFsiTwXggNpE
jcotDRamk90N24a0hiIxFU5J265Ufxb9+wRyNJirVcaigauRxDT1iBt9BeZOnKA8OjZW5f0Wd2z4
oXvltrTPFZDg5C1YyDhHmSH6ShrZy4m2b/sp2O/ty2yCXTIN6/6YiQMvB2xqfTpB7gDJhuGzJnfQ
BL1bxZeKhqA4sLWdmj0rM72lD35878cNRezY777DElbqxqrYG5OHnIrJ0950JvCnKW7HzvbJMqdY
dIyyoxQrqd4nJ1VdTZ68Dq+hwRTw3GU0QUvEUAlV8VRHhxmQ2mGsYRMVp6FWwPhNToMkYWtYrlyi
wqY44irJztKlyG8xiKNq4yyZG7n9qEb4TL659WI5rARur0IVb6KtWUNqcezOZgszEUbpB+/V+Eiz
iqF1JoMENpAKmZEAHVHB3EpIsbD0/LuxGPyrHV8CkenLxbQERzO+igGk495fPDLs+h6X4TVy7TCZ
97wArFg1qG2GonEeICzQMXrQpVV3rD1D8eULURDpPY0AJweUnuAT7XdGUYLizYa2pf3NRYe3xFj5
kMxXHYYCh+bvzp5fpn7avanZLf0s2xIXQaFePgcJhwI2cWwlb6/xIyLGdfolNYEEDCID1KCy0vgm
/S+ld61MdmJBbgFm9DbanTMGbvofChc/RcTLY2YegUOzefzAzxLj/HOYybX2+JYHx9qf2OmBZx88
iDn8UuTepAzV94U7osOr02ATvScu8RAlURCEW2aSitdJko0Tp+jEC7uZq1jpyDWfunOhMMITCebk
HJvWiSFEYsh2PTbXju8XKyJoBRT1Ol765RLkAngilhxxnCVSFogQERLq/RzFvJOYHvlIPkkkCGCp
3R3cApYLai1+BeGV5EUVEm3fKyqaQflhbxki0AtVRJz4j1QAmrMOFOJcEEjaheWf07oUhByTx6v6
SGYCg52hJm62CUp8qYRcknQIHBpNaXzFZ7bj4u6gs/8G6WLq8zWnxNHVhZCLho4j1tcbLTLTbNkq
xtVBqFHai2jKDyNZzBRK+1EqM2/MprDml3qEY8UmJAFakxEoox6keY3J5oIunDPkbFytMhjThvMW
/5RUzpRw8rYk1X1zpXKYEKodAfnOAltVHXOHekGQWVgQ4qFbN3Fhtwuy2lr8/3l5deBd4/Um/R41
30cHPWncvMH+SUjdAUDBeCah0yyVUWXc01DV8IhgPTa+OUYFR/shf8U6pi0YJwTpb7mDP0WC6YIu
PzxJIskaSc5F0IrVSodksSSIRLzZI1GYt/atcy2DRq0Yj4ykZGvG3Zff7loeZJ6F2tKYxfY/+xuP
RXMpCDtNNoBb6tk6HdUeroQWHU3l8ba1XTkQWzO5HvdOZjGquIc75JqekLjb6LyGWrb7hjKd5t1z
FnUGDgkktnHldV7Q6qCLBJNjVEC6Z7Ll/yusflgp9hA+vVhazzYQE0RqpzzVDCXxdjTgaIfAMwzx
GaVdHYxbmloffOXxVbmqGjbJSgsI5+7rQvWeTCIyGXvOsO3/ifWpj/tX4rniq3UPCSpcthR4NFLx
+LzESrbKyFYinR8uZ36qPE2wasbbQMFrDkyKJJPlWAjLXUhZMeOo9TVzgOR7GiLGbMtM9akXdl9F
80QbiBgLrpo0FX613EGLoOh3F0ZRPqlmHFV7gC12gfMBbmHkMMAUpTNi6L3YH82xClvuHq/kAiRY
u/91uiF4hyzqT3knvP8f02QcX+gFPz9rFclYv/ZE4A1CnAnjcyBZLm6VJJEmodrJAyFwH5rmsBe8
ZVxmR1UBa4vXFRYhDzmRFilLCV3axJpGQxswlVGRaeuuBWyWf24chhNdPzfkggfxQHMAG8gDlrQe
gO0W0wtCqxjYnMPRnu67/tmQl814CDt7GzBB8VEjMGE/cKnjQ+hEJf3XJL3yHg2CCxiEUVW8xYy4
Wc3U77Sz55sZVzzWMBh5fhilHHwxSgvwMTEdUiei9hleOTRFhYSM+idnUzIEQkKo2fs53vPQApZ5
WL1JPs+qBuTa+I88veYLfHMvSf6J6xlPXmHxwofq7xYy7tdvaoMD1N8O0KMRRN6vFK0j/1A+F6Dq
/PMCxdEAz/ADtq5/iohY0QfQfuh1NWeIqMA3TBXLFfowFXceXHMPt7+ZM1XtqQcCGtHK+a4ZqEdU
X8VGfWEX1eAD6+a5M1dR2V9VGOf8Vcoe7PBGQiT3Z97vz10Na/gKi6iFMierQdoWzc4RC4k+4cJV
YYjHR79PNTRq7NbsYMLefB1BYG3yFu7AvynSpceJv17ccZlQz2C1UmyAavGRqbmBd6i8segqBw6T
536tZKDsn06Z8MuNk2+V/KcN2OLg96//hqXU6+VPDHOXNwu742SJKgjrHcuCNxRoDUnmMe59IXti
mRrhhTWWd4mQ8XTPq1TL6JkeE1uMRLJwNYsTRFDHE5eu0HKJiWCdfGHEP1GdTqpVfN7sCX2l++Qy
2c6dGlBukP5ggs03BKxvf4axswX/tSSIOqVRxY+ENUGh9eDWdPlVeurqavg8+8iHKOyP/5zNRtEE
alJOFc1utE6T5lDt4BBquzgYClaQkR0d1DIYhmKzkvSmyzVWzZ2PgBHdLInKlgTxFK9WxiKLschd
l+3bi3BfDM0sb6XrU1avtgxEvr1WIRH1tKnFh4r2p5PASx4hegJNkUiSion/2UX0VA6F2LI8FZuL
YgkHInX1iLLt24vUbzoFO2vEVqxyBs+x0NYF9Yvs7z91J4xYNTMzcwxyTA==
`protect end_protected

