

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dqq2ej+LHAswGLNpyi2BwMJ4URtm/h34HwSY5qyFGcps40U3/VN8WKFwHX37+XfGZChHdZC401n2
ZJyf0uELfA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RShplIv4IYGmj4hmPadlbhdpa4eXDDQJnDlnCbKU8o5c8V67SplZMW55cCw83AgbV+E4+0de3dh2
OewneR7qBBfHbEaasIMiCU+zicwJbNM9VmcXiohAYKq3Jg09b21wgUWnQjizooGjaKEjrwAf7l5n
0IFKkSATJTBklshviAQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
doH6vzjo8znCTuVASkkAHdn/+Lqszo8VV/fIaCg6/PKdzVlWSqotQ8QksPb17wveo6mrpVhle1T7
Ab/aaE9I9n4vMXfI/FWx1z3lglwq03QllPp4tizM/2losc/kPKWIjsGwAq1KyC1e4r3jOXEn5vSW
wAG6t+dDeOAro7RHFvJp5WNrqaw9ZsPGHES5alp7+i1zKM2A5fW3oszndsJYrbNt2o0DhzKvTBJe
pWACtYic/6CWArHvZ1hBW+NeExIHbF8agw6nValUyGbrgAgoYKvgt+O2td2xISQDqanZU5ezYx0k
TdAWuo2F+ptoHYLgvzlbDnbpaYfltlwCiHeG7g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
csfgTxr/fVeKtQdd3D1aAHu2gzw+CL8t29x2K8aPw9uZ+LarpUYk7LqFUy6b5Sl1OdJTAvVuQG9n
5euFlEghCMUBQ5Nd/fPjuJkThGKoBDPPfcptYVqHN93OBm3eZXgxire2pFol7b2/KhoVoBckFmFu
z+xA86qPFh0t/6hOrEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iWrYYlUsjF3sHqYa1YvLKfZWmztT7d+xNuYY9994lyI+KXcZqgZrwGg41h1Tjrz690obWegSp1/g
FB0dDXfIUiHiYD2/yK1JWR09FXSTykMHQFAgkUCT2FR64CxYjKEn4kixQsxvzded+m8oQLtN/sKO
huWNyOla5moYPLYi3ONKXIqIpiP8lBsvjVWrmrNv5LE3TVAC4aypQQK4UiWqxM5N8C6AsQZbsh1D
wOuA6RwWzU11ZwG/y66u76tMNNdkDF55Z85dtQpn9re7X0RzPcoTUqEAT/dYJI6s4KqEqLik5x7W
FZIXXtdazPlz9KjsPwx1cFU6reG0ILErlZIf4g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6336)
`protect data_block
2BqmOY6mJLP2OD8oPNabFAfJkGscfnwLz2+jzHhKm9p1jke0TBAsfs8azMo+hbiGeDZyeoD+yxFN
6OJmloGaTgMX+fD89DGcEFEvfTnD7d2j6/CU0oi3K8YkvUiNRf+WXc9LBRteF47+sNgMv/8QdYIM
A0eiJxID+bOs5QkZi7Pb/Fr6YN3ZpHI4k2IUkNq+jTBFh22gkhP5p7CerrC+5CjG8UAbhEGyXHJ0
xtWugo4XUeDtvnp8ts/SB2BAVMtYGMhGfA/oJKcQ0//cS1oW/WL+ncSf5r8GhDkR8slK3xs+jmgm
44fXzRatyMX5fuxTGNoMJH4grYZCkIZEThsETcffl6aExiWdN6qlcylHpGtMRpBJPfHIgxT5hLKJ
Qelzs26GKn4hEv271pXsRhl/qWKqISvpU6ZxS6bCiBaK7GvDMrVQn5o87QaZULSY3OO0ggUYVv0Y
Q6mRStEmUYpa/xeXJ9/kDqVlyoi+pN+GQZyro6wBPjpaFdiBUbV1lgI8h0HldXqGxhsJMgUA4bxE
biqaREraxOz8csTSDAQdWdw0zCzjo41g/dl1yXJRodMT/p0zn5nms9wJa6H/QNZPhc8uLmED+wTM
rWEXcAQcSew39+7AomrjchLVem/+0PSwLIliR3yAN+qaNCIDJVLw1bIku6ttm9xf/XJSKSRWPIto
uZAhMus41IKx+t7xcpOSFtmg2hcbb3kJw9GGl53rJQsf4drvmmLcWDzWnqN8Ph0x1wVPRvWQ0W1n
X/JTqs1Z5EOT6hzFmOkeEu3bUT/S5y4YPBRc5T8wE406JkxpeTw1z0u9DFaM2UHz9A/tlUtrDsa/
DAFVnXzES2L/aZnvr4j9EFhivUsy28iTKCBFo0gZ0Ah07rZlKxvrZ23C7x8jbQDSFQ85Z0A9xBlE
M7IoxhQKXf03LYTrdFwTi34qDCEIAZ6v5y7YIvSnRIK9+cveKi0WoWQ1lbLRrbrwCAMttokXbfTL
peMVW9Lw7wubKdACNwhJ+ygSws6WZFHAijiiUU5M3vtHjvE7saE6EYhbK7a6I30qN77I02KMcsfA
AXx1E9beT3DNE1B8RGvxd3dfpoCC0IbLrzlrSD9aQvllqo9WwiDZvlXt5L/dT9FFg3Vf3dnNhgVu
fIwtsJO83HSMdMsM8qzGNmlhRXj4K/hh8Kd0Wvd+/ZeOeJVVjCu7xWf9io6XcGIwgMV/agtHNAD3
qDdFvuxwt0KSTePl76joMDgU2lewL99JbzOrDA075Aibiyn5sjuKq1M51/N9mVotVV7SW5I4orJu
0Gso7lRk78CDLfZo7D6Gz4caGD1UjcMwPySYicr9u9MCKT3xjgFcLUjSD+vurdoxetXrcfInEtJ5
wrsUZUhhYs6WTNRsCMk+T5YcBHEMXOZ6WqMn8scmSBnkxXrL4y/LVNCSaA1rq/eZOJatjRxfxBvF
5UUnEPF3x23F7ca8SbAvkX/hQladDnVXoloOvl/0GDorYWhiXSAvbEK4ighWH7kJh78go+l6gvyD
C4bC3XxYP/ZwQO1qLurINXXq+ZjVucdvsTtzSVP+7kkbc5rLgjf6hFFPlUROjdEPJnj27vNBkUYC
/d7QRCyH4HPYYbAuAMLJ9ZTgpOgDKsJXa1pvQLUt2Eyew5QzeVx26GrYdTom7eWGhv/i5lbOrnhq
5EILTxBlq7KTPNzx1T/KNXIxfBfEu9/Tkvdf7TzaT6ETiFfqxWVKi6NLioxpYCL4xNRpPFJdBdi9
sDLRRjxh0TPfBNzbV5DaxT9X2uxHKjFCBTwYi2yfXBI2+akc2DdHSMfsA/38e3xE2VLR/qAoVeLV
pPFHHWDuv3QIItoq9ZdVf7AbTVJ1qhwIWW98qUGJltRo/cuV72rQA4wrMhNHElA+JdBCQOu85Qm6
dt9/HRyc0/eJ8c6BN2usHYDNLVa3k+0j8Sknm1WJ51goti1jp6QWMxRtR8p1xKNxuc/Wz05jcdI+
tnVhauRjMe7Z6j24bJFl2E2KSo8LdvKddxBzPjUpVkpBDIS7pAf8aWUIbXdHPoTUicQ1gYmiV3rH
UssoaA0v0Gzb1hfX0/NXN9qp3vkOK5dQbmIWNekYSdgqGZoiJbmsElhh1EOJvxamsu9+2P8GfpqF
3yTg7cTGkwwodonbCSHrl4ldoKMGIXYmBBBpbX1giFCANXd4r/+F+465TcMHwWGIH3PC0gfKprsw
tuLRv1Ll3aAzZ0Ib+b3SteKqJ+tutUfQcg4GSheIB4r3SVLnSH6zGrjds2cCg+mV0NR3bna8I4VT
YPvan9rmc4UuH2gEQz3b1/4IS2dI4ZTcM2ZJEpuD3ZYNxeM8oOBCVZj/2XGxLmmD8Tk20dFs/Uld
KbgxaCV/aS3QE05qhqJQcOlW+7uFJdaBtMyFQ7ghq+rJkaYQRuRzujfEdTwKSHb7qo3OHUY4slNH
fSOLW3GkejaB51S4ZSQqsaKWy/HPjOEb+HRAJ+2hKJ4bI4+wuuFuHRu99GDKxds50u4yiwqLPHnz
UHK641Z21c6sPU6Csc30WMmOrDQjIYI9nec1GnfJbmw1gd3jwd5UXQswiY5VwI7nfsENKVcU246P
MNFCZd5y8iRkgmLc4IB6ps15YlpxxOoAMbnEJr3flIWMIjabAi19+Ibv1A6dRGb7wqASqT1Nucmj
GKM9nB5aLzI+nhInC5zeiXyFP0MT4icY8r09otUGsfGfBoJsjvzwq4GphwK5igefSEP+B4UqJ6Np
KuGs93NTHtr0D0I+Sa/g5TJT69YrDsZuaFGOG2Ou9VQG9jGXVJk/mwkolZMMMUBsYxc5S045epS5
TaMZiik3iJa1zo+HFitIDmx9xjlrZxm8g7t6eNy13B8cBJCwTwNtVCYHI5U5xqym2fb3wXleDDIT
tY50ZqA30b8e0E0JAA8r8q9oiJkwhyCJc6gvV07/3LWspegVmsewhHAN4XHXPmPwOoZdOTSZnZ8b
Vmsot8ptzhAg6sFp9XU0yi1g5bn6cZiwtGSXScqLMkYAXr+VuFLEWzppVasP1z/N9wDo5Yj8cjSS
LB2Wcuo6odz+m+JRXEi4hj9WvFK4oRccZ7+wi/AkRj3RgtxVwErEoLufRuryeqQK7d9KlVLqzMdM
px0Ede+Re7zkEUoMBMOke0SMp3mBemkcF4tFgJtBiYtC8mD3zx/9YG5qyNetA/n6rkRYmerFTJNA
khwJ+/mec95FQ6CFJH9PFoX3lj9LNMEBICX6ryMk+/P6G2nTb4OQEp8kgmHCyrb4GJySIIQmQY2v
uDwZ0hlcOWVgGpuLblgxfy0Bz2NMoOfcGFLGAjk539nb0rvDqthDm45GTI1JZM2dITy7PRX96jT6
dv/K+FibIEjU3k1fxWdmvbCXfzy+Y94TtelouRcIMAJAJ2VnsvbewJ+fZX1Vc4JQIpEuLcSRxFAx
ZZB3iYXJ+fUwKK1UtVnnfY3gpESu/rcNrW362/nbCvhbOemufRhSHLLt0QqkNMrB7u+fDtuD2yFf
YmUieFDIwLdt7jSZtElBdVa7hOpl7l6DRsSdiua4ljsUQSV3+vs8SzVnNfXtLDy+xhF2wxMKtrKZ
kdG4Va0aZyieSmC2mpX5eg9fJx0wvUumnYT7jKnpGZmncUlZRqMm5xUL7sOSn6Vds7Jt3agq8xaE
g8k1OjSvOce/gIBZGSGZWb5VXxz9PbY8OcE0/iq7PErG1V0mN5tOSBKE5Qq9TTv0HqECU+5a2NtA
vU3p6TEzpi4FCCLv+q+SAWoT/TAQ7oLuMHzo35cvJSH5Jb1fgarPh5uDzoHtKbWI8C3LV/UcfBsY
t4xUPlVgKDqp+lED9lNmCVDVTJq1ZTAVfg0xMi+pEgxW9fKbQCrF61HdTyfrthmbBmbAhqL1DC4L
1Yay9amcJ8Sk80761LOGnpZwLKspwikibYms/HupH7FEu1LF3ohv2ce3jw4vvAvhFidlxZTWTp/+
O67onLWLnXBcPbGH1VjxAvEixgOS5FEp9UH1g97lwUuv4hyhDJMwRE8+idQ9obkVSBu7BCb+xvI6
zGMeTZb5iYXmb6nx8/rPIPwZUpb9pkltLn1ECg8eBKK4+IXFjBtKLjfvFjBWPmymf19DjdqeW6Bk
oFiXq1V0XtiwwAkHNssIDZx707lStF3FzuBY2DddGOL4dRqvF6bSuXFhppkBtGO7CDpaXLr7P24Y
tOajv7Hty39b+cqPiiaPEeuwK87+U0ic2AIEs/YIDIWB3a77okrOzRXpbvcoNZ0qHN/+5xj++vp0
UCSFFV0anPoB+9Ckn06m59pu4aoVvdBGPHnIW6Vl4d8P1h4boLPuz79UST3qvwe4ROp1g+WndyAq
m1WPy8ma9Fe2+4E7h9bT4aZk5yKLN7qNIddKDInCf9I83HuBp2WT/aYemrVibfHqgQevvxTX/MPN
BNV2udfeLPvDD2nKnjyIUGBXM2/5CcXaD4Q+aDf39w5ileCYsMSPammUsJZIb3JNNJQrhJca1ZeD
+BJqWYpaVQHDHwr/UMbqnvdDGR8oDNCG9w5KFl+3tfpfIhV6VUMsJkIzScelsRSrbrqgnfuIUIYn
M+IAntdYBpxZJCWyR0H1QyZu88P6QJU1krOaTwS9TzKEDD+cXh8jfhnB2qI4IC1BY7fK4u4PxX4o
IS1bxtDvU0tThO37j2q5Ropt3pvfSEGTztCdU9oBRWF+sqBXFEkevRwCzsfw++0otIE1StBmVwCe
S1wHkeaW182eaVBbLv+4cxXGWbywLRsJwycIu9HzIX1Y0bIEkQ62D98CtOXMxCjhSidSH+ERuSEz
g26Lh7whKW/ibGmRKeoMJGGS5lwly8Z2uOoHdo1DGwZt9YT+5RUwg/yghvaP2VuYm8Jen3DS5wwv
OlXrym8JIh94sbiDJ5K0xDmJSPOInTlywCG1WKkx2uWo8hMSD4STs+xyDRMxe370SuAYdzXikTzV
uQwtcYnaN4oeM5JACiG0s4lIFmJrbr6cSHcOEpXsMUdUk6nWrf4dnHxRKhPQRgUjruB1SNFnc742
lFInppNeDfNUrQNt3FMUcLsAvkr9nOl7Ze7Tv+wEZD2GQCTiHS0DVdpA91o2sEZt5fTotkeU4oAQ
4u4JdrVFd40Vx5maswsfeVEcuk7RQp97zjQ3YPogSvs7+rm5foMjjsueYNQ5v1O7thiaZmGqGanV
hG+LfRbpBvuHrAoAEsqYxt1UuPzZYFSYu/PkNTPceDihw+NNP3vjPVp1LAaHA0u0MitfqJV1sS1/
LiAf+2NyHUjU6IYu6wcv9Qdqpp12HFl+f06JeAadDQW1vZRPRie36KVNy+24G90Ge1MLTAKVHtey
zUdpDBr2nek6tM3VXrzDxITDrqLjJBiXw4mr5lb+fee2yMF6rPTZwjUfAQkVpenOGTtwTCKMb3T8
eV8kj6T6+VuZEmjDB+/RP7lbsJJp9i5Hgrh9JEsfp+4UsGJ9hDjZ4skXDGkgKC5ZhlEKK+Gg6/VC
bTrkGzFyDtkRlvxskZeCDFvYVfoYaan1A3FqjNoqOFqCY7kvZR1M94ysoyYynRe1J+TqNFA9NpSK
d+WOjGKgxwtuVRu4AsjSNmPpsrea5DNO+asYEylBW2AjV0sNI+BqW1qxI7LQ5z7aQFWTOtcdWbu4
v7Lk07tgNhTx9+mgZMu3WW0pI59thFVh7+WxBNXb4thgn65gT3F5lXMa1INjBwx1xX512qNeyfjG
g4iFBOpIEMxIxQChywP7GGEasZH4Fa8jzo0SHtC1OJY9FrX0/OQdWejO85CyijjIe1VOV8+KK841
S5T9uxoxYOXCOrwKKfm1I8NUatH+Oxk4JZWeskOTNCygEQNy8XUPjNj29owRKcKXGrArE1/hDjCo
E1iubHZVoDR7+RLC5UUYgcWjy4MVkWMVSJMTIqSHptkdmgZTaxK0EcDIaVRSh6s9EHjBZcwuWQbq
S9xDTjyXjMZkKPYrEfyEZGakVkwFiqN30A9USE5z5gHDF59Jt5PR3wtuK/SisrmZYih4ZJgP6BhS
Fz5oxD77a2MkoZBfoWbiBVEwPhCsoGxeMQsqeLAuJICHXLBfsrUT7kaTUrl5wEeZVw1+g4wpc5ys
hw0F6oCJY+DYXXDpWDHbKsWd2ff6PdGmS4mlEDx0ZMyoIB1mhzzP846Abw5HfVPCWXS26+FBcAOS
Nc0PTUcuqupr6N22kmaTQTDHDslhdfwkJQvvArVUAGmLUvbuO9f9e1L5KS4M7yt9MVi+xLFr5nw6
Ubs5pLahuNHyltUI2mPpf9017ACbm26x+Azeo0tejoSb4wz4MKtoa2BuFCw88et1K9NCdBGxiVk6
UF/HIZgcKjEHp/LTafa5sCLvh93Z/jUdfcV0LoLvLU6pm+1kphadTy81+WowutPx+nH3LAZc5QMK
2Z1F3PpavBZpiyAuj4gyCc/GBFwH9ZaVvQLGD7xrGyQqvUpqcescU52IjjQKF75Bte7Wk7uA3BY2
21Lt56VqFJX6lbuotY6apEJshGNVs4VmDIjZwJEVpONTf5M//vViPITIyb6l6+T9OH1ndtVHiogS
5dJmGaspN84atzUbYThyJuSD1cMDgpqgbipB0RYn0pplv7xjkh2a4p/qTl2Jr0bjlQPrxkzt4dem
2z0DegnLduL3E9YwbOBJL1Lf5hLQnFMcjaNGebUYisG6QJQQwDw8xlLXvS6bYx/pVfYV14E1BuCq
BsQXS3ZJ3H7QDAYK/kADhsL2uuM3CORYImSWOd4XXNqCNCOLTUf6PnllWUtwzgguLn5Pm7yFoV7Q
9Ve49DDMOcNBaP6g6t/FFQpmsF91waIadXRuEAxvkjy/XJwnndo2QkH1o+NVi1V4lDPs5M3Mz5V2
SnTBwRjMJsUPWqU4hqhuVri65ARwzRNdM+pYBzDzXiE6mu0Tt+czRNaz94MsZFctcNCYyJmkdSRa
RypG4IZjd+QvKF0px3gp03ueHYxlQ2+f/B4tFgdIEwBHgeI0atRx5dSrDqMtheElmx1OSk6IODHy
S6pzERcDaiZZvcqXdja6xIUL/+GUxz5hkeMZ9EnlIAPiPPrDlZxkPpBFQ+nFNBWvUB9gcJmFazCJ
oKO9vB6U4P2+h5d+nx8cNycbWPQh+OzsK/o7/J4uukk8fvnersM62yHM/zjQINzoXftSIl4674eZ
RwR/+V20J7elx+dcq4oLYlwAowXYXgPpyoyZEJxHSgv1dtFPOHZ/VZMNYPwzn+QohWCLp2vK9HPo
Ga0I6R54AW1GNza67T9q1CyWluKUX1zMSp8RbiQpO4jaMwpcfDXLUU99Cti9kedpVIG8JEKSxTfu
LRz4H7JXrFUB8ZVcnS81gd5YhcLg0j7Sj5BrxSF7x3C7hpXEVHZ0TIHdpnjnjMrKCduhjFS7xtQh
BUAVCzmRe/TOSMqqIt/f2xUZADNirOKBNq/gmw2mHWbrVjp8HeI/ZEPK0oZ/8VbutYnt28tw+DhU
3Ac2LA9jFi2EqZKL4+VZoie73RYxDRoi0q2z+2ovDBYQHFpc3It4co0yMZ5mfZXCLpB9fPx/nNU5
FN7j3oombfMb3S5iF3hMGi/DFqol7liJHwBjSFFthScTi1bHbJ0Aif2aQJGEojqo218RblDW33t3
bvn7ES1Vggx/pETURogprU7z5x8JfoBSeBpVMfhu9xWRNClGZ7pbv94h2qiibro14vcQLdv6q8B0
DOkjWuuecSmrB4RkO1iJYUt15GlF8VbbBny87GpHEiksf0k2HywhwAv9b8amXBcGVyabcOE9MUfH
khns0IDoywm2QIuqlyoHOgENsIWnbYBY4I9//prb/WAHlukUHlBtkD4q3XGzLNZE8U6cQTUYESKu
EFEbpJKcPiFO9lkZvKW/xPpaptyrg/jplVncXcSyZ9ClavYkeTEPGkjuH8wTHLPVMc3XeLvpWWUC
0paLIhfgd1VdpmPTcrymuGP/3kcIm0436EwHtm44/e1cdRN8f/XHdzCd7WQE67TcOobT7fPSBRYQ
cEzMoeMaPioyZdo1G3DHyWHlhGgyTpEngDHNZY1LH3G1+G0U1w3MwvTZaRf9auoEFVvMdP1eMrFu
GYQXQI/sVIwFmE7AQg2x82tDI26Qo16OndlyGYRQFbxLlb/NdhQ4oNuLr4+YrJbfpbq4qrpPy+H1
ueCcg3LBVCXFQhkSKlpDOcdj7TseqabATVjm6xDCF2Ryi0tvRPcfY8ROiMDNa45zZwCjOdIKc+1+
ZwlMsQ41Ar4GZj6RBS3sd4t6j0MTIFJ/xLJzdDNneRzIRStDWoEcRK/bx+tNAHnBd7xJ00Dy9bVf
0fvKrFutGem852yk81QzA+/AMZRTXQkKO7OgeQSIh1d8B69+sGzL9zXgBB41oJO1UbRKIl+Ejzzf
TGt/TvV7YwqZQq6PN3Qi/MA/0JSGp2sMZxDZ79PdrnWCm20sf6zSKrWVIzavcKPNvoUaJyQHz5ju
ZPoY+fYT+KgU
`protect end_protected

