

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jm7pyByDrqpI4tkfO/xf7lmqS5TZ7qYRErFr0jmmE8foSFu+eTk02v/3RjgVn1TrEG87GmvFOJV3
1tbeZ+/zQw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
goD6KB7ZGiMU0qIlT7vnAeRuUN8V5+l6EW7ihXwx1ij1lq+kam/gBRw6CNRo5IxApJRPi0JF9qee
YmZeuBwLDvRABMMsMO8pOTJXA7+PBAPaE3oE4emVIzIlySvLHgR5DQiffOav7u7lWIzDoPEsLFn4
h3+i4GX451c4jB1Rjw0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yeqT//HgCoVczVBw9h+Y6MkIiNON6RgWk8BfMJl7QnKCk5MC5tAhfLpWSG1orQ1tjwUZykL1H9FL
vt5Lzozoe3ULrW5fhCtS/6PGXwAnUPe/7jLWtVZ6P4+P9kWHrRNvcU8LXMEFK6pBseVdQxrSpRx5
1Tbl4MLQEnqTeBjM2FtX15teDLydhuY8Jd6Ppe8t2t9vagQsPOJKVFIDZtHrdvOi3opbn/k5NZkd
k4lahNT5G3GA5ye+TMaACFyQFUnqL1lEUdML85grLjNA2Nd/k2UhZza3Tfcd7EijxPuXz7Azh+aD
IbOREYnlP8qIWVrYSQlIf7o1VO0SY9xt8d1OiQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc0H4EYvS/dBH3PYciPsNxaY7mApQiheeHaDQ+O72xOYGYn/5oCOrxdvgcskbJOAKEw1omtNhBUu
w/LFh4L/XwdUQRn47L4SeWFZwYG/0D/ioY6/0sknGV4D/cFD4sRWVNklXJdUchx3ANgXOzsIn5Og
P1ojtQ9StVPwCpo7154=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IereCDRaESEXm7TKAg3i63eV4h3mrNPCmUUc/xXa+mXe3ubCtmOzNc1mEyz9MQBgh7Qjq3a4yKLb
gUJxz/zSjq0bmIAuYI+caUfvWZvM7k5rE+IazjEsVRe2nULXICkI6GRzXHyL2+B9/rf+U4ilYZLh
vpEDixGVhnlaoVxfU6LUOkrXC18tBbHG214sL3j8PjzjPQrckKWiOblWgvMFwrt+U6u608WCyqTH
smIb0RxXA2qqYhbpxdv9h4b5jlGCAYPO9+ttCBDauSA5uc15XNiVPXb61CYsvfXmrgmPJGzSYXfA
QSlqNLOZ82+fBKxRPNdQKbqbEDnQavJAhWD3WA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6464)
`protect data_block
L8XTOMalkmbe9wewWn0QMFOMlgwPq+jHWl/DKd4vZ04vfdZwcrDpX09BXyEaLHLqPqbWIWRGlRoZ
tZO9dzDEHg5K1ynQdbkkQXaWIoqacWiGd7Eyy6CbhsdBbLsNSUEVS0PPDwVGviOo0u/gq40pXOD9
SzDF7q9H5IjIvzX2liA0CC8Cd65EUA8CvtMr7DqPSkXX1NvDcfN1T/T0EdFFYq23ik4EBP31Lqo0
lsuBLznavjsivTaw+/JKqA4gT737O1t8KZ1ZgBT/9+L4Sq3wld+1drRrOVAt67heZQ2csWTo6fqe
14gUnXApYn0RzTy7UFLwIWhLsT93AXgkXrPJ636U90KfPkooPPFBpBeQNxNC9Sz8Y3rKcdnmAt/v
YlqOPu3qcOwav3GRn8UNUz5bI2T+tKI4SrNCoM2ks30uQWkM8JxvR2nBrxeWmIZPzqQm+vdCL94/
HsiarM16HHYD/5ef7myTrRd/tMCAX/rWQNMVRUNjexN1f+fO5Yar2j93nYutotvLE9iJxIKv7pnk
Hcs51ua+Vo2yUuJinIHzk+OQQDg37iZQ0LYhh3hsIqv5By1ZmAzJCubhIxx07zD9KWbgpiEcBodc
L0vw7caHRVIVvQesAmruME2gVND29r6glYN8oiC6QCi45bJIvUJgPTSQqKx7FXn6HouyqfklmJVM
jhQ+K+Q3ddHMofATbqm8fvYiZpl8Q8N9V5gEvz20Csfn4pTcdjXrQXaHdU575bpA6ETH+kJsuXZx
97mZZTTVulqaSNOTcddQmoiEOowqAyO0CHEQaKggJucsYS7XX0+GldEIb8fNqJmbYRjFEmYLtJeJ
bgJ1sFW6tUVzqe4Lxs8Z4V59CliDpH9OPiTx4Aiz1EYdQHoTcSUjO5ErJn9yJNKTpAhoQZp119HO
V8eby+8Xjii0APOcqB7Hg44IgSBQ4cEWRMiDwx63vuEt8nW7BS6AHYv5qcPpDcKG7/zHb9tXu8XS
S7ihpvEym4/gs04Z5OZQQEfnglvk0l+Os9pP/MaQ99aOHU49EAH79Q2GSALaTNkEi3J5GgtPtK+9
90yhpA2ZNzn7ly7TXd6euTu5sPqhmumGUYIU42s93EBrpLLUu8H+xmJUjl1Rpn/Mtgh8vU2m02pU
vYPoBzL3rHv73mzlSzPcL2Ii12lGctaJ4oikBP9zdZq+/GKOyYdC3HrEH+4mpBCY+06RUX12qbLQ
ICflcbTLBJgh0cDqhP6txTqKbiLhe9XF2Gs5cE4Bsio4jJg7FdV+j4hpWJOYRbgBxd0M5wP3xdxh
HZIqhnfulCM/CE3qXxbQvEAL4+hM8J7HGZbRSHmupB+/0yOFcoKR7n7nP8/n0YD9SkRckUHeS3Y0
CHqKSx+Q3bbk2Dh/rIzX4qUzr+o5CnR4KKa8zLrit5XzrfLhu5y8vTAElXddVE9Imo/HpJjMIalD
O16GDXB5S7BsclJGj7IvUF6THBWFLI8UYbKdOhKXZmbAOUePgwBoVrp3x1GnrDErOCwq94XtonBG
7Fib9SpKP5gySQls1+NOtSHqxMaHDIXliiwzu/GzeFCfcio/HjiXryAkfKt1t4K0xUuLrmG8zwq3
02nk8BUDPXhlPv7AD3quYYwiJp1PuCbCf8kPtsCAYwY2h4CDl/StCMXMhq4LsDSyueUSAbIurFYY
PFJkjU01SGMQ6+Mt+0VG0zFXfHVtQhD+Uy1BeWx23bGU4jAAwH8U5c/B+AHUCnRl7KI0rkR6KceP
tNuNpf0IgXdiboB7mWJvS1q+HrDdYkv1JsqEMe3/sg1AcvAQ0fzId96L8y6eX2Q+OtLgkpkBvo47
NmsobTdMZYf2OhjajIevogTeS2QbiGSytWl+t9og9Dpx7B4JbauV+2mntXwqjiKJgIFH3JktJOO1
mPmfc25heQLkoXiUgknON2cbccl6YLgfP/1AGt2zgPp0IUUUHce2p39mQHf7kUWXFT4bRQpaddJH
jPzR0wkOD5SvlcLDI5D2kzsyl/fPuFvzUQtQCwPEHyr+uO34VdbPFYXDZ2+h+IniNStUPuhh10Vf
ZMIaKqzS0QrwCa+brgfyqMvGlmGo1U3LPPnLbD7Mu4UihcWkZTXJi6fCDZaW3LtidLb7xHgZkk8A
gB0j0XVsCnJzcq/73MfCYAPwdgL4ufklxml0MGbpsmnnSWnhoto8ttsKsoO6co+ngDXiKqmysCTp
mcLJO59+OFOXrE53e4jWJuk0YPMcynpr+b1t0KiWnp0N5yXK5L9ZaiEyX4e6MryoXkEw5WnNnzJN
UnVttyPzu1EEfzplg8YA079i3KptxndeFQbrfGI3tW6JLtI/BwfON1bEIaG0u9npmcJwsTzbwIP3
IKXIbLobmGjp14DoqsZosYEmniLCxBKHJaNtJOCRo0TRmNe0t52aVNfluakgajbmD7e0E9aYwizl
mIAQfI3hwkzVDDlA+9LsXrxxcDF13BxrYVIjM9gLmnJUtJAprFzRWRIJdsbaRczcZXwYMouOjF30
2UgnR734cX7scYKF6joizO5EgYcwSXcPkJBh+PtHjj54Q7O32F4rvtaWPSaw+ud9zZlRCbkR6EZg
S0Zob07EGxGYXNzNSagmoPrknxoVv9kKzWaGvdzHirxruB2A3uEKL3h/eeOof+l2tSC+OoZ6QPCX
I5SqAeUUZElkbFv/AkB/zoquVfdkvBfD7fzgvB3e5GgfS06vJDHoyUmKL/Qom7UpFh7pf0x2QX/8
GI/0z+aVb3KLLBmzuCJKyzHcOnkXoLIbsQWFpbk0YPbqiH9MvR9+YntEvIXI2lIXOceY525z+THe
etNWZZLvdnDsLyj1nrXKDC2JrdZmvexqrMHz8myViCDLR3UDeZXZhySy7fo/UsAfWZwh2mnERxps
KfnoGek2hRM1/xe0aJrYAuTTFHDWMZBDAjex/CbjBysVb9KlU/GpSKOteGZPAAC2bHPnibM5zPsv
yMeVM4OqZlxCPGrXkSRTM6gYzQJYvuSEzuhPSQBEp22WqU8MDO1CKMJ8CQ5PEwzSUUMD+KVUgg2X
rvo7tvgDE7hmaSBhHFJQUtwr0XbYmp+S2tKMddHmPgydMCnFwSibf6hgTr6CKgA5u49LOf6eYK/Q
Y1vnkTGE/uXFA5/hDNBGyfFxyJcS+9Zybe8P0pT+W38YGc1vHL7/2Hkysl/8YupWwfaZ6hX5/FqH
k4F0Xrrn8TLVWWl1Rd602e/iwfh6iV3YPqWjB2/sVmGTRfFU6MpGfYQ2UsQuiT2OYgOg53n51/CN
OUuDb8dYfaw+rx5TRop7rnunuFDe5HBrzHXBw8zuhAkIur5xGorzRqR8RN277UKyGQ3E/wfLYoUB
E7Ytx9fm5RZUioayGFPfZQczewyZ2ffCoqkzkIobDmlP34XCJ4jIFc2ca1yeTEwCFmKaXw4Nqth5
Vdxi8Xyf4Nlk6Ok8xn1dACR9upSQFZXwwRUYxQCbk+kmQCe4VriRdPW1xktKKBfzbT5FJYkeMSat
aKQmtMHnyCundYYhXNWBFY7YU1UjMsrtO7Y+gkqj+crZe30Eikcdk9mmzbkvGkpzWubo4df0jt12
8OAFrFPdr5aq9SZ/7KV8SepRceCDYpGaO/FeBXBmOYyaLSNFrxfdHscRiu3dJntJR7x1/E6rFmrY
hTEHQeSC4aTbF53654cw8PeMoi+l6p/An4d9txAT+7RAOHmMQxmNIjSeQSSpL3lRLFk/LUTi+L7d
TY1OLlD6GS/38/7HGAmNuAHvcy9sAciazok6fI6cc0PLFmG4iTAUvCNfB/rMIqhSDq8meNvU/c3O
U0VXqDGEMR0j0CyOLBqrAL6H6BtjVfvDKeYzDzLpXKGNfQC75KB0Dv+guDuqijn5thQBoR7MTpBa
8lDsO4NlOJhGEcwxJilxlSNSj2oIT2zqpjdIiZAbj+Pr89fluriBdATbu0gBjJNBMUzRvc8Rsy7E
qD1+k0uOx3ZDQWSzFnc/ilKjWxxkxF5/FNrHCaxGhd3pKtGVpRbcD6sxZgNVg6KjNgsMcy/RIxkA
eSpln9icFDgWipzDsgYZFFOOKIIZPovGQtJRAe2MPqNQy1ZvYvBRb8DlB9C1rKkcTtkYtb61A4bx
SpawjfyGxmVfdXYpHv8NDTy65DN8cIokasgnqD0CtOwWB25AHgxT65m32j4YrbdzV/+klUde2D6P
7SsbcuOEx27rdIZC4Jguk1ZX7n3lchzHoN04UABNH5aGg7X8wi7USLUjTZuwtItieWzMDzOS58Ic
b1asaurZQqtVkVZqfH08frXzTh0ZjI9uGZ8MWrsA/1D0Epx6sEUadYj6lKK5GiWwxyAHtoIpVRNn
0CXQZgiDaiwaQiqzV5CIasOuX6lT1ghs1+K5hVHpxY/ictOGyum8MnVQam2tEHBAOuys7bwdFFii
C5R96bb0LrQ41/ebvZuWMkX2x6q5iAKUr7eDIliRIR/hFaPdnQw0Yw9HJHz+HwIgJm7C1DLY//ku
wMurHOf4YeB9U/toc9Nj945x0lSOcYNLtq99FOW+t9hMIOBZkwDg3JQ0VF+Wji9G0r0N3R6+Z2O9
dRy7AZ+9qVyAzoSWRE6UlsMhPDUJ4hyYzYPHlA3cARsg+2wizk97x+i2IjFFCx4FTSwc80t6yFgw
Tu5nnyowM+zhGUb+Gh3Q9xe5myAZouUj2c+eu6nVSuEMh+VOd6q3TDLpYLaWsLt7inyt4EDU1FJC
fG7kE0Yd5szNrYaGYj42/Cl33Q4TxvYcjWF7dVo6K2YZVFpJKpnVwjqQCgclwcxFeXq+VbdayIQ6
Kq9BLWmrsK9vu5CzOzLICz/WWAgNStmIn7M7qzq/oTEuOVTSMZuT9ljGDokApozpHckVfSzYEMQw
qWGplOmBChXp9BFiGlTcAUYkl+mhov2j8l45NwpyJkssaltIO9R0PUK0oXxYN3zWZTBhVD7OMd/g
4sLubnY6M2kuW9IID9MB4xXjk1vLARJBiDcxDnUORW8eFRA+guTLUgtL7aVlqaS9Yt+2+TtTSiiw
NikYjtz2Fa2vfOdTK99zVGIFOD60H31LvBYmbJcaxnPMlpvFItnicifvP6vbUwFGIFpGrSnf4UTe
GomBKsAK4nOFYShNwNLEEKeb9s4LBj/J0S82O+chTIVke1VRJE4MBFTghqEhDr5ZSmNiZYuGNiqZ
DZCobIfKLavwJyPMMkdYK/ndMuaIMLJZ92YB5HnEzUceHybFvOUjsD6HyRGTIZH3ezxNGogCVJ1z
j0lqb3XjjLHo6Q/URNaDYWujDkrPsNOF7L0NfpORvNbIvOpImLHolvxWdOW1Yt2Qw4o2clP6sV8o
xJcrjldoJCJecen4ztBgFNjRALYOABV+cliAeKtHrK3K+/YVzvE6N00rpoIJj46u52ZoYNDzrEOU
M+BpUS3bXT0zm5zVOPRYkOlBLR591XLeiRnqwg1GAr+923rjfGfGgm+DgYkYT31cFVpec/bbnPvi
IEXgX2QsdogQdKW9+MugCISdgnh27ul2jBdgPgTqRK05hBdFjdJkwSM4L85BLonXf4pI1luMVpE/
UH6uS3XLA05rhqKm3/OUeUNu8qwbkYIPwaScWrMO2il7eE4hD6jiefREV+7KztUkK8lj1zYN61DS
no83WKjKkT0+RgAWVHXHF3gAVM+6jC9brYAms63I1YN2mk8BCKqKcASZIwqjg4zbQFm1ATKj7Z4b
e0df4xWW2VpGpNLwPBVfFYhNfc3fwzZVrxRPN/rVba3kKeABLYC4anZHvW1J0RamCeWlRprinHoo
5z6OSejqDiP5DEFT67EPFy/Kocr5SL2OhF3FMNobLp5GOMmmJl9xIkEREBYK7d0dberTpYptmCM8
tkrPRnqoCt9zRY0LoHQV7NAgr2Pj9DbH0fSttFCbVMn4d4/ul37JWnSnAdHX/PGmMn/yhA8sEq8F
yajbbbVtztx4X7tLu62HgHZN5LRp1A51g/eDvZ2XBwLJUdCdV9eJ41Y6plSkz4JgMr2NjTQBU6Qg
Sn1ZmocTx85M6supML6Q2yj7nJiK4pdqQoQOoiugXBo2WTqLftE/twVkScN1rh0H8KcCLovbLACi
GUunpc/145uyLh0U0Gi9+TzLEgId64acFfBIVF/zsP4tOXJKBwVNyhcLNZK/k92Tkm2CrSWuCUA9
H8eN/lnidZ0WNXQmSAMYN+Vk940dhkikxdS8ZEo1mSVGPQf0sz2bJVqQ6IWIohXOYAJEJ8sp+yM6
uNuJSyF5xkOdfBaJKTNVyBxPMXcUY0iHVNUjO+X9JdvhNQO/EivyUMexP00b0KWeiswdiv0RJVgX
WzsFSOODvK0sQCeCFp2KSlqa+BN5zR5DNdC6Y7Mfj7LK6slQ68OfuF1mQOE8OPmMgG6KAzK5Uw8x
AqleXb76TuUh2i+0xNKVlnXVa7YFv3Lq5moXOi3o04P3LGhxjGsVKFhj8ROnZftejZ1qug8bpNxh
msU+/TJUbZMStt6hZiKlLjOMnHkZDg62uhCOJN47MJ0KFaQQB0m3Aox8Rm+SlnTiz8lfP5wYz1oz
GwPouOzNz8a+bVeMlmwWIc9zUhQO9FDdPJcM7ugoaKkamte0e9DcTOHsy1YOaa81TwoQMmrUNMzO
hDhIKO2AGg22AJE8Awr+iSK3IM9zrmh9vSF4ZwiaXAHAmzNcnFge1K7NR1z+a/N5aQlFkOBofIL7
uGmUqdPiamKlH8HXSHnWBhf6TC1Qrtu9GB/EaLN+zmPRl+BsK3tNZgaYyZQgAWI3MBGbRJtck/32
qajlfCIS2PNRlJKw1Gr9R/Jr2S17J1lY/hNVgScqU7jOT0Cdy4sROiJbN8oorVB6Y80OyO1uzezK
Gv9NmQ4TFou4OLtu77ukg62vIbpYy8bIkEUTvXJPSjWzJP+fUyWfoqIki1qW6kcB9+Km76uQDubY
5P1PLyeKaNOYCfD6xzMoZCa/i7yVYW0xjiNb/mPa7EscDtqYX2JCkZNvaa5kbwAOctwaOjxRxcsU
F34Rq+vsxWvsAi0w4XLcuCWj3R8iMGf7yBNVKlYHSs7V4uHzJUtZLdUwPhqPNt9tusfYr9SENMB3
25u55IvidSDQGH5xk4S4wAe2nc6jMvS5z8nMb6mnAw2677zDY9CPN1Yu4Lc+sPttpCgHVCe9ye15
knuwgdwylXBR8+kX+7mU9uBFqCQ0ME8b+sMsv+PFi01Gzs8its/NRyO8byqSJECup9ucR2PaPotr
tJyC094CwzLl9UN2Gf3sd7KgYF5b6iNxhU6Ht6i8oD8w0eYsKm7L3H/THDMpEOIqnNogJTvpLpdx
4T/pGiIuGsfll1NuzJvUvlRJ0Z04gVVYpeXij2WS0wen/t/tYSuLsAcTcgDrjblunhRabocpPPqJ
UkKUrttzd/yaBWv2p38AcOBIbljjiNjDku6KgSWKjA3McrCIFZ1sm+s5kXkKXazfTx+jue1LCg+G
BB37nGrEFCXdPQc6SjnkVLxTgnyvZtgdm8qabJZwidocm4OCoGQYhv0iZIFsRFShdzAC132cUupg
laYv/PZIxiqeo8z8oG0D/QxGEEKUV0ovwe4KQPQrsRs4KhAYYZMbx3MhFJDOo1L63dyyYkPcMfpl
Sg0/lXehKnaQveFb9RZ5ej8ZrU4PPtuLgzyQe94zr3Iv7ydxGxh6J6qniXN33TqmBE9yt9r6DFZu
ObqhN83p8HVKLKIfqzQQxsah0LKhB3W4Dx7asWE4u62Y92XX2PuJpnWuYStwrA7kosSxyymJLBjF
9tRFo+s++YUCSBDOFel70LJrnud5w/zu7euUQxofXXKWo3TBebxN84+Aw75JbY3NnjDlWHlaXGWt
ncnCGEcak1/zAduWFvnMyJngT1Sz2Z8bQ7B5ehd1TjfP+L/hZW9u/KlOwNbW576n2RV+x61FuGkt
00RPQdh5p0Q+GIV+rvKvNe4Yz9IoSoMRjOr5r5gM8UCi/ajC5+KWsftAvTSQssjrBK6v+/H1zzW5
KeuG8qohTUDf+AqKSB+gz3JqXAGF+s7lcNBr4VVwlyAw6jzyDLUCCmPkim/TYgItbUsEPaT/hapz
9cT8fw+niiXemFJRyUhyW9pCz66HfJaYkyptOWdDdtJm6AF+rCWIQohyXgiGN9uthhvhTTDeX/nn
M/SMtdqVaga0QCp6QyHMv5SGszR7r79rlqBe3Qxk4xd/NAfu1IperHSqqxOUL1PT0LKxII2apvzn
P7Oux/sg0r59eSWFNdMtKuqDSKwd6DWO6TT7sJrbIqNbwTDcfzmRbWpbwRklA45oJIY57aj+dEMf
st/Yu8wnQjnJFx5dcVDgb7Xzm1o3KehaBFku08ip6RzTYS+7SSq89oIV9fXgHhjHcYVJ6SuRicXI
36htR7x0xGBclQhOLS8kHflWPMJL3BMZcCQr/kYC+M9LHyViQ6bHdEVMqw5O74epQ7tdc/CPoelY
k1orgQfv8Xbg6/VqWf24M3GpclJQLrhsUL3ELUToo2CVS5bW7wshgkCcMXIxsFW1ITGFy1sXQvn/
ISEHErWCFsAsO6EwRS0pgnjh0fU7UeKpgFNqxKYXzfBnXUv5vjhyZhEbMe8o0ZWt3i2r1/Qm2krE
EMJRpcCjriBtI0ohRsfq3J9EKVs+ZbA=
`protect end_protected

