
	parameter			ORAMB =					512,
						ORAMU =					32,
						ORAML =					26,
						ORAMZ =					5

