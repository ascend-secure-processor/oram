
	parameter					IVEntropyWidth =	64,
	parameter					AESWidth      =	128