

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
clQ5mQP6ZK2BUdMhHPMZH2cI1zWfNuBJIPlb1plNuBJGBY2BrX2Eh9EHFkAHZloyrImm7TZHpKlk
BTkbjL3L4w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QNqPt9Iq3rNASjEAWrQpJIWqP1mfCAtEejDgBg5C4sS/yQGQedbuvSUT+uWUtKzddjE/dej2wni7
1xUvI5j8Whxhd1b7WAhp0Jij8NAEarv/P5JzYI5ZsIA/AlbYuP3s8VWemLt7lN3XgD6u6jXpmFKP
UH9BrKE8AY3H9cg4Qcw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XrFMccHORpxZnZgoluicML2HmWGsQakT89kviQJ16SRBA7IcNIf9kiAj0vfWjBRoyQiy+o9AzIDR
LwbkzRyzrWW0zZbhzWXvlmuyTbFrKmGxoqRHqfWfR/rPzGTxq035uMVJyUlsZGVrBhcqBecI101n
z4FGIjwpZYJfC2DuhGjfRwxT7ZJ/UyV6jYAJqGIGTvohZodK+Y5X0tMJ6QjhXRJzGaMGsfXxVrfL
Q2g/2Ptni7AjGWzBUxBJ4cGfgBVF9UPcmsMMC2a1Ll7gOSQ0tesprflenm4OZOiZkavvfr/TSPmL
rAcg/GEA+zY53Xoo/zt08ZjD0MZQ0EmYki4+Ug==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RGdZQmpjWLsG6mE9MTa9Eis4KX7tnw/iM7Zo70ckZTtIQTOYwZ4yzFZKA7IhbfSuCjATnrxrbbUJ
FclVPCReiKsiVz+RKuypKf/OAvQ/TSdyWffieqepOUYqFy6flDRn38322Xxqj+DKh8uB8bXJpEQ0
CMkb72TKR7y9ahjNfGI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nq6UOYsJERbzojA1Ff3KnzkqLI/eDgzGxPCkUgVazp4gdSK/8xG0lPUbuaQ/jzsWKY5MvP7/7mYG
Azcwo1ATzhAAfKtvwzUK8s2eBtQSsNb2y9M09iGTW8Dv+WiaUaxgMLcEe9IR1yaV/TqS7IOPuK72
/2GpEdQOKAnXiKcwFjNjsnVsfgy+TT6Z0cWEYqVl5XjdCeGKoor059pPmKrkHQ/MfobzeA7M4tNx
aZc/yAMTYll8neLmdg6sfK4auBrsFn+76xViNBCGH96W/9YfYvcfaudl4a0uk96QR3K9p3p7LAH7
+CuTtYNquFE5Z9r63rjqm+WF4x39cAE+TfJnpQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11744)
`protect data_block
U/1tGQF/jhOs1qT/slMKAC9MlAV5SjomylJl7GcQlW2a3mtjU0ExwrBxeODIoNc55ApoS0pe/HWV
uD/aqmZhSthfjSUYzh9CRkvtYcj8GSBejTG6UclFZHaEnZ0yRVUL3ybAmR8a+Rs4O+BU6uo1DN0t
a24JWCHC4IM+642HK+Mc6p1GOyHz7wVt1NP6l1xCxOVUGPBorlYe9Tg6IAtazIh4hkBvGG0DvudS
kCTUitxc01Z7Oawm2QtrmHZaG7Gr9Z2KLP6yrG87cLo92IZgY/zIMjIjm0OCX9wxkhHhTO/aGNhT
jbiH3b9Bw98OCLP+DYigPXX+BhA5YIRyciF621XlcDz7KWYe4yq1Gn2D3obbCKATK89dpR0ArwLJ
Pim9gSxJzWzYdm0LRl+iHgf71+Feu1Bs0OPJKhUd+ToT1vWwBu4CAxOrkr4H9TLVq+RPqIweNPhM
C4BpfOfvWvp/lTVyHw1WkTQ3lm2WdibKErYfJ5Ckm68V9iKK1J58iiJIv11jlbpTEFbSfYC8kwa3
YntlKC3Z+BR+RPlCCFiBFMkiShZXzRI6ELYqAAAOA6hybh0eKR3S8Ebb7nfigRBkdyAOFTtvV+KV
foXHc2nezJ+1r+/AMaE261TJuVOZhpkMqODxy3Iw2oz6AnnpIxkwNW1H8m+Hn8vBu88USgTCfHSN
fg/rzXKIAJWSp+Vte3wnyG2KMetjyljKjF8cJxSqkk92oFmlLOIhh8tDjdQbIU1/SBzVu1T/4hco
T5CuvfXFXo23U+7p82H0EGbhzGqShEP2EcaM7mttwDJQsEtgW3H+N/JAP2gZIhdX3D6Q7NdUJSBX
VEMvOfrGeravVEr5kguYJSc2bTyL08FlcVfg72CliIaJh6o3qlG+4LDjr2RhFNJSH9VHcvrZviE0
5nbMgdBOMh5TMMPTDO8t2nMrkmW3U/lIC1A61bEFb6NEu94KAEnRYJbU3+wxDTnXV2sojRNBuhcD
Jf3be2MGv3g6IyFUS/6eIczVpeR2EG5CmkG5QpeigUdxfG1fF/x94ue3i1pnYu5na+f1EGGlPtok
aXKBJBXfeHGSk4IiKhupcrkOfv4PTg1kreHn8R4ahgjtTCwu9oEj4Xk+fYIHRaYL3K9K8pqhAnvR
WKrzzT3o1x8lxlcNDfP8gdSpDULegIFAb+D+X+0nZNbRG7zARFFpVJMEVL86nDefFyktMWwwo5X6
FdE0dIIrxjO0CpFLHFsz6OWyzOi0riwAwYGGlD8lSb3kftvO54RsIXJESydZUHG8UbFyQKjBqDmj
mPjuVFTCj4zjZS7naTqdksYXgFcZed1QVDQyao241EbMoZXRN6xCFbKU+8r9Ha0cas39NgBbexKV
5SXsN+0FpEgudzBfU3PBwo75HnVu9+9N0Wy3WEy67u/JNxbyaej/iZZG85cW6a6L/eVFs5DKibUn
qXL43OOTsLTDhmw4H+rViT2rhBG6x9ENG9sy5JQMUIMk2eppR0+6hVWJngHpR48HwiVLDYrpOgb1
DbAbfmaqJDPcmcZugnlnbEZ6k3h7bs3XzxAsYpKn0y7qeKOjo9mpkMmSChGZGHoZjlSEnZMzH8LZ
IzaF7GA1lWDNY3VaXI4RZGzuwwwIDa1GgMX/2arLz8JTXewyIg30L1XZQ765hXdYgm1q1wyzs7sy
iK9EUs3LEhSbeiOI99Ql8OZdThTG6CfE32btyKmtXpG25wEc6CozKZ5MeZ/WWlecD8XNFhsnx7oj
g0fKdjnZRLuYDwI/N4FfrrKye/TMvkK6wE7HbbxsNXN3uWG0zYf9uB7rZE9yZ9dkJJNFANh0kz2z
v4TRxvK6CpJBnkdWUqXH3TctJdJgs82uFpZp1NwViIA5oqqLPiUwIduranNH+TEW74kaug0vm8vE
knL58fl6vC52qPb27tSrJmnDPeexG9ofRwiAkzZiUHo6e9gp7CD/8Fv0vFCLkzjM6CAsTcFDkUD7
53TCQa5yJjt7yPLBUdMMgNvM/kWHzIdJqtuecBAYVK3InKoIQyOCoceQ9guahxr4auCHpIzWdNy6
TPGwKHtgjDs3Z/+5hFWWtfUp3NYo6rTqknq63laZzHhlD3jsf76UZQ9foO0JmFZK4lNqo8Oo29oQ
levTs6UE91D0VsCuyDFwnPh5eiBLgzJU7fKswxI3tJKZmZ4/lkwbpOT6hslKg2yjCZHGWk/xWSEQ
/TDLEW+uMVmipvarda1lWsZLI7j+1gPGu3e5Ps+YuWhaejfxn8BRyMV9crc94rVahPBrT1b1SwC1
KCQjuA8Lq3U6OsX+2FVI2/Ko9eUbf+no6INYXoxlS7+W872BsV7QLhQBbc6CpRyNyn1vuqbeKY6Q
WOrINrkNfu/ZDCjcT9zqySaBE7pdW772v97noyZXQcqnLRF/W40B6v9f6IKbR7lwix7yx1oEIxSH
yaDLyXpiM6LtOgaiOdjY8aQph83NZ6r0eM8YTod8ishZ/NU4aNwkF8flHCjMPls0GKiq0XKvJHBq
sknTOcXnunrJsxBHLA2CamusM82Ms4i4ZG5TKKjesKC7RZl4HQ/tSR5owXwGX4Bh2Uo9yd5GQj56
DqDHkXbNZWQd9+OcdUcuhZ1P1zCamUyH1gOk8HZ9cGfSFgm3SGSwuzAEP/yZNJWB8PTqIYGe+kv2
B4eyGuh4kfbi1wdUssrjy4NDGdsP/u4Ry6z6LtvxH1MGFdkCeoLEQ+CpybmFXkEaaQ90gpjgKRfD
lV98m7HPM93L06qT6I6FvBMBQdUbNzpEPb3h4F2M/OIRIK5P/CPKHWzLtqZy9Qm2jyoqPoE0JRU/
8B0HACNsZ4KhSfJoQcvJdN4iCeItji5geylG4iRblQdqoKmOgir+n8UOPHFYZmlj684oWRQB1IqH
Fe3wzvHZK+02sJLv0BJfi4y+YE00YDxeuAbn6wyNJX5pDDtKGCb8XAleTbFaPu9WbADw/+GDnEdb
wL2ODOnHSZA3acC7aciVw0WjE2z4dBBtuG6eiUU2ma8gdOWOomY8NX7X13Wp3qaIB/UT8j/1x4cX
pJVhCrouFE2wt5aBZ5SQA7iEIFkMFCsJHJpUcYpj7XmmQ8WNV/OlPusRssjOuVrMEaWcy9oouPtE
Hddra8tbgWU3QE0RfWeuPjcup6NkEBBNxPj1RiKYGhboa88sPpzLhByz4iK5JA8rEcwHE900ScIb
n5XLnIDzkrIX0Oqlw1h8MgFyGw3C+Q3F44Ctdyh5C4sSEFRfBFNgRASfS1P9rzeZO05o/8iY5w1q
GAoXx209575YT9Rfgn9j5iV28syQmQ5BrA+Z9TfW2ZCkfk4Ot13l/1CcP/Zrcyj5WLeez7qlFtuG
h8jSUzdVPCPvzZRvM3OpfflF2fCljqBrwc/g/+ONRiO/ppzFoyfgA4Uyw9X6LNkwuSpYV026pfhz
k7JTy6VWxemER4LhfnR11iJvenYhuN7x0CfuNGJHR2Bvek1kEnc1pJQCDwIa3YLCkzTSOPXargCv
QPo04OaqFLuxtIitzzYZifwLQAyJ6m4t9t9Usf4rc6YN4uvGmBrYmAuaY1INuO5RIWaGhYZuecUS
413MY4mbx8hc3lCHzn/3kgADfJpXmTkf/B7fkPWi+T6w/Rid8BOgvz/TCPFCakXAG4PUNHERvySD
Aee5LVjcPcJVXeuys2kJ+2Fj8ngzhR1JI0dnAAUOyR5AypoxJ6h0CS3LAy6W0nfzEPh1Nr++NRzt
R7+467IarNcEuewqiqvqT6RcSriqfQBIJPm3o7UDIc72K7MRrOEfKJN0wMjTtEo6I9A6cdxmoVW6
mAyowOLrBzfrDH3WIu3U/NOsCjRW8YyVaGrS5ozscCce+LrECKGVyfyhSKCwXz9vHUwbvBSOGYrK
0F1+lQmfrfEG3Cn4cZvJb5UZUt9mMuYEh2F4XieNTJiw51H3WNvBfatjr7124NKeZdShhyQFSCdt
jQy7OCrmIw6wr5vhmiS+lh5I4LD/enZRXIBU9zmUI8nfR3tUM0VlD8O4z0tQ6g6k0XL/CK/06cXD
6zXdScbmTyGj6NzFbovq09xWRs3kzybVDWVsiQVvRVf+0VI3R56m5HtvDyKm/m8+nBcylE9PWL3+
L0d8uH37z05wXNJazhZqc6NjfNQ/4wV1IiQr06qaYSwIXwWgBOCjzno9J0KR8wdx1dPYKDpv4Gzc
7do5ggbsyRTaie0vmBcuWBCNNK9ZiX75hqBPMigAKWvt9EKC33Baj1Aks/oW952Vhi3AQWikc4Zs
93isFfkLoP8jJxIr7bcUV/bs//m1Eblz80GDM6haGKIJ+ePB5LG7WUAJ/IibKyf6MdHsDJb54aLY
0SxcUZulivb8CiS7sCRrGF6StTOQJQkxEoDFBY4ICu6ZfkybV+E1seFiEI5MW1NzFElrqgTRhyiB
oZN9Gzwvs+6gMK0J+ugaIS8hr6JJ8sX8hOSCWlL+cevsvXVVvs20faUiJeb6pjMYjElMAs/C3c0i
nL8ew+nZzsBDcLESVpRbIVQcoeF5EG3WbVNzbGn2o7GiROIsy8RUTPFiDBSSScmW0gUIkfLYm3XY
QXSzwV2kHxQwVM73H9yL8M1eKj0RCPFEApMNMWk14HWRs8HxnNTK68eUvS4DkDDXkuj/Z7y8r8uX
Mwh2Dpb3ioHgkgPEZ7H2mbpLepoSX+LargxFZFm4TeE64nbAtprcQ1sIerx6VaiUpqsvxsUmJyQy
aarv6Il+7VXIJ7aWfygchQb9D8auKZ8jiTl+4Lkc2dGQyiNgydidHb5doz7oKae/6x1C7jt70uxn
Bj48nAb5uEpMdvXVpGR7CFli3q76vI8SHQbrGaqKvRuONYAUe+NC0D6hoKsmqqC9eQcjGkFKoWZH
pfMvww1Qh98K4pPA9ur7tcH6ETTWHU+2zSnZ8oKgqqRh8kqpWPuZ16DGA8c3dUMa1hOijBIZBNy2
+a/GcoDQkuL9LFC8lOzxXEeGO46N30BSP4c+iUZGO2/GMQ0XG+V+OqpZuBI5l/Oz57ZhFsafIEfR
qxhle+ILB2uTYtX7ZKRVh1kdeF8tlzVcxetFC3Otvj1Ujl8WcBxg6BCPJRku37ARRHSxmUzuvRr3
6yuXl3b88RnLCBfbmCwc3wL3YuVra9YVbo1+MRaa6kjuYq8V6jI0nO0sz6JmwsxXQaV/Jl3AAZm+
/qWZrgO4d/7+48vimSS3NsqcWEhQmzWGwrJoRqN7MWU4//YzfM0IO/zxey9F/HlL3lrjTV5WP725
HkEvjD8FOwrNGznGl5YiX7mhNlAHWTOhMeTk8KmcPnM9jnmPHHHs7sluFfVn+CUmhkTPWJsNYIRD
8BLXfRbZkFkarSu/sYkUudhwhZkWsS74cSLPps9bHa2dC21LGaNIA/3tuMd9g7dnHggEutjWMA4F
MVDaadExyVLFh0diEwbEqE1UPSeVjKRwKgZ7dcBCyKxKEOn2DIDMjIg7WjcKXpEPZX0be7jyAjWM
NwZ51SSm7P1jN8nDk8bfIiLoasRLJUaDYFBDDVN/qjIC8Me9KC+bI/SDcxpOYRnOfwjNFXeyZ13L
welsTQ6nmcLG6NmtjbliITy+nqzpB3otkvGBIkC7ZdnC4+Vojs4dbX+0XOAPLX+OH0Fq3WZlsBCR
qUHzIt3Wzy3rhkvPI+KWafslVlkINFx482CONoBepD14PtGLjABXeBwFnejsmWkwdWym9rECV7iz
0zGIlzg4txTxakymbFAgtpbwo1cXRGNq+HxdLKvNdWOBsXTdgomErpNo4rZArmraVjxACr0Ckzw1
722uHlaItA/PX2V80onMH+WrcDlYnL8l1OuJN/5zrp4hpS4zB72pByhMiBfY5iNXqAxxF5rEZkg6
DKtxsCmK+imALtGpBL1ofFP4el+AekQeNtF4BEJB9Q7UIf109fh6qHLDmO5OzQW51SdRt9GufWKj
DcqmK+XRKqwyV8MKEF6BTGhLvpAHN1OlqnTpv1X1rW7sDPfimbxQhr/3lM8UUirRZ4xA0ariUNyJ
+kXU8b5K6GhQOb3P8GLDOoZxph3E66coC4NCJnqZE9VbcqGRk9ysNT4+ngpTGgpoVg/iGNhuwUvU
1CGX197+faRG1yGFDcBSuC2ohz5BirhexaoAMGLn6MQcvyPrS4Lc/i3qGXJyKRuQoyU4ttbMbTiz
fG2RHh5npJLTe75bjmcNJMO/OW6ybpM3XFc6o+neXgy0j3CnwPoZ/FT415q8Y2Y/73Y8yIvsClUG
AXCgVMuwIa/II+VoU8g2rMcgozSsj6NaNOHNrucyWfCXS8dtab55fmWJ4ojvLSW+KgkCc/0xITWo
XyiXUcbW1lkOf63nuA7qqm5KMbjJGbz+i4CXxnExbB9dU3wr5VfHqFCqNQrWRjyQRumqaXeKNE+B
LNhO/jJGg+WyJORXgRCbMU9nEr3hcaNSKjsSBachlh/74T15pjLmPAqgSbbl5LDQy7BLfPBWVU70
AlBR+rnDCYhMkiBF7PenY4d/GWwFLlJVY5I0mIKEStNxbkWQdgwEZ7fO3uT7TS1Q75A7xxXUGjoO
WHd76epxu1LWui1yTHEdFwuLG3TVH5iOoPZtX+q7np1k9+CGQkbTs5VExRQshfdmTRtSeEdF52yw
KbPamwDiNaG1oc74NuV26DYyqFseY8Q5GnHvMjMgQdF7mzmZSxxJuifQwUSBG871UHFP8EHZVvO3
vxLj0MRS59RMdHi/nhVb3RmGxt/UvNcSr+PWMqQ3donj7c5DLlBMes+W6S706T8VPsMjoMuUcqvs
FoAQ2s8O6g5cn8OAZDPoqUkg4f1FGYy+oAyI1F2zhzMpYwDUEI5+vK1BPhdN3z4kNQqv9lCmPc1g
iuDBJYhhKScUQvapVLLYjjGHpB15C95GUZWbyXn4RG+8e9KF74HzH0V5wKYL1W9uqxN8EWIEXHHu
AZ8eea7Optg6zIITX74zCR3XRNxtCXadfJ2bPgKySRYKgvCjPqgdGOAcCE9t2QUKPBs//D0Q77h1
vG6oPf/vWxJqghU0Uqm8v2HYWOao8CBoQF54Bt8R21jpvKkbQFDOXqRTE5zP8r0n/CxABHskkS7Z
7T0TvJIqDcjRBPcR39QupC9XZz1cb/0hL2IvgXQVskwLCuOcvhRigj9rtbC5ybi0qRx98jRdgncC
ic+QgmmE7ErmgCpNptUn5diA+b0pSoz5S0+rg4FY4sqLECCecqONl4+a48R1yg4CrAn7JqOVDDuq
vQWr/AfBipIod22fkUIwEEGA/lWoYwsKvPcwkfWXko8FZhOljYCtKA26/ZAJlZz/4VwhI6sZQla3
4fRrssIDw4z6psHHAk1ZQ4QAF8eo5f3PVaneCd/glYGEe/iCSnXUwFvUH1TzJnP7o4JemInLZuPt
94WPwFk39SVZkVb4jPQoBQEgtJOO5gSMPIvmi+AzhZs1mmwPkLTVkf/JKcuk/BNEKHmTiTucEJTg
3yKdDDnIbTqmG4lgEcHeqLh53mxzP05z/VdPZzv+ju7gSGaqZZM6HuQl9My6doQzi93Ubfg4UNpU
Tw7z/WvPhKctLSZtdoqiOwxNFtWghB/Wt4Q2m19zoRLOa7H5Tkeb8y0szXxr41Kq9P4gxGJAmmL1
fUjAzgVNQbhCB+o5NQs+UBdItQF2ZnbjoeDUv4uuNMevyNCE4JWiEzoTrJNSMT61k55pCJtjGqV1
6YGv7OJBforjQjJBTT9f8AwePItVvQkPNTE5mKsPCIiW7toCWXIJRX0zA+r4WZRNQALdSJ/LFYB3
dwZiBNc3ZXfiCsowmpBALKmYjQCJzOh/1VX0HsmxPyukPUvX9D7yCeC8r9hI6r0GrPXdUkyvE69I
Pv6g8qTX7OGHXWZcQjShroCYDahM2bReHvDNerYo2FgaFhIFQ2vvcdk42r7ccnn6JY7bKllMNjWJ
GZ+j81qqpu3fVXm97muMlOVeyydDFDH4A+aTTIsIQa4U3TLl5kIcpUD6Vh3kaH4168uFylIIygOl
+NkSB5GTUJYqAVzV9tWIzEtQT2wbQf65LLl3axoj5QQ4Yr7+/LNP/0ngdJgZJ0hts0hLYv/c1sO9
ktsOVwee0VWNzIAdRwAcCDOJL0OGI1GkH0eDZeyTHr/obm6R0yFiBzVO11ekWqviKJNW/sZITP8s
rPqFCAeic9RXICUZuZ2yyrsfRQzGdfa2iV4aWmN3Y+/L9Mv3qHuUC1P1zmFTSSA+cRJIgQ9oDgv8
SY9m2zxHjv13T0ijmE28tE9siApSADLV+qJ2nxUUmfDtSJK0nCmguYAvgQVVEPGyVcowkKYnmyBR
MUmDJE2YtVDBmDJ2ZFKm/J0VOBhhYIL8KXQRjHx+ZEibdgiii1F0w7qS3lM8YKMc3pGXX5aIImmk
NNyp7KMdyo1k0nR3/nr7rRvI/s1aNlgpF3jy0E8cRfF25xVYv4bkZBpRL5+bAZgU6lZcdgvsRCkt
FycwpAh2AsKw3NebirG7BXzsfTM4J4BFyPpKB1Egi4VnHwTOWffHD66xaXSnflGdDbyQDVhDF/y5
/MC01pHiD7F3qDEnVl992M5NDYRvPZbTrcMKV1anx6Epktb3MaYzw9EvNgzTZnp7bW85Dm57M+il
koikp66HTdu9JJZ3YzPq/mSkCWxn9wLQ3CeGSty/KDBLnMHT/hDmNqADzNVXwugk2zKvApgMJHlE
cZ25d6ZhuRO6ggw90VDtuH1yMFOjbB95iWUn2iGtg4GG3jbMzMsRV8cyAhuB7QBqjPGXp9ScjotY
Ex126j31nlAfyy+UQXdscY6qEfFh7NRbhsLBVEK0zpNspzNFpGE8fuLOs89RqPb46/6xUsoHrqER
ZwY+zalZTkCb3UIzQJGH6Jfzc6M/X8euXPIYmRek8FNAxjFN9tPuyhsj1T0zbp9J1NZHJUlyb+rl
ZYSGySrvVYFZcvXkW1ZbMPs6r7RtfizvZCZZfF6VKSGQnJrJ6MaS6JP6ckUoNJUpkZR6zWnKqCKV
vk1ldBiqE+kdqhOcsrMoyllwjpdsxIv+FZTylZ+ieBxCmN1D9S9oM94JLBarjWYu1r96ZORUPo9I
d9tQLeMy096yyGF8Cqiw3gSSP673+xkqTp44YUFJXqyhckp4th/s5bswK684kjj+PR7jB3KuMq/D
qmdP/vcw1y279Om0G7VsZZoK4LF6FXPGA0IuW1+8HHBVRhJBsbRChCFyrM3+ar697xIm/N5LTGOz
yiV2ynzTYluCPSarp1QU0rfiyz9KdO0cdUVI8HV1acXrTqP1veR0L/8rkXL+iw+05+vJ4a0w0mkG
XzSaB2np7AF/P3/tLz7a4IMGX0FeKCh8thRGC69r9S58A3pPs2s0RVxlpE9DEqAbFR96dyEhheiI
nxxN/EdAL11SHqPncjK24ipivjU91Or0awkFY/JM21b+I6NONl2e9dXxSWgVmPR2+jrDtjdX8VK9
qouqh3WoyUjvMxmr5uaqQI65mhlzXiZ1Tg8q+tkCdJe4tKVJFJp5gMxN+atUfFNCvxjoBPx7dRbD
jtx2jPPHun3IbM2oBLLAQ4+bWUJmawNAF5TG8A3/GC3Fksn85PNjiP2R9mkMW+GBjW4Uq5RoTKZd
zQYqSJuYcJypUhF/R/q9Tfb1NN4i9mbO6r7R5QQAo9jixBi3LSTIECj/JhZ+6kGdrvmqVbOuESoz
ZTE0AMkaTT5s9xDqoBX6dUOF36OFiWDaOu7DFsGDqykCnzZx28i23OmCuRBXrFmpt3mqulqGBFiy
0ZvYwAl9jUJa6AzdypZ5lWxJFsf8oDlB7rwxo6JwbGaHJ/lxsko4nC/aTURLcJLK0tZ/+KuAIYy6
ZthjplLgoolbbvpHqwgcyFVx1Qmfw8n3Rljpe8TCV+Ny6syl/oLNvIImw4zKdUQi048PHLdu9KDp
V4o7Rz+0PjAdb999g7qSKW/ovnlRhpdx91s2ncYL7BjMKq7M1O3fCRMkkDo8xR2b5MhQ9Syozjti
LSewtn+I4uzIbHNJw5O6Va6582siTp7BMoWhQYJZfZ+bJuSXRRDxf0klp7DHJSf47La/VQ+ILSJY
YJH+/EXR33NZG1FPtEPIeLDjviYrNsKcu+bs/+023aJToaVMGcapdgWb3iaJb98fepqgj9Gp0xcV
IZXv77wTsGAImU71NvGOV4to9zRs8E+9XrK5WaS/V+pyky7ArfICJzD8ri503NmOL6KmWEnMHXf2
pivrG1VtRc+iXc3DkKB6jb925FYuww3AQYDxgQu13y6k9IFGTtXswXWHamB8yXhtlxhP3vVPL6aC
JML2cNjk5v65miww79C2mol7kqjPAtVlDp0tycrZhq5OCggzXqN/9nCms8TFuBinOfm9fGIWxBPg
yS1/Q6eyn7MmrEbD2wDygE8Bx1MKkW4RfaLyBnSNTeaJx6jHWGSGrOR5zkZgVhn1GiwZJUp1uNlF
/oNhHE7xP+KOpm2fxMlOytvtUT6Bf3xVWBBycu6Em/86WLXvxB1C/teTfjtHNCAJUbZuaUqctu70
CvOKw/RQ8a5tORAKt/DRj4h2/nTIeqj0trH4Xnsztzs9QLD8P4ZTNXQmtF4xsiNbju5r5p4rZgRI
Qod23vmjujNj3NnPrBcIZb1ETkNVV1kRZP1Z4R9njBjIC9loTo7c7SWXcozLWKhnlm2DM+8sQKXd
iKN9fw7RUY17F+vttqtd+WUOpPsxJ4RKrLVSatKFL4i+8rk/0panXuCLBtjlT6FLT2KcXxrF9SGc
UMTXmrbg/IIh8eOlCEnr0Lby2nNRjrzKKKw15nzChDGqts9QwU95Y4vAQm3G5QGSW3CopYCmhc/8
+/KooeFjBi3+jk714mpJPboND5fENB6bTfwbHg2BA55FAGdD9wfLKtRP8AeA3QCEaYJIkFp+6vnh
zhGgVDW1axEXrufsl4ZKOdGPHtv01TtgaDYx66zClqYJDZF790cr1yvN08u/OTrDTE98O78abyuV
SAnuZfsyJMhEVH6W5fJ13JRKsoJ4pVP/uDdeyGlSjkYid7V8gZJ0UEicSDTaTeu9UDNyXn0PCEQC
tqxCJZIpERKng8wJ24fLv5j8CsmpCfObMMAhsshcvhdr6Ap7ioy0QmMqQ/7vHl4P6+sHiP1uYa1s
1W3P2Fitmz+uDsSIjNIBlceygkIfWql4fuq2pMvWm+JDTw4/yBFWApmGd+wONAbfOjRkW+Q8Ybk3
xssJxpPZDDi6g8r7IQ9b7QEJLlaORQjxIWcL7Rwvp/cCs7/eW7gWWlHX2Lg/lOkbQtzQ8nuGErSa
JnAUfWdlY7dpuIjZSpyrOhSTqpjSfR5oHUw5YJqO40xa1gpFYjtZYsp/t5r2HhIQKMaSr19qDCeV
X2rx2TfrJJrSZ9FpZQ348SPVaYlSCO9vwQawCUP6MzVb+/4HalFhXI2H37AEYnU2O2mEzMoKelGH
nKzcrEX2KaxWd8SIFBMH/Em/ZlJYV999R/iRnK3L+rIxrYKS9atbtnKsNECwnkYCUkjSMPCr1M6j
jkR5CxINkj6BX6UeJpk1zjt+H5ByzxSMJI2SX5QX7kyC5LK12uM7ssTXNzm17GFVNnP5+bndLxPN
w402r4S7YDfqG3c7bPvEib69O+0A/4PxUdD9cnR1h2l+MhqE1LAOCdKukElHo152CsKNij/ocgiZ
E9dKszWucJQiuGfErKlPZj4f51ddDGyqi1NEANqIj6deQyGDYZ4XuMHU4Tk/eBsfeWv580U9bHS+
EtpkZNhzb5Rs2qo9+/T6T+H+guXTe/Xyq2gcNmGWCUpRb2aOT6lmUSXmt2xKz0A1bksm9uIowpMu
QNxBo1tkNzdZ//XaVRHHEXDbr5xC/yPabUcWnqB0eNR6vjvIczT/pRX2T/BZjY4LdhgWE29lA/n4
VsMRN/MUGynzsgornV8Zy6x63N1W0J4SI50lv3Nk9C6x9qM7YDvJM0rRG+q1vtLNfOZO9h2qtR/a
SmT6VU3RsdXJJFv20Y9fjx1NGTH9WSac1D2JoBX5ZDLE/LC5OhykK78II7M//SYR9giwxwq6QZRh
+RcuayO511LsY8ANgeyGeh7Jo/BOK+uz3Mcg9GFCo4P/UaYZ7lPemU3Xy7/AvbR4vqr9P1x+sc2S
XZFA2bx48x5YY+lgMTllNAoLup9cdBj7cEKuEwss8MwqslBY4nbJl7XzD6pAlVfsTViL8ztNUzFB
9vvTGc8j8+oXVasr/bBdLK8JdfMTAroZdq97/L+eGbzfsEtlCm9YKMF0uD0Q2/U6LGDtOroPDWnr
kQ6g6Eote3IEEd9Pzbx2k9IEY6d2wFH7F4ZZOqfB9NE3QJC5L2vLYGOjuZL7b5ci2TkYJp8PiNbk
0JBrvdpewUeOxNKi1bDcynF/oYKwVka9SPX/Pp4TvoaBEGvnIJiLcwGeg37biTM8jyeeROu+9CfM
N8SA867C7J0w3VW9o0EzesEpXGzxRo+Km+OB8Zw6kjbpobNSPldt3P5PstueYrxvIaxLF4+OlADM
hPX1kxy5OXa3bKjRVVHpGYTn8s6xeL+Afjt0y1HkaqJDLk5ZnG8e/S8ckrAVc7JJyZyYzV8pUWl5
TkZONL5c/MK91BWpiswuavYuGlwORag7wb8YuUe5BhlB3DEgJE9muf7zC1wgFhrZrxmETcxtNsCI
8GWInGE2OiI7tUioBbxmaVVgFAXKsMyg4TvKWmi16XzPDWTzBrCkRcl6O6f5Q8+4Un3oGAQsbL0h
oCbAScztAAYeezorbl5l3wzVzyJHS3eYo6jWdhKnCFOn9AEEsDAN6bA3pfklIrzmN/9lImcWh6Po
lLiqhl9AXooMVBEeDWqF32buBA36yAlBy3GW3xo0j5ubjNzMjVSQ05aZgGdSLKUkgf04myjNZlTs
mqVT+qxtBJuB60ZWuYltPLl8LntFGjTaF58n37FcQxwuvyfswFImrP3C4aUV3DQToxbgl15zaUZL
3fdNEDOBA0hRnm/ZieGJQJGc/zHfbY9HkrtLKeS+6DfiIf3hLU5/+HDgNzq1W3no9eLSKBLYgBaJ
0g63bnLcFAO69YMeFR3RO8FDfzkWcJutsbvVgSvxxe8eEq7JjNRVdkEQ3HHE8A6bft43DOC4bQKD
ZkZ7t+/Ky3O2FH2c1turv2sqgXEVeqN8La1R2BuBTRFSn4SXBkTpPDpwXWesth9T1zyFaIu/i2I3
N6cRY/vOejsK1Pk0fWeVPZ1bR5pb4O+Bvua9M0RM3MpdZCY0IqoTRhST1p4O/7wQ2jX77ePOFyrx
3Cx209KkbLbGZQBRtFRORHuV7VxZGHHXe8GFtEZLK3w5FxkCTPBvJIx5TKZCcybaLmmD60nMxIFt
oo2TUpMQ3hThCAklyNhtpifKMeL9J2Y+O/SDSQILrvkCM9Xn/Ce5hpuCAy0B78drxppu68k/unzD
1cVwhuoXGaPWZq2YyMT4Xqte7Hc3wkrqL/geqMqLMDn8gGlbIIfBHA65s6lZ8PUYDbKswODVN1/b
W9F++kxp/AH1Glbb5ZRn98dp6YpxPph5aDCr0pLWaMfns+4w518tiBPeIwVbkpY3gssAkrF0d46H
1VJC5856s5En5WHW4TLXi8K5QhAa5On3XxZ7rmXX2tZ3VAv3pZByN4l7aGNkIgkur0oUtn2pXoAs
Fpbf87W4kUHinndzN1u+ZN+FCdRE4Dybov57tkIeL+lt41NxiLZV/TLdZvsJLGLpuhTjQCBuynnz
4w6i2sRkabQRsl/UznabBxuzfdwb6xoDfQu4Lbd39ut6KXtWnOQxjIOEUUC1ex1rXYmdWBJ15Oxm
P/3Q0FOBKWwstFtMm5j0XXx2A2sG4yL/YWzOXqF6mDC1mworJjewdpNu8Xc1Qb+3Rza4Y7wiMjHq
BZoSp2nLsYEHkNbpBYL68bWtQO8WEmw8AxLIKIc+noVYOIjikcasm2LuVDfCe0DenVBKBPsOd3r1
3BoBftCCbefNAOHvuShQPUftFkooD786DhDlSte4DWvp4q+cIr7GSl9dVOvj7sqd+3PdJS4nXXcX
YpWZOe5NzldM2s4RI0OdajhO7iZrSl5R9bwlrjJqSfwGF1JouKKySjYyp0xW3jsT6l00Ef+TaiSZ
HWIxwklbP51dv014RfV5VNpwG1TkjagLTtCj7VJ8S1uZkCDwJ06h+Y5Xhap1Jk+x7QWytfSuZPjN
97rAR5Z46wfTDpSqiDuwK/zeuITfN4rKojQoutBmCfWgfLy89YHp38iBY83+VqYhBrtpvYG+FUTi
KzuVJKlT7PSSwnCR9esPrLik1z4ICzLMEjSxS78u+BimqUFcy7FCghCtH1rXLdJW0baLtm6LWUzj
xfeHc3StxBETygpvByvYyJLNe0QGpEtprGEzNBh7l9qQfIKWxhWKcHRLEd77Y1Yg0/R6LLB1HIix
IvM7quSJpLcTiQflY9D8iWXsrkaBwdTI5qBJmaLmy4f6waKvTkpdXBI10de7A43AvDtCaVBqbO4j
ecTFDAAzBQ0jG4IyFS92ttWWzs09UPOkGvhd0S6RgbG1eAvlDwNAHD9Y9IzFxf2Mpd9b/O9aWnPZ
Ue7TBokwnwyUhCbyabpEsBUj1kFFFUC9hXgitob+7WShkpVxVL/mevNkrnSk3kkNJzgIiirbW7Xr
wR57Ir30NBkDs3MU2smU0a89hWrysksebDJu9yB2wEt2Qpd5L4MVO4reUYfysiISM8J1hXp6DoD9
3VQ+q3/nxSO8bM0SuJtUUhJRzAgEueGtNE4po9LTLIXrL5+NxoZ+caDZTKA4EKqKjY04HLBTn+2q
Ms/n5ROvYKyfmRYUfhnJU7zmbrxQtLDURvS//CRsPZwAWyhkjC1hmPiu+sE16MhOtxHwEp84itH9
kUZYgmG6ESeV3Kj9pSEeQQlzmj8VziZW2oJWDnSbzZEoKR6keT2iOXPEuIZnTV55EeJanAdgLamR
5Wlk75abe4lv8IKyPgNFD9VKIa+L4jA9upiJGtf+JupkEXQ9MgAWERmsYmDFdyvrnK58HbR1ng4l
nHgY7B7KgD2HJ0zGicyQG6tDX19hQbt4DQlyvGo0EOTMfXiruTL2enUTe2LNF+0FgoPd8p7mG5sb
zF/CFb+8rTsbUtRcXPzxf2Dn1unWYlUUzVPL/zmmAZMTr6GoYcOygjdLGP1XE8/bnzcnDcOj4xJr
Dh6j8kuyxC9OLsF0zZjGWyOtnKjNyBdQCrIaMJcF9TkJI+PsCID/D7ZOY8f4dgKzxTLwI+tM1nlU
uODZydUWsaeHTH3a1e4vpJZSu2vwTjvxrj3eZdm7mACbDPx0r62LStk9mFOl/7deAy5yy8biUDEY
+BzszVztCdmjOdoU8qv8pISlTjIpQ78uMqc05iQMphufXwRH7P52r6mJIJrle/Sh7mFuqCu/v4GT
hKEvxjcf7VDGa/ovNDfzYJ3AKyyznpKYVfDDeMC0Fw2jo42qAj3qPlohS+2BHhkbo8yGhNOLRRTi
01yx3cqDJcotTA4YoabuezYzTazBrhGNk5OmyXcjCoa6+k7/oiXA+SwWJGrlD2v4vaENpCyHL5f5
/w9aYeKf6kPCOW1H3OR1n7yFfOcYR3d0aB2Jp3YBwa+tritTesUsbeJvViUSJQw+nY5ppce2Hx+l
fevI2XKL+v+uDYBRxLJ1lYrZWA/4PyRoIG/o4P3sbhUEuz8lFPbAjt26pL7nX8qrTHjAKOP2HsND
Idc=
`protect end_protected

