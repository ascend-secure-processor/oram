

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NKBA/jFNZlBNolObnhgZSN2glxkea5aYh6Oo8fQjSGUHdU9GhW+6qyv5320jK/wYO9oAjt65aMRm
b4KUTlNnCQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OIkv8IIW4TfZ/RAQLjTLJjF4suwR39gvZuffY9zX/a40DVy1dx744Lt0n4QOUxWtBv+ddQv7bWRu
Gi9JKYUUzmGhqHpepWZhcTCuyRZaCKURcjuOftviPAtjt4RSuDhRHO117K4ELJ955V1UtftzoWPm
FC19h/BIc5UlO24EgEc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ioUk/EUJKwhbASDvqIN/oRQm61ru0fNEPgQq9oe4qPeeXJlhC5lz8+wNSGa6jqeduGFs6tdBWJNy
nhrriGkIBQG7T+xQzJHCHMGRfKnEt1sKc6QiwZ4wvJhdXVTvq0NT+1r3JgZ1d4DJpO9xIXGEOMcu
i4bS/7C4CndxGT6mytHc+AHLCMkmPpnOk9pGF9DzfMDG1f0dITimGjR05GMpjFaqQd0YQy6zJ2y5
WChnoXQkQGv0eQs+IaI9Y/SgE6i/me3ONEuKRKdTP7xisrDg2ZiCsebODtxnNaXNdVE8oNIlp2Xz
aRSNEVHqapKMDyoV2FylzwF5UABaV2Si5Jhe5Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iKgXaImcxRij4BKGfHvzCeK9lCz7PAHUoI9MLOm/LQCVJg8z1EqBc1tE/pxakoTW8hCYofeX809v
tuN5vfsOBvFeqxpuY9q+0Z2OgwIxl70gTOZiH14PvIOfDkNAP0KDSx9K5KAbcjr4muWrKIzgZ2ze
qGjUcLHoNdg6ll+76ec=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KzN2sDexjIxvhNejON1nSxkoQviWQJdwsVejqI0DrWt5PNAJyZ0jQlJXGDSlVcor2DKbESCTzeC6
2W3yrAkFEUMbAOtWXgYTfzerK0AxGfZE1vY1cb1uD2LtmxgpdMB2dqTPeSLXTKv8mIRSj8YpH4Di
X6t2TCoDNcRgwQIW67UrTcO2zOSIRnnAGbnUHluhm8ta/tfeSvDb1CKnyv3FPWP7Xd0A2/ilzKKS
bhkYi9oJjGTRYubl5ALRrhLKkCNLABVB50lRxd6P4Uwu5igzMJ7n8Z87V2UTBOLae9vjUbxNqAiV
ISknxH9ZFocY0ZsKp1U4TjLP0oc8XqpRivSUOQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14272)
`protect data_block
mJtArJ+eQjnDQM9x47pl37DZJSDOGIxmC463LRGUtie01VrQNWsU1t2BaaIHcX6oiyckHKRjT+Vc
YWIbfW4HYanI8wPgDJnaSaJ6/ERtraGe6dQ0AS7ZKkdTL6MBr7xMlEWEnPuhSe7xkmag6UIi/sQX
OiE1mDKX69/wceX4sFJzhNYDxgZjXbHiZjFeIqBunmgX2bGdhVWvZ52MYmum1vV094Iuze7sNOv6
4jcpMUy1ADq6yMgczfBtRHktjnxmIzbwtEXwPC/DbiAQH+18s0bQyU9NzCxqWE/QROp/VTo1XoO0
3atwd6iv6dDzoT2YlnCKArKj4xnExHJ8jDYcpnIPydoGQh8vloNiGA4gIf3D88gf8jEv+4os8p1p
nQWtwndNv/EB+L4OUjvvbqTuNfksWqDzBJiXaul2ZAvIvqUDCy8dht5ci6Z67m4nNm2LFtbi9X0H
PoXMcaXW/4Ys+B62++/bawEwRFHiNaC/MMQUUNhUQy/+Sdy7+LPXS3Aez5DxiBw/UdVMaBuSrTkT
whybZ9qvCNUb1/fBeDP0sOpsMHuZiLmyRsCf+R0vw20rp8YiB9z4wlJwaqkv0RVcB7UQOlgzxQF0
cQxcDnYm8fKWzi5701uCV2aitz6zTWFAHqR8JyOiZpWnl4rmfpTnEmaMInOK0ddA8d1U818QZGOD
1sAQTBkdDIIizFDDAZTnhYGTUraoBn+XtX56FCbSTIlhiWjZJAxstHT/jjl9T0SRaDQt/520ZwZq
sNcrEMUJ9ERwipHg8z+1l0qzzKS+ynu9KTm1ObbhfGyunPjdLSYMIn0H0jbVjfr+ItdYhZbNUr3h
+4kg9jt/jMUlTG7D00ka49QPN35OZktXz0V93RogH4XnJyOLCRCoBbTVCf1JEdK1clh2F7N5HkVU
qjZ84AMCGOavaz8Qk++iUBBjNmW5Egqw4TxzE8QCzMXY9+y0MmEks9eMezb6UByOeIDAHcqC7D12
+QEvmlOITFEgRRrMZTBgm9dHtPMUFuul6m3qaQ52JvRO6a5KmLTszpTl4Y0j8xx+h1WnLoJcKxCF
ZL7nuQg/+bXBZYBiKPabtNFHFB3o4guhwLVk0/Sfn3wkhGrfJF+v6MDeO414EgV3anZvPioRuHTz
0NJWuVhw0u7bC9nUpg5zm74hzrMxwFkWCOVZ+jOy32YXTlKfxk4oBMUrhjUH2dNzzheIvWC/tBRh
67EY1Vzx93c+NBGTkLsyDw85xPmVistFfDim4m7GvopIPZU9S0+0HhlWYgO+GwK5gcw9btA1N45O
T/X6A/spA//oWKGmhDbYsjHsT40l55U5wgQHS0l1NaRQz3YoaizaddNyKHjkwkaVukMAMFg9GMTn
97LkW/HjLp50G6XmRO5eaa2Lht1epUT4OigAM3ioxVgsjKIsm3V/d+tKcwJpRCKwbJfD5BZ3ujGW
P5D2fEolKp+ldnTY4zq76qhN1UU9K0m/uPPoJi5P9WRisitqIRslstSrG5YT4ylsOvKQ5FXsnAv3
K+x/Vi/3gqzpUK/AwP08LoicIgf/8bB2S7pU+9WQbB9R5uALS7xZagaBow6BdJ4L/pv2yALrbSJu
KGMpmuoReef6ALHsbt5oxJHZNfxSxZatmCBxUdb9cps5c1RDdJY00BRmxOLkKRs4BJwfC69Rox7L
AFrcKXVRCH+6xVUvRcvu+oBDUloy7NwR8nNAoz02iZtFCMJBs/owOmfhpyJ4oHaxtRr0DBt0MZp/
el+z3jrYumMIhFCBSj4mam9w4t2rNx6YXCu214YOb8ilh+XFbOuAOLKRw7TPOGfrk3iPP+R3mU7m
hQDKJXm2fpoqiRNcto2Z6HbSKidNMzxp8b4W+ppE6mKOv7wSaCxtQkrtPJpKoLbx0/Pyb7ggr/jd
2+ONx30NQVLsoQ8P1EOw/YcDfCRQ37dxt2KWLC9BoMWKshsA49KA8AZMoeGbADPkqWjTTkdWh4on
XYOYV41ol1U6Z9Jf+gK86Ln77qHMvGU1GkX4LyuTzUhTKr1rZ0fjkqBhONKhGDbmqDA64m/4fS55
hVsph6TZAqfQB6ZuBcCwLDkp15150z36Ok9ZhdJ1y4CVnR920o9n+/a9/rLVmRsrLlywlWA+BtDB
RNzzqgjq7oq5mzFaHkCQKtSjHAulPVbQC1MytCxCe3QNxDaqoLVmcvB50yxRQgZjh+WKiyiuQTPP
qv9PYJfW2DEuKceTBuewv5ECF8LsRvaULnZoEoKYp33J5cCbhAIWFBk6WU05jh1I2xjugrBHDh7+
CJMYEuO8/GnOwS3Q7QcOkGvKYgbx/wJxa/1O5N7cFhegHSiqLY/vxILN2onpRrorRHB1o6iTyfIZ
5NMdYdsiEb/cKnEWJlGe8fcQAsbX6TyjlP4ORwwUSjJxQWgaQH5qH++csKhDHxRjGr/KrjvHuf+9
MX0F9EnKk5W+ZG+6SV0QGnFGBI+ylRkqNEGtNlu9m/UnOy0hgWEhZ3AM9Qr64ILu4pNaXyje5X0J
sZCPRUJefrLOj/MLI3atUUipr3EoKt+ATLzTKjnP+MKFio+fyKfnDPVzHPSGdbX614338GRFR3z/
PsKIMybdZf0+TcOQOp0BwEwJc67/2ClI1xeODDEiJQW5wdPfzgekQPfaqhJP+0RsvCxHb0E6+LUO
uK7sXmczOwSbK0qgKpPUgMwhebbOHebhau0F5Oh7XxfTLEAkobGXqdDTE3HRqGTNlWZyWBJHL553
vCjqmrtsw/FExjrPPPJDVG6XcziurPTveT3j1CcrKZiserkYyvURTla3CYlcBQ9iLPThPrOxUdOX
NPYxzqIV4GSH3hflKFlTmHL0GD0dk/L+YIhpFzUQFUH3QXomVt+RdEoHpMQAUmYpuuGnU+JDn5dm
16oyQcWxi45ctxnpu8JfOxpXgQa785nZVAlfuEhWod4Kr09ydhLqRGzoUE7kt5bNh07HfeuLxDc/
BcjwBd8msp40L/WpgP4dlXtg/nsaCtXXs5hAjsEsPgisJOCF9htEEOG2sEg8vHiL0ob4tp2zUvAa
U4kEYe4mn/ZWezN1ax/etJ3E6X1jwFIBjpVYBkSIo5vYgQFmA9A3s5P8/6xOkavnoxTvSLZ8GcmG
rTDKeHp9W+owNnkn5sGsneQPWUMmvdWi+Mj1tIkIEpT2K+TlvzZC6Ha+ANpvjqvGkC6UnuXmJzMC
XVZSYS6ANdK8yi+TM/goxMoSRRwS30Ybb3Q0pvmR6Xipq5NBMgW0W6hlVe44tW1SKCGg/SV4OGnN
7jxCbErGx8vWXkY9NkYDIKN4VRtMSifljMfBjF9fI3jz4G1rx6N3f2+1NGcGyhl7xruUXSa0sLlG
I7rikM+25G1EbeMD8CS+tu1F03rGt+W3XIeo/i3ayWA2CsAU1l1f0D8k5iOvhKXg1Z8Dp1uZpurd
RSicFYJ55RQ9HQ1GvvuwakpBGn1WmL7wDdtKFjL+damt1bCxbLzZYLg4MUCJd93UfszggYUlYESq
aE2Q2t8yPFcQuLA7hDd5oBwRLFUEsHvLuAS86WzsLLFYSUyNmGA2TJQfnaaSYFFPEbkCq8QQDuln
h7eyTbOgsZX5oW3knXFElRV5HU+2rqFOBltpmMAe2bKl5R424IUDd/Vpq2RYLe7z1u7U3CzCAwvn
HCz+fvvEyvMcDl3wOUnutrvrOG7HtxKVl8MFljQabwNAQZU2e+viO15Dx8fkfkhGzTOIollqllPP
FjEJoX7pu3W2x+APZvWdV0dy4epY3rp8EW/oqkGjVCrolXWsDNK4yPTPL1jsjvDSxPm/TvbTlP8r
lbvIeJr/QdrlgK4qf1GjuMJNsmw0Oue6xnC+DGsntSseCy2aeFxkyB0M8BAjrR7j6anH7TCXsRYe
mD6aOmH9gztwKvV/F/btAwbTc23R+6Y4rXHBmBs+51vvfhrrK8as8EBm8oUPaR1++AEULdk+M0+X
pI+sIwjYg7Ca6+nR8GIUgbn8enZZZiVZp0LLcK31cFVhd06sY7Rp4yRdgkR7YdU1TMGCcUzodu/u
o6hgeYIKRh3LLDUh7b0P9c95sff4WJCnY4UfMP5M4KdJmP1ZIUTHx7UL40n3Jv0aD4NX9QWpP1BV
E/mBmBBdzEUfPNe6NZ43vHei2HeG3SFiAc4xtxyTsheM/XjY+6GYoLe7QtAuPVCf/b96+n2GFAk8
xO00yUVE1ydAgbdNdW+WctmnvFyHplH5R27rRGpB5hy35ZHoVTu0jteHrOiMnGnfyOgcIQtR0APm
7zhJw+bWjGIsS+W0ncWCMl5r+HbsIJS1Szmy6sTs3qvHgBwdbd0FGnT/h11S6Kp34Q8rBUioP3HE
ey3rV2vRzfshYIQ8un17i4nQMEU485Ke+nE376UKML7zkOxjzbdZl05ElM2LfNZxYEiV798T2aGn
ZWh9J78uLfI5tvAtjSpmZxnSjaRwlRiSwxw+DvpJ2RY2wDn6KpG88zKrMy2NvN4UZ24QBnYyASxF
OeSYkXxbtI4YJ+FEf+nxbokCFQviXLgHCvZr/M7q4Tmje8zhaz6DKy//iRhTwp10FMmHehvPpDQ0
LzKpVuS2kj9VTp96wTDIXRIRyFfQqg7WmFYU/PWvqbm2OSNPH1/IM8Jn8D+Lx+WvlQKDTL5I3bzi
5ytN0wwRPwyNrx9TROynV1zT9Tc7ZOOw4Ah0ERgsGBrXezHvADIfTCr56DJVSnb0RTYfvqO/nsMR
dfvQrWRofizv6jj+2rYjCC9bG54ODZmPuJYuC9rq0Go4x0tLj2mMj+iH5K9JDL3tgJQj2S1wRKeb
9z3hDignxOdcew+nML3Cc+Makr/U4gkp3OIYUr8sfuvu4ny+Qn359lxvtvm+Dw1cbj/vJZedixhx
TEZ/1FBAw/NvRFd5Y1SPlohaMXsyq3IrbwHx0cSEHd4MRR6rcbVYGLWVTM4+yZ6Co2uYaHE/DuBy
9QUMQ2ArleoESOZqT8J/VCzjv8wQvyX+2BeSC7nbM4aUMweQcdaN4SgHesU5it8dc1CyCti7lmif
HNRotKqCi3N5X1bJ4sxmH9ujlazRNnvDC+dCN8Ib0WuEUVv53ZP6v1r++Qf+w+9u7G/BITPJ0Kv1
74Z/Jm7KB45CvpFC6mdP06zfeFuDA0QLgLtlTLoTCymlQ947Gf38nGXA1Bv4SlwNyj6+uNLgCN+N
0Utohr4qHFXoNAkZ/aPfbd5zYJc/1u34GZsWK6wnhSjJ4fVv2nXSebRx85pVuGarsMG+2qnZwUbu
I6Bh3C/XvzNXLrCCt511YlK6Oi0AN/YAi6vKq8VAsSbAzant/iNIPsk7V/WAM8+d0ltRqETH5zzD
LEPDzDXUwjHGfT5C1byw6nBGo9sGz3xODUGFr9Rwc37zpVEOXCTdst+i0Ti/PYYgRYyma00Y/Cfg
lSH3bTSslUYhJivNzEYoxjc8EN2RouNTKqMnYU3YCNnLgwas6uo4q4axafjMzqWmwkav8wC0A1hD
A/mq/wrmlK9gKRIGyB0Rwpap+vo8BSNYJJt5xMh61AEr3dxCnRNqS8rWCc1oQenAV/uIC+ZLFxAj
mA/+ZTLf7LRjM2FoU8QHRiI7491JIe73Le6fXgzRjMupwTkHFQOacUdAMfvphQs8QROqQkrOnHa7
Cy4GWPuo6EifS7iT38ZfeQ30Nvd7OIQPXMzQyGJaxHb42O8drNF93jCNACIi94TQ//JM1WETJTgV
oCuG7R8adCqiJwjdHae5R/N4JUXu/G49qQ3gLVdSsOzDrKzpvfuqWXZF+u7ueiZKLhgdyg+mT9Rf
o8Z1I6D0+mpkT3YVkdNFH6Zvnxp3PoaAzmHbwr9WiBn/v+97FInDA5t3QA3LZwTbUNonoQdKQPyX
p0y12EHX7jnQ2hAxzDN0JHdTB8qesaDvc+xsLbPQy7RZPk6Y6Qhjs6nDM8anTaEZsf1hImHTTRM5
sGtZ1+rfn2/07x+wkbkWH59c1KlsD16dmNHlEzAIQXwk4K//COrxi9ftVdoZqjcr8TN5cOCx7xd8
R4GMXkpaCPmloj5WVarpbCNGnOvcQmniZhFSJFCugpiNGhCGXvw8ERelG9kpx7zFwhaEUgn3dlMl
rNHj0J4qw7LHS6smK79nmlGqWaLfSVPmNEb2RFgbuwtlHdUQXH10llveDrx8ANoPoMZ2PBMV+/Hg
uUlMMim1ycWGNR9iZ5Gz6XFbKWeYInDyqE4URcfB9Hld5U9qtg5lmDOqFhOWz6pQUFHI2vqDtMbZ
SZNt+itZk7kt0vOxObLu4YDKHwr2kQ1enzaldRBIgPoPHf4e4XBVw7zMM5vVXp4OWPq1rF8KF0rn
6C3eT2ZpFPAONlI5U7QrHvrfI73Jrvly+DrCm8vm/a0J0Z3GSPfXQh6YCTqCy5EzgBy2ujoVNtl7
BLRNrDu2lFVQeCA4SrBUCF+spmn0e4oTw9O2863LMga7s1nv/wTiErDmv3+k5ZHV6ReXBqOhCJdD
a1ZKldP28ELQMFESXMGhtgAFy1kPy8ehdFCpFo8ubvytKp6L6lA/2+7MsJ70CrJ71cVHhXK0rF36
Z2GAxu+ayacqFRDDrO5nW+0njawN3+1oJoE/5V54Fphd1Gn6HjqfQmadNd5Sp9Jr8kJ1aeaZrpDb
Z+t4VAz/+MFFkNUWzfzx2kXEI/ZYq7DN8ISS1vimXFhoK5jcU8qf1skeIrn3B/YCLsjRXdu8DthU
gj4JTXk6sDdUq3Jek9E2reDWXH31yLjoiIMiblhpdYHw3X+vQWv2MCWy9Jqb7Kp2ZZTNSC2hkEc7
G41Ki2W19IrleJCYNzR67jQ4DfAzfiTueOVcQo/cOWkQ+x44GBC6q+CzD1Q5imYY8F+AMWxPEIYI
RU2LA/UVFz4GDDooEn2HLoD11wLEpB8yX0iQ6FvzpMQ48K/XN2gz1LZ3Nb4JY291EPPPkmjoOVdT
ujtXAaBmy0cNxNRpAp3HZztpuxPhv/LOY367e3h8ry8nNiMy7s9+Qdz63MjQjsLndCImcmfirYiX
qoBCE6HXZrjTXm84UO8lI2Wk7HG8CzRKOl9mNguNvqm8BvZ0JK7ztbChc8jUhfqpBbgJqvwZwNn0
etFoF7iVs6C9UPbvBgtXQxOZk55nUx2D/1ShApbs773xB/dcrkRlBv4eyFAvtkHwQuljUIRCBfDE
zOOmFuzTNSsEZySc/CejA/kF38+c8iaHQLuPAkCNki0tWZPxEgpKbdzVdyaN3lxl0fMNHZUqnIZ4
gNb2xvN5cVGOa7IwLnyERLpBprwSameHH89Ue7R39Hwd5gQqFe2sRRaHAlxEZJZIACd0vxFfHOTC
p2FMgUihRaATRytjxTCCKQ1Mrzx4FJFwwXXgBxOHXSmBgGNT/i3QOlnjjiymSqhoM4qk0TxJjtuX
McIzYcu4U+X1BrZJuCCvSw1TvbthM30eOnvHyOSJuPWruncrfB5LauzZLZa02GgnLrBTNihrWbam
W2nWzx10GDO5jGEQXoLeGyllBHfBGVMf53t5W4OCJa/RhZwB17ZX8BaN+zQGQ3/xTk9vV4M1lb9J
W1AZ64ZT2R24NBYxRtK3x9ToyLTD4VUqSKzn+ZhH2GyZjd+Rw9xSf8ZKqCD7KXotDfpzD1Xlo9kP
YZ9HXbVN/GNmoevQEP8//0dufBmtKEJuXmRcJwtP/PsLiK7qVkGLh9QPhepzXA9TCGlYMuG15RU1
BFKV3fOy3OoSb0mFOqgNj7I6snyER1TlLdMrUnAwyE2+IbMYNNYxH20Y2i8ZZ0s6T+LSlVJNjcc+
xhstjEw8DvNnRnZAg3hRwSHMmnySFVwqKD5+pgyJMAucblGis/ce3IuNeJ5Ka7yEc/+95zOMur6d
1CjmSSZjPFev9mAEUm3LcCXmcKqejg9bkHtfYr0d8YlJRKC/xsRVBqTw+PPrkH6ek5sXIi8BDpcO
unxBVoavV4NJ/7tNzumNQVCQ1MQ2Y03Jiad0BPE5hSBw5QlLyvtHpEMqWM2ZpY1P8hXrjVh3dEy8
xnPHf3GYHYnqidb53Dsz6gazYYshKXVXGYzblvTfEn6BYYAjHTXoG4bp03kPf9vd3LDdtP9yQtV7
LJW86YYcnqcGBs8/w9TzrftPRr9ZcltZTfGlQvxP8B0TgIttvpDoyYwhDzvqXSdHpsUSt9QNDP+i
KLaxsjqbNoyPof9S5NHq11amAit10g0Dogl9sinQ9TEzjWlJdYRX0Q4F9MVFsnuj8mefYf4dXljl
ydSWFkYCqS1VHLoZHdoRM4Qin727VbpXvYytwHh2G5rFDeEyFqagsFRA1flcwPcHNLBjtsbbJ56O
GKw5L/nc7SUMsf8GToR5vnKBND9eXFWGFXDqFtcqc/HTD8w/JD8dvPtu4fYMeKopQ8oOBzcPD2J7
T6rXtCNOqxWumFA8bZuipHEw+y+QdwUtfLoFsz1DQNl0k30JNF7uc8+7Wu82wBssnnM0zv4xqEsH
SxeC/hcnSZ5VskbT+kSbG0MHQVIN6GLmPRRk8X6dTGdrz7eTn7JwspztkzM1E50m+WheaXl1qguW
VsuK/ZxarsQvB8xFYukpWcJKf+DcF3Ac4iwPrtHTIE0PN7ZjQrDG5YtywcDQ42iA1kOK2nlj2ka+
x98Yl1MldYclk0f7KkZiUrhTyroczR4n28kYvLIdyvIbpTjS4jjqYCWcQ0JNQENicdVumVZXnWBy
TShICB0VCwABVQjvKdXUlvFp58YRfXPFsMdHS74eXP9TSRAbZmN8oYxNbA0J6szEuEl2qKVcxofk
UtvLesfDT1pugK21HPqS1/dzkOFUSaLjAoWVACljBBgFWVek7gjm4iyEeU/Hra9rgITr4bWxPcL/
HbBHYeOXx+fA89i2E69/cX9xsf/z0xwX+Uu/rDb7RCSE3sFqfminhuU1QnI0FZnR1c+96FzCMg7o
TrBPhuA0tl+AR3X2Z3mtx94idtN0JL44eF5Ihxmm0wUTLDKcVWm84W2WsD5ALWRhDUe8o2V/4Rrh
3fHXY+9qF+VwW63B+i4NoouhXsbTE3zmxOURfxrAzTGXES+3LXo8yqvvz1YSnY+aTehvSF8Wsngn
1EIha4AYHTElWb3SJbISQQCvbD1j3pLfxrQDWVfTeqgRsDh2gzHswUac3ylOXsHU7dfX7VYqh+WO
WtpHb00obpfe4qRfa8Ub/GakumBoq454f3mWzEj3+ty3z6AHSw+gljdD/wC/fQZOwRJsf4PlVzG7
Z5/ppwOlUYpxDxCCW/ZBv9BWuepxATtxgfaB3zxVx7E9Ub1DM7QxGZ0edPaxMfC9qpYB8vrO3HGt
K1zBIQj8W9X49CoXKSAJwFc8bOV01vDgmRziZ1niUKhMls8qQNQ6Jnr5e6KUOFgVDeCYPjpO3Y0h
aBxKHT5UbPHN4Vo0GVhQIaYvS6dCneMG1AEhekbI3A4Vtok1RF2KhDQF2D2IfSPZ7EK5MRsOIBtb
FPd3IUz8HbVGhAw/X9GHFqjRX33WeCOO9pYYaMJ4axkaX3fjsVfEcfWzM9Fleo4sjdf399ycwD8L
BqEhL/y24pSC6S3eW01MeGh9i3l59ljT4FY7udnA12IX1pNmILLB3IPtPQyQGORvLq7sV6FZqaSb
MlZQ5kNcXv8wNJ8kdHr6q96/HmqtWqbT7FS3tzsMjTbI8N6sa0fkw8lt2McvAndz+8pGrTKgO/vB
ytFEoAQZBrMWsDqTpCM0Sb8QuKXQ8aw0IXU/mcNMr4np5T3aW630UHxLbRT7ZnrFYpD+lRXwqqfR
oLeEzTyMbsoywhOXBttHqtP/mh/NsGUA+Vx5rUkkLUH1ZZiU66ie9EdT/In/u8bhoSrq4gfAt4MF
MLMcVcjzRIeSrqjxkchOaoYDVcqBd2zTsomYR717T2jxLqRPzItQ2CB46d1LnPeeDET6+Slg2Wn7
tai67EagzFAl8hAgE9eRbmxVuZnDJUhFcwY1OBG6dEz9hnto1JHLJQ+wJMUd+GV5rW3A92F2aPPo
J1vb+HFGoYvhmOZGnaLqLG/6AlV6e/yRxkG9hfsNbPVTBiEeIg0UKAjjQN/McZIjRD+fvEDjpXFN
wwXtgw3lCQ81T6SlTVB0BZIYhrDMMtUEs72cpJWICvFCnoL4JAYZ8n6GyJBBmi45vsLsh5dQ22iI
rd92O9/Vrh5G14ydz24Nmm5EHFVPq7rFlN0i1WFJ4FO4x2QjNoLgjfAK5OFZAaPiEev72OZc/tyi
D2EIods2I7L3+WiTkT0PA/0kX5IeFKIgnyNQfBB6EPG9P2Fr1vkhw3ilaEFN1ihVG606U1KNCCtW
K7mz6QbrZom7McNLiF1nj4YYN5q3N+ewW2QD9Lmx+337gfATeMOVmNLNwsjeHY2PyDTdKBJvHWam
z/szmVT+QnOOifzC29M+qEaYJtTWESI21X1dwzrw+0MngFAObAAv1kW3ENpdXNmQrVvCrzaAF8Mw
LoSFOQdJs6RAncpcF97KJTFXedSK9+EX4VoQcmaELdEhNxUo5dBEI1fGTLTsdDz/4xCi0UIjQuCE
JzIHljgtZQtItYtaYuvi4whUm+JShsW1SH2f3Sel+xrCcf0PTVO+lNJSVgZsaYlATSurt9Ps3oRK
E+iWzLm5Cb3EFFYKvI2zwM+XARVDM6XgQmpaMGgS++vCezfRM55ae4BGnj1vPLT6ySTp77K7Uz85
3mP0oZzeMMXz4vQ942IYrYe+6EEyugKLpF92NlprWxHLM8elQefAHOSWUwrxPVQzFZvexf18+EUb
ZVMzgBa8fJ8aA7th1P2QEMUsgCEqYdw1x5CcFPGZMdF9ClyRBLf7O2MmYlVS8vuC6tdZzQqogcPz
w/zBEeaD0QYzny1qf+6K8Q/YiIS51g+eqLufZ/jMiS5eFQtRQ+L3JCvxUGaV3r4ajTe1YgjlzBwV
VDddlQwM8pGDV1bkOiLc3H67AXmE6G+3pZML4bX1g4zzYe6xMahm+yAOsDpsaNtGLVOjOQoX2S9k
o9y8KSTymHkWd5dhakRhGrWc/bTmgM9BRk8ds8jRODTUzK+6/jbR9rBX7VJw8crN0ALNAWgZorhC
YJBdXF84WJaZ5FPhWyqJbMBjPAmELNqwmSenbb780CDnPrZYMK6MPcJ+tylU5G4DZUH1zW2rWqCI
MRdI1D4cM/cxj3mfdsc69qCyRMW5vf+m6MH/uyJMqHPdMzCr2N8ZFlbmv8rC/bKEBH2glNAbYCdY
uS/UgUqmzWIzqliw2lgGMsWeOswsJEFG0F/prqIFKefHGP0jw4Rj3tD4zeyEvnzt9kJ9io0nlv+M
mEKtKxOoVZeN4lb2PzzbuW2fZlKI9WOxqFAvggL10dzb8O4lvf69G1JLL+/KqUJIzlR77/75wgKy
IO3QsDPWlZtrcR2A/6Gzo6W0dBIFQR3ZEupsPnP/uZggiP31oSQs4dl43kn9r3OtZRHCHelYoyP4
PCI16snuIoN+G11HbisFz4U8GEFXCOfNRPL17ZBQIXDQVrLClIkmW53BWyueHxaguU5nVejkxiJR
PkV9fF9USIMT5QUqR7hYHkeu93EPWvMLUkyrPFI2TVgVNLKyPnWYMmcIlEcUCgb1p6UPhPQAJEXY
nmsHehz5dzZ2j3OCwSgbYVJpZ3gM6nwKwyVBlqwbX1meWqYblYpGS+WkxSoqagtVtUCHVCoCUbBV
qZXcLCenfedxXrda0puSEShCsFv9gQUPP/Ph8wEEBqXGGqxSbjcB+sFjUHOGCPUclCyTXX+rBGI2
DN+WNyxgd+S4YKPIirTTdgqnpVnDop1gdl59ykN066jTvwOffi/j93Fm6gP8Lzf2RqvXgO5rzXdT
Fe7oN/2MMIirjAzzSEEiOx7l5zL9eDN0axYxn/gGnk5g9uQA/1lc7vqo/UFYLrXRcSoduRioV6Zo
1deQMOg5W+jSDfRGIW43dE2lhSEGv+VjRRYKvxy4T1AhuGovXvMROjSgdgbF+UIwIo1N0ibJL0N1
NVagVRfsf800cJrTR7cP/0MAZKlr664raCVGFBzaPOAVUp151u6QGg29V9vZREw/NZsLj8J/PcEv
DVswBjVdwYuYGC0yw1UDZe9BeGf0f0Y00dPWlh30Cqgajd6oDgsB6EfqNjMEqjdmU5AbH0nwl3xo
Hcb5EOQT+A2DegJ72hRAb5ImFAkcNAzv5D5u+2TZujQAn8YDlHPDNd0eMzMJ/eaTvvVQjO+cTeca
PH8vpodxE9REhY4T6Q9eVvdv6KncKyWG7ZZMQnRLwJElBhrY5WFCL2rL8dNOqJOTcxwXLq/heYXn
e1qpnhlFA6f55X9tci8fII8WVsN+aMeEytYoGvSHFfYE87eXz0W737I3+FYwQugGB+qRB5KbmxUM
dHcuba36/ZUEwQdyk1iZL+fGwI9DRGvknH+50KyOFgRBioi2F3mW2nDvq4W5da7jR7hXyqexupuB
WCalhyEUnlgM29P6aQExnPqO0fzJIoYIr1rJdqxR7C1rdOM83ZOfk+8zTx1VCt6md18xtwSPtJTU
Lnf+u5OjnpTwEwzYZjXFRPii3HHmYpy9cRtyLyZpa9eLeS4yzx8xjIwkY5gRxFhgbSB4c16Ef7zc
iLvR76rkMYl76g0dcMOTWGDP2QJflhELrN8egiz6YzbuFFL8avgiPSdZdURu2PVWR5ZiTtAStM3l
Ac3k+e3KVSdFcJIwekLNSUHgynM4wFh+V/ZmIpVduwMuEG6/5wlNbgx3L4DugklxeZEE7iSQDx00
U63ETtWi+3VxU3fQA5log2tXIoAwNsSUuEh2I4/qcAQPuoAUMm1PuKJUQGn3hR5PKpJPR1gVW1/c
G3dVYT12OtYTHDFeKAZd4t8h04gFERrA5nggWq84PzIwghXSxrZenXSYD/xkluMvJ6OApWE9XMZ3
Tsk1S2zqmuw7TrL5s4xm25fnBWwbrdqfGP/x0zctVHGvAB6wC3HpmNPevshZJxk/SeeTHqUCVm82
n0ONx65Y7uI4Bx0V16CeP4DZwNH+p9Wd8QQanha6GkBrqDaQktScGJjdOtExS5ZKjruB+gMhsu0Y
fFRJMigczcaVHxC+B7XAckqULZUTKl1L7yBBKADhWmWNW4oA3Lv8xIe7mTzj5JKKN9DlBjOybD8P
9NTEv+L/TLiOxS6VBJwcXysEucjAitz6Eg9LTbJHsk4PHv5kvgF6kznzrkr4MS3FzuSxbkNpSHBw
TAJmf7ZjB9mTQ8Z1vQVzuLs2dIM5nhRk/Wf65Vux1Fh4cfvHY1jA9W4Ey12vp1X7ni3RtZISMNAD
uupeXBoZLnYAD92Sv0XkUv3SLw8mAMKPTw25ylwvGc0y1VFHDNpR/0J3elSv2G67ZiSYu34PcrVD
pU9FXs9e9MzrzwNpG34lyfoWM46ZJKU68+QNRs/7/rlXdo8+NCIaE3Zr7xnj6SFdjwY+kBCBcxgn
Ix3Hc+g0x3ovO0mPS+CkhjGqf8xTczMN1qTEH5MfaMhSP+wyZDwdaDrD7ZKWun0keczET7jibEvd
wE/mUlMDcidUSaevcbOmBQcSPMij1nl8d1f/7540iEW3A95O799rOtDEqrU/qObtCn4S/WJL0E1b
z5snNqfW8yvSoLV/+YFi+OJ66E6grWEwCqcW5ricgffPCUg9Hq+CrqiPRSS4FpEIuw9No6xUStEN
5Qq4AsxzOfjflowBms6zM9WBU3vMW0wa4I6+7ujOHaWGfRS4nLnEliEiq2JHD+DWqs+N8bFJslIh
ueksGIJzoVb+/ZtQXcRavI9PJMqssfQm3yHpM28kl7dFloDyV/3KfGKDYkPxdtqnxDnurbTMFOPP
ZVkcNtvv583hP27M5XcBjJT7O0K1N3NiHS21ru9WJVCWZUCp9sAx14YKJQ7/f/aNkpIHQRTme1P+
ATnMn09hj/g5mrWgTUIM8PynOZEw5AoYyWaX+9FqRW/rLL5+Nh5VRIkiwd6EmHjn9xZVmIfs4vdj
FwyxMhR3Gm4VMhjl4KsF0lZMJiy7HzhGrWmGQ+NWWUSKyS3rtHh15z/F/sDQ1aZ59zFcmlJoPc9f
jlIX2aMPYCz9yvWEHF4oKSWPXgksgIk2wHHiBcWw43enh8loEyExJ7W+xplHCxffM1HLgf+mZMjz
1aJVAL4WrSBOO+wW0+1vLh/yubvgdJwsV1h7HYw4YNLFN6ls438t0OcPDP0TzZIMNE+Lz7C4d2zb
3oPkBlByZiDu/MvqI2oWDkXqGCjGs8TCehDtAmVvfQTkyQKvttULbQWUw+RXBWIpoiAR/YKZoR9n
A4CS2H9fS4obIKnS5O7lcNnYIyvWeT+oKfVW8HRV0wefC861xAb+IDbYqNJIXxUyPb6+KOjGCfkx
FZF7JCCQn4YMCq8WU3c+22sv8esLmghQ2FGHHhkg2eSl7Iov6gyTxRK4VBhD3foiCUuJOlKi5X+L
9syy5Gcqvg4TD5cWf+Cx72aeWZf0Vi088RqAotJx6wgxcs8/oerXL+a694oOPxcOJrJP8ddAmqqm
9HOAios7bpI/95x/alam6WdDVdFQ2786aNAzRHx5wSVWgtpQUFM9DJzIvl34sFHde285DCi6Z2sM
5RxOtfTpdP/K9OKhzW7yhvuFemempUQEzh5aTu9nLrb2Rfo/QGTmFmO/7PeEk1vIyrudpl4qVXyj
gp8kmMy3ZJDQ3SC3wXpS26syCIrbjNPsUTPK1txVgeGfjC56MFVpyj/Pgwi5p+V6LwK6tbF1/80P
0ZQXyKh3p8mNXD+cdB798t+V5vkCC7KRzT84QWfNDQLUbd6MIaVG/maZUnkEpunh4ND3vpmKprF+
J9+NogkBxgv0FzXg9u0OoMvEN8spw9XMqcPQeMmBwzlKg8i2zcY3eaLUkoEbV9F4jYMh9SZ/s57G
DmBGyvcLKktsv+q10df464bmEGIzmW68+0ofhFhzIL4OWoqVnDWnnebkwVvuAmKU0hvemBhJH3Kw
tAndV6p815ejp+CeujE3oHdWUMGsHAUBNIg+GHgnkz7l+EigxFvUQYLkFVulDJLTW/wPFKK3tWoj
muxOVDtusHVVXqF8eDhR27b7R7kYZELbN36ynN3UKxTOdYEaP3xTIOCYmcP3v+RKUIDbLA4A54RV
CiPBoDaKi5lrsploMvpXFpIwiDnRdkb7M+XYRrvwLpGSpAMmroq+TAaAYQKgJ74oIjtu1ie9Njzu
S0rNja+i1ZJC/Bo/eTZYbHVV0DnR3rkfBIeJYQeEOORYJbFVsbvlgjj7Ck1DMXDBdQ2d1UH4/kjW
V+/0Nnsbkzn717O93xaiyjuhmDnJyXFvz4EN/Bf5Oq266HFzkFFa6qFTi1uAGHfLUpu+pWMBr4kG
XtODNsUTdvy1ZjtrEFUMFp0dCzd+5Bl/TkTlNqjNO/Dnv0YZIqXGG4fM6IVIaYy9Pi+OM3R3C53E
LRnz7zLGwe6AhAnJWN9nJSTAcV1w3A06i14vE93FKPxABtFvgSfawJp64IjxffGahTOwkBn8SgM0
XTVeg3sahKkkc+P8em2hBJk4XXKb3FFUJulwtVXOg0MLx9DzFHFabJSHgOPQ842po2xpT0BrV30h
w+Mp4xRcvJ0BaazU9Dniwbk4TdHs2rc8FjXrvCy1b5+8hQG57H/vtTT+O1yRJIuUEpLAmJt2nVwz
hMLphJJ9XLWMNl/59TxchgZNUV2IYkP+nKSb0zeWoHw95Xb0T3eE+5jPlPCV2oh3a9PNCR2b1u1S
zaJRmTGmLY5nUd/W1q3zomvqfQys88ZKOR8gCyP5jTTeuQHfkLCmQyCc2m0W8dXczEilrujZsYeW
qiyrbaO4FPd1PeqIfJxUchzZC4pqeXZvuoskBPOjV/ie9y6mKKo9/KQptlLqO3n7Gn4iJsy8Q4Li
H5FZ24Co05BbxaQ3JAorN0YUpFlcadcZb7FMUEvjD+BbVBu7b71aDEfSz6UnvMlqpMy9jQYbCmul
kjAE3aeGpDrnuqMPiy1Rla96SV1eOaLzQ5GNI1ZfnH6UBKkwqk0OJ2/wtvrSdZ3uWYKQJl6496vT
VYDdrzVLjhrB6rnOZO6nuu2cuNdbybuW9o9Vvz4/fIaQs25X6j+OoagwAZaoCKMZTG1B1TCq5Vw+
ffMbAMo0wlZ580P67RnC/ykdY1tg2M9glqrDBtAdOEpPBkAn9olZyRgdwPu+5HJsz/QQFHFp+fuq
JmLzr+q+OSWBY2s6rZOLT/mBZ87wnGPD4oovkHGMiVHpL0zt/C06sboIBEo2V6RzrE6mPjSzjClG
5G5Z4PuB9k+4zr82aRllslFJnn3tHH1BeKYmpxJ6Kg3Ybvv5vU8xfTIl/OkumBAgSVI7lovMudEf
0y27oq6zNTOrTYoW9t73xgGdM93hi+yXqrzvI6j+gWa1tXUEn6TXhaYnp4KPCkewZ1WZD1+1+id5
E1GJf+bd3z0E8o4N/cfBYzQVy8VGeCUi5WmJELoB3YSTWBEdvvQCiUerBqzWwD861Ya8eAn68Uhj
UkzBCWyr071QuyA5pmfcazUBMeLk9Gnv25Qc0vgYpmO4/1B3RhGVi/gdKsUKsXDUJzax9jlPe3Sk
drKCy8hfGIyYuKY3epsIIW6NsADWNBKuhyYYYW9zJu8FEkZD7AbyPiEaQ63SQTVH5utNYmIRZUdb
gpN588O6OPIawbP4AegGNQEXNSkPuhiL3CsnlD1QMU5DDwZx6WW2gSMH5jSJEzcHduTK8oavKkvZ
9tZe4gjyg1YkTCTooxw8iCJchmWNsfMBb9JLQ4XKd3vbXYKm5SLanHuRsh64xPJbl/8LVxK9kL2t
FEkHM/6IJ9MAF1uIIz/yqWbepo1LJNFc3VY3tlT2JF8sPk1YDHenNQZMb72AqK2DWq4LezDgLwAh
8wn6JslWOmouwPGBKvE3jJVmJQDyO+xTBnVRRx/ZyuBoP3zxyQCzkwUEvc6CfNW9lTSFcZp7GiYv
sQvibK7sWDjqFWU+Ko8KjM/Y/S2KQU4gDVcnS2C09W1WF3R+1Uz3+7d1h1CDIx2E5a6MnLDCIf0f
FTOu8HqD/Uk4VQZ6UYwjoM/YsAVTDbZ70bYJwhUC07A6aZBDpA8ke0DjxCj4OkEYc/hUhKudpQlr
7NAltQ9WIuVUT3dEz9xX7X/l7dHMprcgM+zoO/pH41aGLBHkulMWMgukkPp/9w6bC7DXtLjziloB
RSDYtPQR5tm94AZrbiH+QMNyT1gbELprwQAq2UoA3zpjfrFCCKub+qgfdZYcf4+KzXCGq31roAWa
muUjisZJhpIpPZx4GmutBl7iwsRsSmT70w2MRBWM3zsyRHxJv1ewYH2w5AS7wKVYWo2sVzym4i2L
p98GSCE+Nmt04rQFAdi/RBJn54XtFqPzEhHDAokdkTa47qazo+imW2f+iERGoC7NzVTVnK4D7elG
PAH/agQa1CQsMe5xbfZIVJYyL1f2A4Ftfzkqr4ViVYu+8MqlZJ7RZIuo1y0yEspykKOQQZ5s2WZJ
OOdAXa6yBE+ik28nLlU91sNC2hatLgGkus4dDUvgvlN/q639pY5/HzSoWQT4bELnxEI30rzmIO3y
O4aRxjtRB1ZmRsfquNnAcfWsE++WNuDeuDILpd3enEUUFu6FKCvo5k/cyhigeuiu4wTWs8eODmkI
jfjOj1nUYMaJ/DpXOiu+ZrVtPIdJabu01/kXtSFhB669UT4uwj32oLNBSCNl9rFgOHgJs3nyKjr0
NPGYjuDe+fX28nXeqc4QGyzyG8L9kwJzLKzmxyZhXXNoKn8GZp3d5a5J+8Po3CrpFpIYJaUdiRPq
WNtI41ULvYwhq+ntyQJ7Ogna7LUeMjRrfyKYpVdGerZuPocQ+QgdPLAmkVgLpsSFEItmp3uCmer9
znyw9dax/jRxFpDZXoBp2qEJSXDyF0CoYVg8MvVbOYuElS8CPtZoReEdtS7NDZHuok6oB+swnTPa
rYnLnyfjHkBRCBBckiJBlUFP8T7AZCf508S8V+fpuIVQ77mH8chG/o+55/zYv/9fQh50eqrxQ2Ip
13k3C/bXUk8EzusDety1cGj40ccOHqfV1QpHVF6CuiGaGOspyERNPN1zt/DoUmEFw2XGy1XheEb7
dzhV6Tm4lYGZhN58qCV5vHlTQ7Z9l4jAqHQwC9VOqq7a7MTDaR1j5g/0Ffn9RCoydWVHcqQuPewT
PDw7tP1utnHmJ1gC4LbtBjM0/Et3MIrJhT/13L8es0NnAFXGvhZQFNI6EHBIDgGZnTx/bOl0v0yL
iw1ayF3SYtJTl9yPTz/21/N8FqJJtMjE3xQyKWX47nrEudvbzF+0ds+vXAFSOgIBK8miXpFpETPG
5yTdrMjXOJWF3obluiICZybYbdf+jedYKBmUbtK4M1A4d1pOxcRwH/IjJyWYJ6juaQ9BkHBDkuS/
h3160pzYo+jR8Ckt3+aQT2ofwu5z19WML9bniC5Trauob3WWWswBodf3KWdajLHDnQTjSIOoCOro
aSNJggXWHMxFkUXhF+xdgtwB76TsK/Wp/Z8FoJYzOXJl0VSu86g/Dg+h1tY20biLF7IHClJzagj/
H7cAa2GTu+Xw9J+N22j2FVL4CAOjI18xgbZhJAWF2hjPKriSs3fONbD4H75OvFwhTcIX82TUPGfR
aPxYpyEbIfKn7TE7wNwqKQBjU2LUHGUN3Fhj/+DKQrCy4sjne4Z6VxCcY/2gLnNOO9472t4c/I3k
FDdUM/5XtgDlPoGxjVIOBAsxe/JEQfkYX/WhjEwwo4Gl68CHyijmiwlx2nUJ7Vo1y7bVaUSoq5bC
WSdtjueI8HmYVjNjn+8HaaaAXOPZ1m2BScQ30anwuueaBtTBX+yexiDSIpB/9huu3VR3gZ/sEYSn
VYOtyILHk39ZXuaHouXy2VP0HmcYKne4k3Y1SPR8porMfnQRfRNsQXAF/1Y8N2Ec1jXqk4TdSnS0
g0R84V1WREpCiu/mc4KA33uOqq5PeByDleJhFrmxxn1YSVP4gMqgyy1ROCoujpX8lQhle+3T9Lu5
9JnHpF5O8rA+1Vw6xz39hwoj2zOUlZXE8vzxrPm2WFsro3Ci8y+5A6tgXFUn00fRbGlJmMtGaJau
p+RyksrDC2XQ92XQJOJL4HC081Y+xg==
`protect end_protected

