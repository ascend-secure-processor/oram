
	localparam					DDR3CMD_Write = 	3'b000;
	localparam					DDR3CMD_Read = 		3'b001;	