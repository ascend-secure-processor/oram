`ifndef _SHA3LOCAL_H
	`define _SHA3LOCAL_
	localparam  HashDigestWidth = 512;
`endif