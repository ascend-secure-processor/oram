    parameter   LeafWidth = 32,         // in bits       // TODO is this just ORAML?
                PLBCapacity = 8192     // in bits