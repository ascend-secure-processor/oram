

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cLJLYG+eQT697weLGw/M7+ydzYpSUtzrFP6PHnuIQ/va48SWlGG1JfVbKOSSCc8ukA6oXFsdqmhD
LdTRvoKWhA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FIaDtJzqf8jiUAUGWUUVl5F/7pvXp7KagR/ry0lA8QMgkF5BeMrzQu6f0u+TbZYtPsNNuXhzKycs
LIm23ncOzuPVNPpKtv+L+mcKrFOJ9+5nVeXlCh1AFkPa6Nlv5P+S7Zke2oxqFt4lcMc8Ay4H3HG6
XM35fRkLM4fWOXU8CqA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nqjD6/IVuqiOLnLEQ3VW9Lk2KqpTgI5rNOnreyg5CBREOW5kogNwLYR5x6wlNGtcwfLdC9flDvW4
npW2P44CcAUXLBGZDHj4GVIpdJddJYVHnYcEuF0RilfTCn4aJHEoSZ5UAyoB9qdaCSwi6ppTuN+A
ske89F7VT/JHZOwgeP8SKYPvKqQ2qjtbfv0gAfC8HB6u8EuQXJ8CrEty3ZkGcXfZSoQFoUqrmm/J
eQM5IzEDZ1pa589vEXTMXSxr2mAHJs+u0CbyOfbwVZVOzwKD8xoydrmkqjSsNYqorNcvhqwE80g/
GiYKR5TiLjIcBYgEDyo5ux/1McBdN8wEdis8TQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0ef1iaaywoWYVFWWA9UDGafO0ilqoJ9ls7n6vou0iUbDAm9sd6/JgIpjkXG2SKSSl4Tp2ec7lTbx
CtWZK8Dmk//HJMMNzN6DqFcvS63Rz7CbcEzRCF0TExaFfzqB4Cy+huT6FkggPlnSI+zMqEUtJJYl
JWhj0a8brwA3SW7O1RE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gg2wghmvoRzjJGOH/RRay/llr3/p/sPIopiFDld4hlS9GLvrPwSV8yPxrqaZJGrT5BR50aEJgRES
0PuiiRekrcOK7Mq8gTMAvy79PhPN07RkpT7I7qLVNqQvhJI56+ZvzSR1T28c1TNzj0BLLXXy7zQI
V9ZS3I1FI4UnTIhnyKZ+ACt2C4NIrRucqgTEYUCzNh6/3MORC/QS22Q0MWy4AOhYT1sZcrD7UK2F
9NMQ+sNY+yl22M6Gyml9S/uuIxZdFZqe94Y0ItPFndaRemLSTDo/SCcDb59qSqPut3lELhdzY3rz
+CXm3YBlM8pvzxWPG4FbPHDnTRHy53pfZTveiQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8032)
`protect data_block
t8vOK8P56YpOmLB5Y37A8sKfiSKs2sqh/goAEEGI0/F4EV1Zv9z9d32sKuWEienwPpQQRAj+7ZTt
TS41fzRwJuuNA855in8+WkQMxN49UIDIXUoF9hBCyqK1FYaqPQiUua1XmQ1dSmO6HlpaxBsLLL3q
wXAloF4nQSG06ffqBuMsNNrC+Opc5kTo0lLqUFBibaW/0xUYe2OerC9JXQDpP2XVX8vOBYm7kHqy
QgX4KgH9ke4M4W85/qHNOtAU+PJEoy77Pa1NIrnJKYovrh6c6qwDD319ZsIhefOxg85OnKbIJ9xr
d48yQMlDLLTkUOu53FQpSslDHSxQ1ZSN3KnkWd2jOcslHE5l5imNY2rNZPPjStlS5cO+SSBKf/Or
Zlo9NCCsCnvXXJ21oH1Lw4OGXG8CeqkbxblBevggMjlbY480wok+FSIliIVk2ahvf7Y3bznJBO2O
F3dErXtDF2wr3sVoIDQAgfqz3Ct/XEVdO3IbI/2WMKqN2GUxNKt5/g4VgAa7KJCD9/q0Lui+0NIr
BDECg/+unI+X55tl4qIeH9HA3b7gqai52hCxzoK7Ys8NxclwY14rzyuWkS6S5ncU9LEHIH67AyUE
anlr4+gGblpB2kAxn8arF6g8c1Nz/dnIBO5koEYt5sX9y+dn/Ms3mUTWua1FzpGKI0dUkncz/HXx
eRhdxI8G0IAFfksoNw86y0vBbSznp2ooEWTvqzzHq7y9a/EnIP+hk9RGyzx8uyd5blcOb8pQszhX
+680dXwXRHHgg1TLEA3nXxJYQOp9ife73KVuaYvwxLbxQVcK6VavzlZ9r2WjDdVhR+Tka1H+fdlq
rc/AoK2jIk80wzl4n8NR6HMwPc6ZxuGOM5HJjltyG/xHnOiMeEq+eG5djI/AvKCiwXyVs9jfCW/O
jAl7p7I9MhXLHC19Fe0YsiOLd5cCRMg+tgFh7O7ClWrDH/rsH7rrXjHdNGk8FZPJRCYos5Mhvy5O
3wsRekxl+K8YZDrUja9/miJl6YQaFq1hnXDfdVtru2Q0b3GxLSO01fgnzKrstS6f+rprXXf8bxm5
X4zUXiuXFWU4EozMxy2Yl7sLwVjscQqldobyOCE2YZm4KFYuQINQtSX96gbuVZk3HNUSXFXlgD6+
zJbKEnxkkg1LSbCFkF5kOiFN9pCN4Dxo3XBdG5cdFDlXmxAUq/gxrPb6lu/w2z+q9txpuCV4UnWq
SFzxn4s3AGLictEy2bboJXqpyXA8VzBtxkw6BD9f/nDTU25jIy57tGSSMHfDoF6EobOhL/y6E0Hm
5Bx23ndaVEueav9dDtvghpLV8yy+62VOh2Oxpc7lrXyFae9Y8y+KfEct3HuYMSrZ7nsxcOJJq2nC
/lrz4vT/HMAozcbmAxSSIbcSX0m2klCUiSczCSRtFOyoJPLkSYfNOXGb1NxJHsKnlZ2tRDEnlCya
4QqaTEBAgPosRVj6fGF93PJchBZaqnc0weRWCJ2gq9pMEwwYZIPYHuNzl+RANcemjO/qGgiqujdp
FW0KhjOkJ6OIdWWjhMWZiaeTGfGoeo6df6h7NcBJWuuIRUIDK3Y/XTQoYYFsKNH5F5cX/u3iBTg+
1JDEDK6TUByJNGtqa8jcR3Qvu1LZomQwqRTq3iLckSid+yC3/mf0a1ErCoyDBaJeF6dEiDyqq4bF
KDQ12EhgBeI7LxD4QeU40HevrolUQrp5xP/ko5JWk8Lxjms9bbz1098HypLDPddGTT/T61UoRejU
twkQITr1j5u16CxYzS1JM282JsQZIAf3+uAEto03ZychOwKhGOKEA639tqafQmQCccFRnM0WeiFy
dtxDzsH5Sx6kTIGs38N4/y8Jh9NK0sCn8N+X27Wo2OLStqPa9GvccGn2h5zO6gecdEpqYX5Y/grV
B30OMOsaFWx06DteKksrI/zJLr9yF7XbrQbsCysMT9LRa3sy/Ilgy0KyyKtkKCFfYv6avv/i6RmP
0Hs2vzePXzsl00p2THpjHU0Nl5hw8X9h8CTj5B6EoVKFoUZcPnyjJM+JlHyAV95gb+ezgKKuhDts
E8hA6MnE/yZ2Y7RbY0y56YUIfnOpL1M+S3Lm46nv94bIj2ccQicMk+NkkjKKlJG8diLmG0A+veaD
YabCnKWIyxSdG3oUuiA3LjYIYpflskCfiJkO4xHORXKwmRh0zXlyDKcs4wuIzZPYF15T5tvBklU3
sAlxjckJKYrRlldSj1oWr/APSnyxSlEHUSwNh/RGlVhMW9SDN8kqp//IMvlsYqR9SwjJwoBJ3Q3n
unYVtxiJSVRwSZRUsxvWU1NIa7bJOKxq+/8wZ+acqggZBnq5jLj3hlTIZT4Q7es+Py+paYEd493V
qMfD8YTRc2S1sOVQ7p//kTp8Mou4nAtbCrcFm3sb3GaqQzFYshjW3cxjqCA8/kw4U7/RQ+xvHqMw
JBUFXckbgrmxx1vECmMH+qr613DtcqXqVSnhg2Vz5KLkkuq0KUXpMCImhjKAXI7rUPZrJhsLnABW
gJhH+GhkZ1ElV1uzubTBCGPyAef1Yb50BPNs0DMWkpiaZiAe6XMc/5TO4PzvyB+nixlqdQ6p6DO9
R6s6jFDxynQgsgv1yriIPxP1MR+NIAzr/CViradriGKRItZs7nL+npz/D4foM++DaV7H3xWXh3Sx
Iqj8E9ZbiX94NeoIX7CISwvzvNZ0Gfx4Yykfxdx5YJy8QrWhSkKGLgM+mU1RORh19GVKHWDxX1Bx
9bVhohXyq02iap3bctARBiGGWkAxVwwQn622wl3Nd7bPlMy8Wc4LtVnMXBHQLor40pi7xdKXYj18
lkyq1Bhe0iGOlWKPDJfVaOeyu4E8opNul2mLfFkVU+xNMwTM2hiiFBWaW8dQo8JfCC+zbMQRrdvO
cnvoRRjYbAQH/LV3Zc2ev2CAm36i6PeI/D4skvQGV3kIy3Y9oH6WQOYK5HAT9EmQXHAgDS0+Brzn
tbHeoIS7VwJqMA++cPBcw0r08qNx8Vw/0/L5Za0L9k4RuF9CEdZiYAKpBunehiNr3WEJ/C3uxISa
3J2ur+xotq0gwryOp9owqTV/MDRJQQagj06S2O0WymORYs9dp9xb0+uvKCwPWbt8I3sIKOqcXkhr
AL++BYSGgCbNHmUvRbh/SGmNSo90ZplCM20UGS5bgwwN/Ic504PdTRTWL9pe3T/9uh9q5lUZbLes
nE20WWJA17aNCVPUglUq8CHts+G7L0/1KtfpOlXQBmiCUgvbPaoVujUzRO0JfH1d5H5xmWDyX6Jz
dffPcIH0XU51RMFO2Zef165Z8FS5n07jcMLj58XzgefAedLCXbR5E+GWxqVsPE/SwfsZPh5+XGa2
QDbpn0wBgPVKwfAzc5TvaTqysINKdZcVXjynpFvvjEnRnjxwhinRG9vKTYsG26s18tUx8saKmesA
Z06Dx/M3fJgScxUaQNoCdfprvvcDMG85LtObUUQVs+4tSAl2Zv0U8Rta0CWkfUHcefiFBDRA8+mf
Q1NQ0DziuJqWQZWZ0T4cckqQkZBk04447Yur1Pj2oURZrpHgcSC5ktUzRQ9sHKIUUjFLnxsvreW/
47eHjtJzU311gOMk9MPUcoqzo/Aae1pWfdmxrTP0NfD4bBjCz1Rkqw9pr3sPvzmT0o1cmtT3uJAo
1HZUvLWmRYi9uMunzz3BwKsT2AKjvgl1F+XZ2brKezyX3WWRLZ29z3ngST8CvmJXBah0LMDXehJx
H6bccjo73bvzCDZ7r8WioKLJJcPRlqX1RkHXGOXylsuy2DndII+RPmILmTUrM7sIPsO9sKRzuto+
6DRFJUUw3S3u/qbzCezbqXr6GV7X7fQeuIAjQx0GpGRixYosZBvA6my+CNi+rMvu8EN9I0GyTrPq
yPHoWAu15SZiLEKzQw9TifThnUEWrRsNGUoaIT1vySCfQqNNqsMUazhL72VajoH5DGDqLadB/eeQ
9IweCDkzKCaURJzv7TBlz1cA1S3kUUfcazbWWiFGCZv9cfxAU/j9bIt45i5yQmvS1rrax0Lpxg1W
P8cKy5RC4ZD0Oyem8d4ueB6sYioMm8ycUiZdKvsWZMvgWwVvZK9gXan2Iz2QIChOq3E1Mv48vz+l
QPhSOkQSAGKfFEMfLh+J85Exy7sU7nkJ2Rx5AMuC/KMi0eEIzcp8HNWgVG9Vg9TuRl9qwmCvdmuK
5tCsX9WXi8Xy/p23d/pqDpPM48eNlwDWqVIrqzQJTX7DtSjAYAzKN6E7jwYvJ5mSmkbp34Gbns4K
Htcqda+1o8ivbNEX/FPhhKSb/1hD+uvbAu/aIgOxuLAoRUsh6b1eIsgrxw4Nb6hSYhhrbWZo7VEs
qw2jRW4pY1YgPLmuTwenkU4qK3DoO2//Nww1t9AeTXFAphPOvIpI5QAPheood52n1RUMYMwqa3WK
zrA3kYbUna7v/barLhTryBwu+M3Ad2XIpZ65yqDeQZWZRztvoSLERN980krgGyzYYjunwW1PySMx
VB7HyhUqbbcpmP+PZT4FxIeQmMJxslpUyq2aLlrtELfioekj7zJl+uDYO0PelgLBYmetcFUwbFom
4+CQ9r/pftJOd70aqJYXwsI3vnr6kitH9LhccHGKlAVprn5LAVcPeB4oj+bGnQAfEe13iyUgPO9V
57Z1fSwaU6hgK1LmDXgw2Au4EKVKgqtZCRrj7jH4YCMYKp5pnDw035o1ns3S4qo2VDjIJFc24FMd
wqcUr/bTj55ILIwI5F+Zq6IuSA6hLnTP2NFQHkwB5gl4m9EfpFg4+rPPQIym+grLGLvRvAmho90f
6xGE1MzX6p02tRd4FlCCtJKFQD84hfAh5y1Sd6A6uakcENusjNvx8mqgdsOa+9GMpbsM+R9zRvtZ
lBCb0HdyD1/H/jgqnXGRK5R3FWbeOZpOxtqXYsD6aqxBPeEyF7QM/NNqmqbwC6oac//mASlBjDwe
Y1Cay9aXUJ8l+2QIHEHq7OC6aqJQ8O3Ws95WXyPQ/7IyRx7g5owJ8z7S8SwAnH9q2NzAJwu+4Zen
8fzg9dnY++CrnkhQsMInuzzdhJLqmoox2bsIoWc2w6gPrHkECRvPYU90WW8ecPj5o1yqAevNFs7N
GU4YaVI8rpxXPVed6Oj9xDUJAHDY9kgJflEiyhVminhkn1660mrk9tJsW+8+FO2uqiPHV8cnfbji
muk/HIJwyYLTYSG648Kji2/YIMfqxgwS0PV4BnYHpEeh3xZxgXtOqRNy81Up0ofSng/x1/zaruJP
9h/wfgsKgr60pxPDxKU7RPq1Vdg34qBYxNTbijbVuJoCS8vSkBPu+NJ0n8IljuAlkMsh2QasJMpR
xTzkVmmSQ/tIl6kIMTIHWOcsIiGQPLBLYu7nRp/8GchgRueIs5Ju4BvkQKZ9g/AdTjLV+hTZ/kOz
GHa9MtFEOkTVaN6P6tPpRQoTS71i9jjErYgSJRdPOGvSWCUocALeyQs96Gv7qDNELOwMcXXVc3zS
tF4BEsz/4p29k0pNGeUU4FosMaNS+0hXsgD9BJf6oCKlsgI8R/+xkDRzfcm6plsKQ2UJZ/opSclA
0yYQ+cKdl6b3zJwHabBmMg6vOvO5WNyCpt8m48kYuvli5W6AqEM73QUwps4mbHDxh6zSa9LMCcvm
OIcdDcRXBMXBRqR+wcOXIJ58c2vGxy86JNazQaUazvsG7akTkSeiVxxKgT66g398mLHGp9TUHDZr
PqTFH+BJxnDweBUVvoitFpts3Nb0bf7lLg+r9Pw2MAGLZ1QHD5YjT3rLQLkHFBpbisp33P6hKE5n
Z71zK16vgaqC3QE5NcQnkzVnkXpo0bzXZARtn5xpqVjtFFBmcpQksKsUVAI0nvOCve90YOXzx1o9
gCGZBplOu6+YU2BzpoQTmKm1toeH+QM0woCD/Zop92UgaXDfhL55GTp/dMKyb8SsFcT+0RKO31m6
Bjk/JWWOLf4ejDTp48c0xFIqyXnDJ0ovLpjub33eHA71QdPCR1zlbr+iD9bLOIjXTj2x3DwFhbyd
FqOfNbq+hl+JrSbaYSTbSRA/IvzcTag88UEf5WdJ1yLrCsJC90CmacV28AqNRHwtKUVEtT47toob
7dmscDsmI/s0OMdnZg+PrQ1mx+QltC3yGUuibU+1kvE9fWxFfmhVPuHKDYDE4g84VODbIytkeFgm
Ga6HbR8cla2/OsmgdxutrA7o5W2uycdbiGo+PEVkdjYMMrFs38eVgp3w61+pEFS/fhRw9cwomXNh
+eESbR/RXj3qwOMma3u3a/CnzBWyGOlApAO97acRcYZ8NgPXP5BhpINrKSmCzpNfRrqV2knYwVhy
1J6TfUM9MxZBAjtLotBDR8PFYx6VFMBjmz1pFdzgQNeYK+rBrXyn/NDYFtjSBhNPlG4B4X4bSv5W
oZqpww0PwSgmZwOCYmPWxxN3YargNXy0ww+sz+moay4Rfx5tRv8doLhCbSyat9pv/eDZfn4MEqZf
/f0sQqyFRNdIzfqV89Fn6NPWuPe+Ujg9AWp6eZRlk46FhoZozHsCJzB5VAp+TRVMcga9aFS8gupC
ZxHCA5Se/zEas2yAQaTI0J4wjAAob+fL02LTL7ziASX2KcohwYywc82bwCU8W5NljwuQ6tDMNaQ5
WsAlytY1gMAsB/U4+B2pdNAGgQ6WVoL+RleeWYvID5qYkyYgvkaN0LyudQgacKSfhcbl3K5B+uS8
CLgSZoujeB6kLQa2VSyq46Qwg1AAKv5KH709n5qUjndAYInzGV6Ti4k2YU/1TAmuane4Wu+/nJHb
3KvrQHD2o0dGb6VtDtwW5eOMsX67izVjxqS2fHqG2xRv396afsGGuugWPAWMy241WUs4wnJG8hK7
n2bLgm91m6GYDkXzLD6qwVrZ0wohN2XiM1EkdBa6mAbWrdm7HD+lwc1BJ6GgN9HpEHObXIBb2XIt
loJ2LeCtUo+AqGvku93rOeJgYXidCXmrqEDre6g2+GCnP1NiwHbz2fwaJeBLyMfSo5lHmWJ3iMWB
HLJrJR8dcKfi3bUyVTuhK7PUfFDRTMZMzqj5N9PGVITC3TAYeNHHvX0pOJXrhN/l1E25QcKojOo9
1jWzTGSA41JDMKJP1JBYNmSDZ/F/4KjksoZZs7AyY5Ot+cCQdDSbVB79zB5fiBMGBiGy8ktTQZYQ
YXx/0uw/U7OrqWY+9NMPyBTruFJ2f1c8lxs5TD3nnF6ChHeMtmW752A8A+kiw+L9gqIqa2OOCYEs
KKav9E0RBBSJjY3CJ7Oj752YGhJoXXLUR70VzF5zXW4JQh06HzM+IQj+VxP/Pq6uQ1Jf1mvG9KoT
zHhEpDMKAIXLQOLYZWMt0n20XPpLgkPJihcY9pM33T87U81Jf9h1GtcVx16NLXbv3eJXdMadrBYf
tgHoP0Pzv7JFWPOEESRXCgT+K+YphBKi352QippyazTyQk0mCpQGir23QlIfQ8ZrQQsBL8FuMuJ2
c6LxFj0vkyUs0/TQZwxgHVKjR3ysafKoNBQfxWUxmP/hzPE+KdEGzwS1qVOx4GYv8do/p3JPcbLq
m59jYvx4KgaM5eb40bKbGCcnV2r/ZjzKLEzpkUisUPnzwjwdtf60NQLyKmC9oG86tAqc+R3xt9Qt
ai6J8BUaDaA2uVdLocF3cBYdAJ5w8U3NS0BGJAaPPL3cl+HtVCb2rGzGlkEhoC3zES7aSml/SDC5
1C+8YZtdGPVB/O8MYHXgpdaSLwwfeUFP08Ig2khJoqofWd2OcWrPKeZpVsjj2xWKfudsoFmtOteB
et8f2zqfcki2zPeE9BO7pe3OZ65UAK/nifAOUGmucL0RpoJGtOeJpmzFb1Z+vVvE02gBcnkQ0c80
uBAp4vzlhkgj1gpDk3odf+2LoU+yX3TkmPOCcA7K6R5KSCNb+Fvuh76aajvMtdxyxU8Q1qnwQ4QL
KviUbeZdLGsWZI/w6+0YNeOzuyhHVwY4BGYIzj1DVD/wQTuVAHi9BXRKIN2bUIO4rG3Uf2dsfdUd
IPMthDfHOIJxxeZkaB37VwpPxy31KHBuSOeQQLIIC6yu5TcxvxgUB0YOwNwvalaHHj09LkTEioFm
C3v6x8IFLY4vMeWt1aR0kt6r/UixraspNG5eydEKgDp1JIWcpn/rLpoNV6ykLYPi006a52J76mpS
xS7SHxkGYFbfgQiuJ4R0T64IRw14QdIamYhvSAxKZYPEPaFPwo1Q515z8VQbOXl0wqGhQl8Duykg
ceKCbGcOmLvtc+W09dlMzbbBBzElvZnBb5CWfigEgmPsbZ8xULm9Vw14bIRj+oq7sBVjhHDhg70l
eRffTvfpMVrG8vIijK9lHUpJe8Cb8gB04PtSuSGAVot/2NreGutM6IcEaPY12wHMa9Ftp5hgk5IR
vdgTNxvyXzKC8xhAwHveL8CTd/IgAcEISWLgUeGHF9ZKwKAdwkGfFRf5x5+Btv4ozxNx1zGOc/S8
5BBau5Mf60n659KbhdPx6aF1LgS9wsjdL0+igf/EiITaU2cxdAix4AwQDEOj1bVJgg/33mID/L+h
pZLS7H9Q/UtApCE0xfOU5MiixvALvc7Bvne7g3amfc+ySBdW+edh2io4/XBsqofqj9kymEDgSP+6
rVPqYHLq27B3hh9rQ4DxFOw/3Nwsxbtz0eb6vPJrZWunGovgvPKRq/NphmHpucHp0Ax6sRMHeCqy
siQzsMLkZKcm9YRps444u/hSgl23O4kp2WkM6bLsVvtDJTdDPSS9xnr+fjGU6HqMDbvKx0/hzUK5
mZQDE3iHyRAsFj5dXL57FSOZCwvRl6sHtzxPu/HAJMfS8xT9fioEFVf66UiqPt4w3glwrK/btL/T
X9XCbkTD2RZ9Eobcvq3yX3whpTgYl0rS+7PK/LDpf8zqiKWhDEYEby1LMCkAPvdc+7rg4d+CX/CU
uNL0yZEdrAYaGRngubd14WIl2FqfkkBjA6MAoVJaJ/3WQGqc7eqWRNn4e6AgKvJQlLQ0kRernw6f
J86Da5vy7xWAEy0BXmJR/TZIwSmacheaoWAQsGL+nlJJdoB7HCD5ZDyGGzmJw5FZvC5zurMjjVEr
cK36yfuYAs/zhr/FF5di9pa+gg473CqvfdduWry01eT1ZiXD2mbktx77EKKehr2gEyQWT9aIcZ3v
Ht67d6oFdADcUKjDDbA35cojaVb7wFAVfEhjskIRiJjKrV+khp5vj3E3CBmvLDoehXLVr8UA+HQe
0CWHBGSppGtrZG6tHOiMtR6hwXF0c9aVcNyP+6ts7HYRrpcE6lhMfdE2JC/SK+YfYzTmTJ8LHcIu
EXHDAvySXByBeuRPWn67R3i5XgVnId1cMq9UClckb3l807g1CtF9MGt4bwoLtqwjSq3+WlCGrZ/I
7IXtWDeBpK0/YtA1Imq5tBMdxrtq6i5jsetTTWuvxPHW+4khssXDTiHos/ntkuSsNKz7UIytkwlf
mZtFrfj7vc2QGw27lSS9r450YfejX9wgOEyMYzzrym2l4TGRZKLftIeoqPW0YzGwAk+Yp9q5MwSP
PHJYgkZD86gkFuyHanWmgLd+YRLnBdjjGOuPDkhTinvFPD94I1SVpK/4rrH4H2rKG7qJoQDHC7M9
O/Cu3p9ARUUK0XNdyh9b7arF9V5mXt4sIKiImzBIQnVNO4GHETCyE4JK+Niv6QV9ex/ROth5Okaq
e32fdKbbw/xBkW9xdIf3kmq1tArj/UZD50ll4nqfkWJrE782fXpo9kT3+WjPMJAqP48xHZ6E4up2
QK/Xe6jPaYQB8KsHts3W5ih8JdK6qnZ6Nz8hddWLMK5+L1y3OHEas46yXDY6yOJ00O2F4RPSqq8w
ht1yuvX1u+4cWswksCjk5FPf3hDYowmgrJMSHy4ClE+8SRC3+Y1tCoEysOxpUWpj5djZII4TlIKA
hZ7uLYSCdw6J8TECTAdH7CZ28fEgSq6nT3WC4KBy0/FrHX1qK7mVnBi3RcikZrV2X2HH3BVEm1A5
X5Axnvd8KVlF5YiGCBUVIwH1TQu4QUYIcgKznQxoHaQoTacYBrGp2vAfNKup7/1Z+7HmkjKGX0da
e5LtxkdCKmSw8M83xyBEPXjkZvLbUSDg52SWSQAFq9mCRNMBuNDwA05OzP6Yb7uGo4oxw/MF+8Tl
FtDHbKxH1P4RTELPPsu2dKMMlW9hbd8eJEAQvUSTihTRHqDnWVGmYNZLfrRG2e5pUkghenn8q4BI
Lw3EVkZ3VErBw7i3fqolWRVEsrra4LyOZAPeHkaqmLl1l2FVP5MUaQSK5Tt1sh56MxmLB92duG3O
8eyVtmXcNxeWflKkNP/IPraCARBHKyPmOmiSzwwWfeOvwpWZvfDTLy8kQSLJNv4ygi2kQNud1mrM
l271HmspwJoaoyaswfrcQUnNV0WARutzWkY2QudC+E7tT0fPPOHFvMlfhDhqI5M9Xj0A5QlKBreT
tsBqNQUytNKznnAE22HOcDZ+sSywf7u0Y9Rf5YurIOalY6NqBqg2PkbUz8pC63NghC9nPv1BHVgO
+Fgx+7Veq9WpdyKb+4njn+zITKEXpsl0GMstQjXDC9tDxAvPQ534OLnkqhXuIJW4OV+A1l+m+kek
EatCcTkp6Y3Zw7BxuY8WOkCoP8Q51dEjk1R3iTP14XcD+OnrxPtqwxGpCWHr6aQVsdOip6UwgnTz
tNFzR4SkQvUJgFYKJhVwF4O5FPQNrSKcNplGmuBMhhaVHxKfQcFNF9qj/+HH9mobixGw3Q==
`protect end_protected

