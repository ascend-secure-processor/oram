

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MmHSU2aymsPkZXc7ZYzxwfKva+xI10RFNyTiRqijQ6tU/Bc1DNhEdxb64oceqoEx24pqLcUoY10G
dqj9KQFLNQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k5bAYD4ecQyGQiMvnBs0mw4nHlGHol5epAlLItdjUy+Hki201+9ja0Em0dAdvrYJPpP+4zjBvNJE
bHZKhXLm2SY081BD4RdPlFuoQfQnoe2NJyjgCNN1o4liEt/PKgyiJpsmyDk+hqVXEykyxS/lmr2h
9CdFQYCAhEVEfkdKLOA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EwiVSLKCERe+Bjcev8JmoT2f6dd3LazWl9zAZB3SL2q0SUqfxkHHlBSPNw7OQZsHG3eE/lotziQH
1MMwwT/VZWEnxw/DiL9cvqDbXFSq70wNMdGGPqOok83kSvw4+cJejlbB3U6sqJFEeftmCOga3qxF
Zlm14dARySCqXDEYiu8tasB/PRIpcgDdblYOMeZPRe2fzbYaeLwx1+GlkreO//EwRoqFDRDjohCz
2Qh9WoCZc441c0rH9e0Ua07KBhOddM8GnbQuS/a5EKcniUPMxAIZPeCcPOLTWTVXLzFHo/rVlVYD
LvNTgnUJPam6J6IhqJsTKVTDHXO2WbQUvdtXQA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LcGga0Ps/lJvIfWMgrQ0Mu9kJ1ZyxWqqQswpigXUOnHjoUCBQCBNE+wJ6qe1XcQaKijFhoffX7oD
il+KpPmVSGsKgRxc1zNuWP+f0wOHsh2ofUoJzXkmyoxtNzjJOCRucHlaMaJRfx9fXlRMS3VPLbe3
CI4HmWxUenbN5IpJMAA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
otgARbXqljeq3ACx2fUr7TfjeBoSt3TlOuI+B6WZNv2WwS736+RhShwCYxZCGSTL2WocYZ5jhIwd
Mo7GIy+2jcthGOUKUHhw2qpPzwwBsda0A9oIgmSThoZlrBcoxx0AO/KOjY7yxbfPxM4bznVHHM9q
tRX70cyqze85n0fiiOD9qcOnv/0FvbU/IPfSUld1G0iEod1J+nz00fh0QIZ/09ljdwLnzPSQg5Da
hg9sgcCDgeEF5HvUPwTwG+Jx4aA/zd4CCwtgEhQszB6yovkPrQKWwaTj/5BUpSmAlacieA92TXUD
eWhbCTpf4DZBYhdDz4FcSH+eQdmAGHj/rTxkaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17008)
`protect data_block
8QmXOV64u8vv8L2sdGCOLA6eGH3eCPDG21Lo2yXdgFT/cG3fmMSh9SgXZj9dcqmVavFejhiA20FH
Z6qNLQqkJVi8PFSl6zMb+hUDkslA6/v8zV3TZ6bJp9hNkGIc+nYZ+8t32hhpFceZsYskdac/l2BK
ikdq8WuziQtlVHsX9WYNF8tUnIZJPme13wiU/ha9QLqAgsktrtWvdYZg6YSAr1Aly5G18Q90te8+
ew1b6hTadvxK93vedqYhrjVfFRFBpGgIi9LJUKgK/F/17QCeJiOG8aQrl4I1kzkBEDgQaUG/O2kI
CFJJwlMFcM7QXra/yto2ozBJdPfmxSoCOQ6qOtNh+1R0cVowjMSG5I8/zz0yppetRSZs9YKWs/dy
obvR8Zi5WjjNGu81xKPnq0b98ug6/Yr34/OSpq0GX4X0GDyM4LWfkHIxjBbxYYv/r5PnvnmqjIzq
wzgX0f/1VaWlNyaKzD8sGk/R/HAFG2wNUrN5NwKgQZYYkJvv97Z4pdF0lKxHjxrw5vRFE+PUIW/g
VMt4YKcQTO9lz8b0TP7s1uwiVH8135ADhy5l9fyj+dbDHYC333NTo/QwDvcNPkyi3o1jcOCJ7pmk
VYxMJyRkGoqsCoiKaKgplCmisPcJ2fgCy4O1SpvTKEXsbKXYiDuXg3krvKBIMpZRGV0NlLLb6ftO
X9EBN3iMZKRVxsnPdsGUvESKb8adqBE7R2AwOxAntQ7orjPst6Ey8+iGHMN2U/jsxKidrKBx99jD
xfT5yImzdmDzGdoOYSXe3zLu44qXyK5eZnkdiBppGOQ8mzFmesvu43cwpN/oQUk+T7c4yhsaEQ5d
VpR3ViBMVAo/Bde7jWbsT741XDk+Eu3ZgRr+ry+TTj39sBy4WEtxN40/GhpKS7S1F3fxoNQXLVfN
uytaUpqKukBj7XEpHHt4lvpgczFnPwQlxatjGvadZ7MvZRY6DfuhlFzxozfrEfyUGibv5MMEpQ0k
AcnHBr6idk4/mBgLvNJ6fOdB2gT//roTYxiHFbL8V96gmkSUg91TZc+dNekj5Rzbf/Rc7QnUbjrQ
crdE6TrBAjfEjPD0q5iiK6rthStzukjLXTK6A+jRs7pYkSJThd+9i/wBGaywQ4TbUIXDEVnvxXkm
WjeisXeNPIOngdCmY1Do7WJFFujIMZP/jjpeMJLAHEYL1AqxRe3e1Xmbn1fkg12gPMr46VsRTkH6
+/xGT6az5Lgq5iTxHDHh1LuhxExXfH+ukl/FZxcCnXKGZIGnn06yI+2ibBNET/ctAFnoPsST5u03
nruRyAuPhJbAjhL4VP3txF6DV/FomPTybSQOeZoFDaNoH8WaFpojcHCl4uVdI0g4vXAQ+150Dfb+
LVF7VezfUpV8XXgLLQx/kEEd1mJBANc5KSGHQLMg+h5zjTkDV+mJ+Atj+1B2vTdq/En8dmoW7vkb
1xJnKQs1ftwn9nQvZ12weaQwZD9mCmS6MIBc/tXW3JPRvhpXJChz2iRCmyP8tYP38qWe+g4/tBtH
BlNV2JmNR9/Y+UR1oG1rwWusJYmx5H3CaSSLj75HXsfCPK7pzhhtwiCGoechHvvdlL8vfFOWojqT
JfNnlOG9Uwnc22p3m02N+w4FQavnIZt+gkiBNpMP808TEYahAlOhcxEoEoFMThnbieQV0fDj/HrT
LnKZ1jiZpGX7W1xgETnQfUtf6cpfyyQ7vCumIDIvuCYSaieZsHU1SNBteIAM+vdpUzctYExwXacH
1RhesAOLUbPCo90qwORNilESKcX0q9dVnpAhB+mDFe7rsGGdXdK8pYMqhbrooUMYc2jyua70h9aT
jri+ejpWUFPXa0DhlWgyXeVqyc1US35Q7coX0fPtKOHq6NZOqVa8FH9UqZFMTXfbZm/K48J6umdN
Uc2xWr5z4PyI/ic5e3zJPKcwVGcw4fgbNP65SesdVYoMPqOAI/aq304Hp1BJ4xRtP9zlV13zrlkc
T8++Sh0hhQPcqSJ6cgf4y7gx8JIszZP7/igr71vRDHPcK96W5POZ4yMGFTDCDpjeanPaalFk6OLC
sKEw/A4sqLM5YBbbm18vhrnNAAYxxuK/gjx+52W2G6nAn89MqUlecFOBG+XvTYssb0BYj3LkxvXg
0osJHoRn7HXqSAzmBZhrJBzQPf6M0KCr6ppzhtxVMSYADhF0ntEoEumSlF6b+z59fhUyvpqVdr4p
ARBT8plZxG3Pb2XIQ63Fm8PHSjIhuLVTEf7FehKKQ/u5pDDltLDOMt/PdodC1uCZJUbhs2Npj6FD
canr9LGewRaoP0oKHbye7uoXYxWg8Y5hoT06ssLoTvAVXyRHjMDczaj/rxknlQ7pIeDu/3AKCVQF
td+0SIywAXSbRF67PEfs0efIR4Jjgb81ctvPj0O2HaSCLtne9XtsnqTMTBpwmswgVOf6QGuYb3q9
AMbvMTmN5nY8pnE+DW2PdRjGGtHTSY3RfeLWy18JAdEqKk0pg5N9o3i/ZnJRZjDsE4/M4d0lDnfN
I2UR48a/MkcvHG9GioHJ6ccBPygJe9G/llGuoNvlaOYvzWFEvWxos30VAKN3gNHOKwBnMD5KtuvV
hwvvG9WOXJasHfG2jdV4T6gCT9ofTqFp6Vg/Aery6wNIO2Kl6hvK9Rh8Rdm6ERiwMdjqbf1vKNwH
Nly72pFj/ikbrieMmVXtuJFl32XAkAROhehmOR+qcOVtDRuEzUwTYbVqmeTu9fnCVhodHybRoF0F
yr3rfcxxHD+9IAqDtygv99/9PhDjy+xveJzV5KsqK6tsP+gUIqckBH5b/0RezqTg25EBELfs6F5s
1xwP0Bx+V8YrWvN8hAcSGj5aDdJAZIf5h7sokk6Pr1LWOeVMKHOF4NlgpcPIeBBLm3GK9wQMLQQL
rbHNh9KtNoH+o/stL8wwaPDYIfsXHzqY37c8iklg+jpPBVv/HSuTq8M8HBsMTNkUTZS8AYuuvFrU
nldO5wTDYwcFUg4ttMsvR72JIOX+LyU/GVu/8rx4t7MQZp0zBnmfK+DRo3CGwv3O6qU5w8CdnZQA
UhoV2bH0wbOs+ln9eW77t+RYg/C6q5iOgffmBZKh4oBfq6qmXtv8oud1OdLjiooqDs8AjaQeaCmD
3HMpiLhBJU1lkxsxLjsjgxti5Kvp4k8zV9Db4kJIe8LiO5ienr3e9gaeiC5247aKSQH/PpdGltLM
DuyJLUoIguO4MBFoMYvcNEgPRVIEM198XoZLi8q5MlOK/Md9jiBfaVfhT8wQt4RcVLfj6Tkg+Ojv
2mExlO4bjD3KH8gaCGjEuO6KN0+Zjmy+oopvBK37ZycxFQKLBe5aZnOzgvotV7PbboQlfsV5FLTG
Hn8Nn2j4fa8ubK3V4uhr7sFDfW0ihYJxyWHjg1cxpHkXFMQRxZhYarYS6HjYZlJW1qZCiUHBdftF
hGT9gpLLQH+rhIePBZ2f8e8pLUSXxr5Gna/2nMwozEwq960YbFOH/k7qa868y3ZS4LfkI9cZmmCJ
++/mxhIbBKFQThgmsKKisQy+xKkCljHDRTfWDLJgtuVROdNKoqiJ/sZau6yAMYrNeMI8FAx3bmJr
D1Har9VfOk6JXf/7vY8D4T9hEw3LNXLJigTM+Asrz81u4JRjzTGKh8HtvS1jowjNJMokRkanOdg4
fql+uoHXhUNcCTcarEcqWzhxfK3Qpz98PCI/Xaa27DUPOLkAvtPpD/c0G9IuS+zcand9ptc+8Yhc
UzbNXiff63aSNEYDZKjEOdvP8QUg1Gr79bLDukTCXblAyp6e3cI+FyQiWZOncVe/dVYpPyHGeNL9
hwXm1rZdqScodQpRhj7R//cD8v7gMnkbi1mYbaU7vH1MPcpvTpdgNC3Yk4QYWiURBneLNy2Rj6ks
JNThhFx6vqP9a98b6yiMyWdLJmlaqTM9Jv361w8osidr0iYcfSwCDe/uIFEL8xf+BriObaO8cnTS
uipFwEQhrU3QBMR5CRhCNfbMjfIO1mNViDbnjJsnCaxq71aK4upCP8g08b7xbfuWPb2VHK0wqCeu
38ANS76A+PI7E47F+pZnFIz3KgN+IhcIy/TwNYvns1RS/azxDNw5NM2MWXTCR61/fA/Kq8kGFUGa
jfaGsqTIOTN1QwVm/yW87eL8O7h5UCMDObgIkDlh3dBzJ9j+no7KIwCAxukoC5nSpyb4PPaDVcDF
GfzA0/IKl4fykqvmtCEg0dZkFFn7Ek98yk9iiNZkXOJSgdBWBN5E7wGAd3aoUuijdkaZ0C+/C5sG
nfXK+qYtrpzTarSM33nBQna0tGiyWemTkigbpc8qJzquAjtugzCQ6kmQg7mlQPp4guIk5jt/n3qa
BCFiNc4ipk8CMChXshzBtqj74H8Ul73EiDBZs3EC6OlOdj+p3Q61xdxLjDAQtAuAc0kXoC8zrBPw
8/8aK07AMwtx6HcQ8R2f9OP1aXrujz/AZMcufz7of6SKWDMtoKLR3QywRII5XgdsCdISw/yWeenw
O/vjJFrsiwFNhVLMNCxPyp4cPDX1N8vnse7Mt0MGMCSrr8aUtrfDpgnwKlLdNd0osofM3Vhzj7zE
8cFQaEpKaJnyLl5ma91MWnfUvFh6bVt+TOc/qHxBkIWqujEng4TNmk7YnX/N/Ln8ydTz4KHJzqOP
/uiVfzseajb0sJ6qNELHUL0pUFbL8UWw0NmKv+4Lcwp35TI4dax19pJImT7GSaUw+ne/zo27GPX5
ZL8QoIybawJWGEJOQlWOGOfnR2mYdS0/XQzkqWMbHypKJZwjS9XVFmM5jJeFkVxruIAe9B4OauNl
vwEj/niAZYmUzBj41TjaHzDk0Zr6E9bjZHuQc0StlDcNVWO4c2k/Qez2NSvAkrq5Ln3VhNTL30p6
7BVX6/NMEqv0Yu21IEYZNbJBH0VFlMSSoTleqFl++ZwHzEmkwNO9Zds5Qi1HTQTsvajIM7Nqoqhc
bR1S/jeDOH5DrGnKKPVNQ1wuj0K/SbNe1hUEn34H6+Sx5V8jHg+567oLk1VX4r7pCojLDfGU9ber
yuYarn5f4FSho8tdT+C83Zf2+UjDVcwhh3ijzJhI5ZbB5lVEylpdOjieymx3+BPHq3LX64FlCfZB
6d/m8EvthnViDeKNn6Pfr82gLy2ACH0GYIHEuqhUqbUTl3d9dO4xXnMQDxh1tdRrj1ad985McSNb
Bb3nEBlrA/HXisg8t+4OCHgBq4VhUucOlmPHHxER2lgUjjs/ljAgzDWS9xHJc1GH3nfQiEss0YZD
wQfQELkPhWk5w7gDu5Z1QlmZ0NOHaMmECS0VYFJsScB/h9OIQnQtndYy5vYJLnBXLjk1s2hmbrh5
Jr5wjbXG9hrKbJ22CzxZVYWqR0ut9N/EhzI1+VgoHNWoXHdB8qHe7CxQqDwa2shd55woMesksoOH
lX3r7Av/95pSOsfAF8M8UsjZtJh34NJKIM/i35bGdz68wjZjFS1OF6Kzht9NahSt9Lqb25Ov7nN9
78ZCmkHJfS4sjknPrKiSSN/1GcV77l4UV3UYjHnUtEEXE/8qMUiHggTFaDsrBRqyfSjbqm+kVncl
tBTJFmp1pPIiCJvCFV67CynhDFiAB2JrbEVEzXAU9SHkwIOoQ6EnTd+RpMSz9FHrsPTo1X1Kgdzl
BKRm8IyeR39mU9x6JYci1Wral4wokWg10GfyJ1WP0P7g+zFoCzXuSUjHD60Z91ADVXnQGh+V2n+4
nBdGsF/OEfV0sco4t4KLdUZZM9v89788FhkoP9j0MAKPrpT3Da4pCrgMJnzb1KmEnP7ZvuN0oanC
Q34bCgstSuHCJIDpwWizm7JEsYIs3IYCsr64wzwvkrZWu3bPNoGlt7meZCCAhhabub8N/bg78FTT
vN2PmyIn/sIj8hfoOB4sVlOThfUYi1uiwGsCau7OFCTK1I35x16yEC1+jR9KVe+bzVwsClgrrJqw
fC611sDVy+0D4iQisYXdBlxo2BHRVn7kwmuM+xZyM4vQsYvHKg4kNyx6A+bV4tmyPQ2qXwAylF5K
kxZIbS6AstUNdGat3wYcCxoLtbUyrj8EsIt9Dy80bRsj+65gi2zKrNzEuCGFx+oibPniDKhx+Miq
VLoK1S2EFHNS44c+og9smmrMDwktGUyvmG5SE+h6yAnz5PbX5wl2y5/0c9BJss0BRaFnfWVBwmnh
uw+W/1t9YGB9cfPUdWmjQZlHyRZ7fNb7tgA6lTE7fs/s4ek1mYHcu2LLZ3GzoNzsfT6ooRGVYHbU
YW3AfIGIgZUB+bhUlptsfX6p60GiM9um0uTG0ueZ9LZ6LzTVVvcebxW4KuRsfuDBsG0IXwvzCRaW
6qNZPQO446i535qJ517BvIxGbUNyvheiym1izQAzGbSrRStErtjTRJbeTaQ5negfm0tBAnV4UGfJ
pOgYcAziWj50g7UIm4zMHAomxRl8azyl5rl3H0F0VfWWmQeO8lYQtrb2p3+RMwqslcMyV00xopXt
DWFZa/Fe7r7Pe4xytbu/6iziZD8uU1cOVsjhqDpsL9h3AABHGPj/+D8AbHx/Nl4UpPwqKgfzy/ha
RT86aHRSJRcvNix6DsZiAOT99S/gLijh0TsTwxJKONld6NOTxAnCkh9yzMv86pP3sQ6hCCIu5bWs
v1nbCwWszs5BqjI/PNrypeCN5mtcKdzm/Z1moc+9cuHi0OOzL5iKwZaxRThCQ9PJPMdhO2A6TnTO
gXELtOgaiEDL4gSJLykH7+AxqAS0XgpEwXW1BXfEEnR0cAnM4RcoEUVqqzyIDdxnLHBUjaXGjeTT
uCFagB11uqOqhFjIbPWk/deM1aZZBXk+g38TOAbGySFe3Od+Kjj9eUSKxoDcQuPcgeOPrp8lUTwB
LqTk7/CJYktCnoJVqGIhCeKOd52ToPsTrRxwSNoHM0P1YfXb82MkTCT+0jwJ/daMkC5QvHWr5Gld
tswolZKzT3G3ixtGFpv1Zvu7Xyz4QC6RuXcEsIeDNr0Iv65Ir8SgfFSl8H8KIvNOLrH5zMhRiIBA
TE6SDMuLfrdlZqaHE2KVXKd2/xycR2zxqkD+KzkKf6gk12jEqCENU3dOzCPlgzEaUIPWNx8eNwTN
TfbBb/Kg4XO40T17G+YQ/7XqKdWE9kc5o0mjTcQkIgFrvnz14nwJfqAjQ/SrmcoGzO7s2Or5GJIL
OaNR0jUwx/IwjoV91lEi+nCgMIUaMhE4JtRnucT+N9Qdv24jA7FCMKgT75hC14f3PqvReRBWgfqv
pjcTyobAqp5vM+MZHX2ccOpawQknjDNsNlGyfHI5Q2UL9sZ/HKV7Fd1SnYCjdQ66UeGXuWvxPEUM
DSH7w28lULQhaOonmL49QEKNxAy2eMeNUqenHgvPBHLuUIrs6IPeHIueT2p+bs957SOEnQ6Rxbzy
u5r8pvOGfdmb14ty029sPaNBGb6WncKSmuqG0FJioUh11A4DScIwXzFHuw/DF8NJMdv99Uv270e6
dMXeiXVV55J2vtZax8CWAJSJOR1F0ZYo42IryTsqAzOSt8JJvW8dm+dmfEm3fsMVkcSDrURRyV7u
oSZw0fIMCuj5PY1xFka6btBgXpm+3o/XQVecOZZMt1sQUllPqj4O4YOUKIgo5g7saEEJX7DLqg8t
ocyVLDbFZo9ie6QHvNIapIrw7Se7KFKXOPTUMFRd1uayne5xyb0UM/TIwDxLYd9pDEpkck+VYIS/
t+7ylUdig7O37aRslhc5RMxNe+JYv8N42VZesmMQXjxOBMvgAXGrHoZjsAjF7RN5NK8AXoS1UTZV
6zjDh4v4Kr67PAiGWWsOAf0/ETb/mUbMEO3rlV+0hXu/3P/aQmtisu2EbxRs740vMOIaJIYNtcG5
/563KmbjijLUd6Gmpet20VFwF/RcqHWy8LH2cqbHdXQSnbuUHmxwji5ZCItqkxxXbU+LtxGU9snJ
yixNnL2YcnBnM8SZonSKxmV/hfQwBCl8aJNCrNUtQ3CoiUJakdJ2+4V8LafU6wmEj0Vzwv857T4L
uSYLtx+jg4L0CsKkfJoHK9nUvC2adsgY/zSx5rcmRhwFtWtaeHdO1E7ZZ7mrus5ZhZZwhtzooENs
TrQaHYkMCLbFcMd8zxUt82Ced+R2ji9i8kblcGVWr+Rc5GyykvdfU9MhW5FXafU/g99PpKsLlOYc
+AmBrT6fTYh9X0wXw73/cGeoS19/UQVLnZYqG8/vI8qle6VOekFK65DGP8hbWQHrzgUiK0Xne+8h
VJNeNlT+7sDOz2uPvbVkiR6wLGV9jF7f3waK53FmKlWGobyqGWqo1138VNd6ixan26I8S8U6ot/5
xRavgkqbYIhPP28Jhgx++lpUzqtaRXuzrxgRIAwNVloYsMA1YmmOelmED1DtULPxByCHECDpPND7
PwFx1Rc3JIcUhDlxy76Jef/XFZaAFpIAjEMJZLeLynpte8eEnYxxvUbiwRd3u/cB7yZ9RqI3Y00Q
g1IyMYBL+2+i3fd0XqzKyR1tgI0sIQTqZeAjl8B2zWld6ua+SurqbY8ebgfblSQbPER0CdMOi8Df
XF5BZglEIUVIq4L7XNac1/+ShRw6tQ9UYMFxu1tcIvkZf8focK912uLpMlKoRX2OUxQSFWg3gIE7
B699IVReSBoPbFjbueEYQMGVrAFHWfL/xoShJxxC+RACIIklKclzqN1fhAHtDaTe4I6wJMz3A9GC
pJlQWR12lrAZPFMdkuRK78jdd6kgUOVOEsorktRw0G7Ot0WefjENiBkSSgyilNraaXhqVU1ysgpR
HmEBu8IOM9jfHGM9YO7KogZvnoYvRk7GTl3mBnj0WO6pxgXnDUt/NZXOUttH7JL+1XTuxlKujuKU
5fyBsHz42DjZ4Umm46stfPMdyJuW3UGpqw1iGgn9ulbzK6/0uhVD98QTb+AHQWFMB63vRej8xR1y
dxdfFrgaT2d5cfGmbWKFmxu4bty483sUXM6sp4YeKrVHTJv+lYXS/oO3dqwzITbQi3l93gVhFmWn
CMI0XV3o37PcqtK7ZpthSj2YJn4roOxrdjFPRoSNNeBiV4vK+G9PAKkM+CbHjHGAANP63XrLo7KE
mYs0sbYBA0zKlANlCLOIjV13HIjr6igMpIgYwc6K4WUg7Bkj0I21mp4HOzqO3tWxPk9obtFfyCkj
pNuXLftnCjjFoMQRGo9gf1bTyUvEmJU3I72f4xQINAXevXe4NxT1tdfvfuo/1IjfIQyZKZbz7Kwk
cXiMGWQ+hBOWxSZnuMrsB2nyuhG9L+0hlny+6jGe1cGDE86yA08b5w8P3YA4NuLkLxmBRsO5G4Hj
Lfxv/RWvqiFjmo7HBxgJNIZ8dYtO6phwZkpz5+WBPp1oovuhbGp9efZhotNauB/Jl/WIqIr6BMVF
J6lUSbaS8bbxAxYZxBiaNrea5D8nwNgIthDFpwE4IbV1jF+lOFmuskOiFPemy0W0pGHGhyLp/GtM
gzZUbx+qDfYNQzDuozGvy+F9EOqD/F/LmCBfZ6R/Fdsf1HdZlzGTruN/vLxOkOujRwjidlFEtMzC
kUi1NqOsJiJpE2reG5UPE4OH/uDMK0CShS275vR/bIQhCvbkMh5nkNdOTIHb64LmNUvy9KnQaX2W
QjTWHWnHCzTZjTK8iRH8fhb/ChCaLVtirQ4wReD26gqMgQ3/nVC0VWO5K5hS/HBJ1BaZBncGfWDx
8mnbjeqHZFgwGYUcDUJDhxbQ8GuugrJHG4zBvH/TLjPslnEW9G074relcgvT2tIBruRKPt21bk+s
k+iOAVNHuBkF14VblN6eEKYJdYXHeca7o2EK2m8hn4Qqc2a/fji6UDt2PMGtGNESQOlrd9Nrxff3
x0AQSdkVsCUvtMJLoW6ei/QR+X20kdCBCOChFGQWFupVVGu0Hl0mH/Bl/adlWnmK5xIesAeGbIrS
lJHlLoYefgI9SuHilIi+nXtsryPCc+4MfZXRFTkD+DzkpUQlChNMtTZkP1Dc+fI3oXJBztCQcl6z
xIauQ0Vv8KCaMBWd80wbH/0yPrSptjKBUXDCGNvZ3uTr8OMR/l5WXXy5b+RSLLASTYWqhtdzubyf
KoIeYi2FpVY5nQi7KCYng/rUcLwwtlyr8jgk7x9lThlAyo1nqzbbJcrsbhMLdR1xZdeCT/T4iYDm
kPuqO4gxEzuanHIquCeJw4svDiav0D+CWhxw5dSD/feC0HeiQrLAixGIhcCtACfDydfWpSM7LbsJ
1sv0xB4W7Seia4dSI+idkCBA4W+i8O6w3KP6Qy+8wst/vfLS/I0WWBRSBT7PLXh6KOPqsfGqF5EC
Ek2oUKpvgpd58G5w5VINiw5l1prV17kRGvVg91MZPefi1P96HKdYhyhsGOFhu1qfgoysbROo0NeU
xgSpzPyay2icWECr+NbmCf0uxzaFZj/OwEas1GCgyEkjnbAoNOOd6A7Qb3N9gRTODx7LNWJw0BmL
5JjTu2MSdAXlZtRTn2SnTSjWa9KS1kZ6ullYrUKX8IFk9NbG78VV0LXqEnqCWqj11xeKFBj9NAi+
sfS8TLFgSPxojPvjPpC5IT8ECkwsU/bF48B8JBdR/HVgycXRvohDgWN69qKuc/RV6Aomrv6ocSFP
xWcNucvG8hk3WJb3MKIUL/Mdu7aMxfG9mNT3YAujeQlrmuughfCBUWyW1OoBZLfCxkA1ilRE7A9V
2FgRtCwqbJGFz7Iu6VTmZgU6SwIG/RshDZ/sBQS2ZOW4ypCzSBJfCuF2F0Iv9sE0q/RSmqc9x1QI
84nvGBsx9C878ljgx4vCuz/6lq9M7wyyRVxW09AVl1p64AknuiHQL+R+kLbgQ+IHN7QYxsOmgca3
sYFh/Zfe7j+yWkOl2QR5yfDGueas+3+p0TGcGLIEFmomxY1DgStlGr8DWFc7wRTmgSaKiYY5qtE3
SsVvllkVwWStQ8WfnarIMHpaBVQ3kY7DaaJuEeg1y2O0I3vAdUfsPOIL8V/StY5ExKEoXkVJJUIK
CKYHgTVnubrqkPS72Mzk6WVe/aEmWOoLZR6Qs3Z3EXfTgup+3g9EoRS93MRHkbYrnaw9+X1MlyNb
5qKNa8tSUC2m7f21azPgE/0wtczFRh/OXSX7kU87i3rPsHv7VgTTRhYujL6ycDrby0ftH+LSIlbw
KSn05fCY7Bv8KRuURqL01tk7Egq0P+i5R4I7bGC0xMNTxxwGcN9PMGvlh5zeL+nTSlzYeQa28eUR
myrLSsSiTsIIU9CI6XokUeWk9cP1BprfwKR1lxxnrK4GzZHNuEGsnW+3CMrjArqj+OWBNelOE2Va
j9SL9NN73tyNski9SqVDjJgITo3lurhMmDv8GEkVZBEH86J7E7N9NHqEHPUuqGif/9SFsvgQUfJn
S2uCCTpa/Am9WQTKXObOGSvqB8I/Ap6Ko/O8rB9d9xlJ817bgW+tXA8PpHES8h+Wi2FNbVoJDHz7
nhq3PawjFDQe/DOHgybPOmq4F1rOQh7wk9XPOzJrwirRPfXnNPkeK55FT47BaGIOPH99nhx8Rd36
L8DLNc6CPSfEdvN160/rA7NnBTgy/9CMODUqeBLkwLd7eHBkO1IXZDBJKMTMz8LQyPKbXKXByaer
9PQ9sdMqeGdwTTDKCRSy/s/3hyLGkYfPir8xqDv2MaYYnTgoRHo3r0XEC9ctnSLeh56RY1NLYiV/
tYigXG8pPeZ4pZZIgakG8vj33c+In82Jp/dvfaGqnedYyL55kfORI4SGckZn0pQ17cKwbX8YNu+k
v26fYPcQKWuuRmIDqn2FfyAlXg/yW1rTKJ/JJeg3lHXzo56pKBM3xtyyE3cw0wUvAd9RK8LiW3Pw
lgWeeQ4D6I2Jvvni9tzYv0VrY9Raoa/aKUYSRMIXjQNjzb3gf222NyhNUF+SZDtgM44lZAjCzul/
7VG4faGrLafc0fkg9V9mqm/Vae5LzB5dS7N0rN7aNtYd5f3AsF9aVeHoQ6Atmd4W6MH8tj46LvY4
NG91PUve/IAvgmSMEHbWdXtnupZ0bJqE2WGBzHOk1QE0xwoO/ocisWiCzPn9OYuFYgf4rE+9CEKu
cgCFcHVKaxc0iZBYOgovuGb+GFjYX293Pt6BtMPoAbHF5L1du3zfn/HCHekl/J7AcjYH1r1efdlg
gc5pEtJJmBDnv/0bClfLachqPXayDfOo5ZcLO6xm9AJn/Kj2jIuXxi9qNN1elQ6vEcinjum59keu
uE9IXIL54yMbyE0qfjmnW5P2Nr2CAtBKZASkI+HV3jQ9N9erpnf6dIMkiORBjS+rdImCR8B7dSD3
9Xqov98pF9/+wwpFi6pYPMC1+1BcD1XTnPxcRa2PYVo4gHOPXEcGsKb8dZkRjLwzixmbLfmEjKbU
77LFerxPckLlGXw3DmbWf83guLv9EV7H/ko8/bcJXHKUrEqHffAM0MtYAUlN6b0glaA89OtnulOP
JhoRiB0r9QDSCTAxdpdlJ18eyTDZr+S/vGjEDMle6vkRng4ntYiJl3kIaIq3kYKEd5+9ij/OLWlc
nHAcy9gUNedl9J/gRVe3s7Ck1CukCihBO266lXjz5S9I0WbQ4mBtE4tue8CxEbYK1M7AekG1oYnU
TBULJFlJUbgY+gk2eMKXbzt48aVvf68/RAmEpwRgOvytaKiGwJKk3pyWrCo02y51kNZI6gKzbw5U
jZeLu7WwvigrC4REk/x0NdvsSV0UsCoA2QKfOjTwr/5QrVLMG14Amtn67MmruUloUmlM7K977EV3
RH5QA2jBk/9IiN2SkApJo1JB5cFvKEOUY2/02o6jjMzq7l/EQELRoS+SV64a861ZREfQdy+SoKOx
dmt1wdzjLOWFk0QuOnyMRbhgqW0MGqoo4oNPmxx3rQwhUHj+WhLcfc9QJdZFnlEyh4kmA67zhWhh
E8jBlf0XWz5Ife2NI75/YZicwXI9wqLXh6t3nX9hcyXtDMdaPqZfiR7iGtmQAybYwP0UZc0TT80x
14Fb9/aZk6D9EHvELGkj/wjr7XO6GEJbmonZ7MjdGOM96eiQ1dZzYmtpMUd083Zg1n/7EgdaynY+
WL268seq+uhpx1tkVvA/L1Si18qbmIr7bPXtuunmTKyjEQoZ+HNI2zON5cdewhrGhdb+nU7plRuq
4/Iw5aAhHzH3UA3X/PlU9/a7MAGN7JQLaCr5/d0cGmYRFT1wa85Q5UF+p342vsgXzawg71ttX4U9
cyJrULbPFQ+0pfnFW62Eyw7pCOzjDemaf9msQqSc5Lq6TSTJEIL89ohDa4fGolS3hzm0hN9oaHX9
MskXIF5kSk4hvcxgmXDqS24xy3D7HpHxwXBcC7kzD6/EfuLWo6nyokB/qQGpa8Tp7t2zlnmQp6r5
/i9e9dbXL22TbN9e3VNvmQwFZCIPT3Ixdx7ToI3HG+BHGs2/d4AQKk2W6/+cBshVTB+54OI7WUnb
p2pnoHDDkD0AqBsTEnLNVjQbqPLqdeYekaLA/8+mVGacObyxh62/Z7nPKdGpJe3Ey/Eyf+dt1383
fYpZu2WNsc0aCo2t6Q1gw39gXTiBajEowOiP004sc0eIizuZ4YB1QxOGg/2vORZ/DH3U2rLNEzzX
GT7OWZpAj/XowpieI2mIlTl2UTtPRHVfY23/X10INekclGQdm5eabMAq/aPa0uG0AVpI8EDQVUG3
hVBMisVDcUHUUAjhbMScEpbMZQ0xDt0pZquk/AAFDu44wnAHt0Le64EScYyIZmwAZtRCffY7i6FA
h0WuscaXdSArA4zKraWy5bIBgFlnECh2YJkVybg7A6NXhWfrNoQEA7196gurHBsyrmoC/nQqAh8p
avmRUB08GIuLquIGQs18aNVSKblynYvj4wEJrq8LV7DbiYZ3bbl4xtkJhNxa+M1SvOkKCqL8FFR6
ZD0KORsCy1bG9kL2qLzrBVVfzVN6iNnePL0isE8UX1QKujGIdHdxDFjPRnPVxHfbcK2Y7Otg79vp
QOFsbRHNe0+8nUo3xGy38cXUxGGQVc/s0CqUrY3FkcbJxynr/hFKywRzmOC7vSmC7oNO4CCAk4UQ
vS1lTHMzElXDgflRe/qrgQsjzwianSqMLdF+GPnpaiUW/9oDU9vs5MSvIxuE7efsQ4Gr20qg/Ru1
uKD4+n97YGDjooibJOOvkEpfDirSrlDCQ+/INKgXu040LnOK/2alAF2i/RpYUX0sA7K8hmdwlM2d
GUXC7Kpt9E7xCx28cvlv4SOut5IGp5bl9V158TDdTxcAevoBXS4Qv3D6H9oxKS5vey7lI7LgwKVE
Bu7zAHhlm2xu3DK3JTcHf6Goi6O+Ti2MCelOBiL50vV00NDnNR6d8uaoq3HrPtJNb4c3iyt4WClf
mv5lk5H95yilWZvJCdR1ZAstJifsQ5Q7ye1awkNidxzc4dAyfErqtaMxt4FMsMPzalc1tGD32aOS
KUXx2A7SUoaDAordrZyzmAv3qjpgA385rK5DudEeR3PFARBftQD3oc5fU10lIc7tTf0gz3ZDRwBf
kJVv3ip/CUnejx+eUObdeEroZqE361csH4CSZTekHcpidUAv09bWKNNZBFoZDHDv2FPULavGgPE5
TBORE+M37LYiquKzgZCdb/l1DjQZ6VnJ6WucH5MaQUuyphZcbY/u2baMUizodtSNR0phKFnr+DZg
WmcefY7u+uy3er0r60btn9vfsVEr7NQNVc68s8/Cb8d+HZxCUTPi9iwDXFdg5tiE8a7BNtD8J7i8
5c4XHcI3er3NpcUVVQrPUD9WppGz0xfidgg97vR7UTaxFrhHZID+86xT6x7E1Qc1ucl1hVOyfvpY
3w/iZwwJ1buJ/hi9yap6DhDLSdqv8wSGJUOhj5pSewIIXbusi275aNI1hb/2RYVesM7DtCSXVikM
UiGNz8XdvhfoR+fypM0I3KVypaBvPn7jP/5xBll8yEKqPaFNrlFTvmNMInmJcIOgU8K8Dp0CZueH
M9eLRdZa1O6pEaimB3JIFW+qncwMzGWFKAHM+h5sBB/pgXMo0WwHKr+vJb1ygKSO7QW5eZb/MTOl
2VK4e6mS6M3mv/ywX+WTOFfbBNpZgXoNdPPY+zyD7pFxcJO25eF3cTBbVGVWAwxxf2kEwR5j9y1/
oiV2bQfX03zX27q+jH0AgtEKrtoittoTDAejPkyq4zyRS6mHoDo3Q6M+MyuLYaNF/1ksei30PLjw
Crevme5cLbfX5V3HL0uwCZ0oXA9MhhFZxbEinO2vyebz8+Vq3ieOlnLX2+HE/u4fqzmZIZ2XhIe1
k96tpPJk4DcJbNuGtc5KCOM8qS4/gjtsXb5ztFLUi3jpoRYfOEmfYiZkjsw39vn4/CvXhPesGLbG
xUK5WUA9DIEhR0ecG8PjOuKqq8ID5G+8APPC/T3VX7QMLKTmxMyJulG/7zv4caCBpXMd9L4hxfrw
QSQsLcTKexN/ZFS6kJR/w49BW972SwT5J/KuyjbXK53S81ELh8H4m2gQ2zAoY5lfDA3tzZGNSJdB
J0Jt7zSlzs+XapsUL/AhTYR2EHKVb3CJYTOjufZuFNmxdd9DKDMSMW9medBUbm5fH/9HTDxx2GTq
gCmvRk8IY++Nu2UC7POG+ZeWh0GodnjMG5zgw+kIiD/USJ9jbdiQ3fpFS1o89Nwzgcx33R0KhaXc
9AKgG7buUNVd7PGFagOnJNH9VUL4iwA9Pl5LKyhBJ0cfJEgUF0YncaWp+0KSvBWLq3soo022vX77
GLvfJHRL0YJ05h2AmVdAKMKPzELaVszP8k5uLf7dwq/ZPGnqTPYTPtUU+kpN6lsojt8YssZuO4H+
AOPnyaSZTtIphLheh1YY8r/0VIVJAlHwC+ITISMGTBVUm2s2hUq2QvczA0JaGQH60GGUuLFvt152
z8tW2pvHASCOJMmb7iH27NKlazTNAiL0frxyzmDFYqeY4lbmqOlh+6ev9M0zDLhTvNkAVHgEWVTr
+Guyln0HekOTVSL2NHNdfyt3S2fudJTT4Qz0npKLm9r01KeKHs06uAOiTW+nHTOCeEyeQROPO/Xu
1a1XHkxqfuaYiIVAhSVs4HjeAP7oZ1vXrLak6prGy30ZDGuq0GKumM2c8Ses+n5yTT/RE157JXUL
aqbykZqGh3DJSmo8sf0xYnff2lLg9q6sFqhx+6LkUZVXk/rjzvt63lUJHI8Tm2VrGtP5s9CRwMdo
mZxxKIJySgTHyD1Kyascrkcj1IF3hL4eAWO+RZljZu1vEMz8cDAb3j4FqE0SLS/Ae2UDn3C4sRZz
X8ofu+VQBqDi+wo3DJE39O1/SIWZuLYKDVuzJgHdH+x1aOQ2UpG56wx/+KbEcTA+pw+n5/VAOvDi
cI0dsfD8twC2N7m7/E0cVNix6RxWYRF3GWm8iIm2lmedqhpHyKrHzzowEo/TSkWVTxwkKDh0uf95
CKo2trZJALCZtVGzl+3ZpMiKF6F22w+IA4DqIuVhDP724ItjATVZUlHb8BwBxgskn6YMtpUBQNOT
lLQ5ZBFY6w9azeFXyPhsoHkzC06HeTpggDE4v78QLfpwiHuXqcJGMELwm9wL/esIxiyjfQ+n1vPO
FGdPoo0irn2XuK7jrryzsiNUOfF0Y7cRyQanqU8IEMkVkcyFLRJ68k5vFX4GyFJCcyVLLT5eWUvS
xnoZ4MSQvGO7H3+nDImOGWq3SA6Su4XpewnxJk1+MeulctJrcXbR2pzaYpzYwGrxciEuv2MXr+ti
KDALhBl2dKnH86vamZxnmhELfx7PxryVjcp7cSz0XTif8zYBdI9+dYYTt0xl8+hgHUjYYNL7NHG4
hM4vB60o2zzIq6M1Px/Pn28KXHnm93IOhKY5mDQPpnp9gFRmIM6i3gDZm1p+CwOlxzQwOs+D36AV
x4lHN9TbYfMmervzDioCNKfZXTqliyGF6Pzi8cqgOFafPurbcCj8c66e0//phLNU7bQNdQ2EDBG+
CtHjE7xddQB/vqcWJCZBJuRoFsbJ8GcMCnh6r3YEuYGIqCXhbMveOkugOOblgbkJa6Ab55kQlUhu
JcSYKGCMuHdYCiqfRl+BfMOP2xPuO0hKGfGbaw1pTKInvJeTkEfmqtvt3Moc1TE2uOcAeTFzBKGM
UtMigecP9RA44cU+uMFiHmp+/PcbiKsumhzlMBanrns0/9w/vs+RD9VlQZE7bmhytZiBSedYUJAx
vUWHMbLH2Izh8Oz3KlOA7waH8pAaXF6ZoE0d41REQyCOyDjpCfhIQwTfsw7Gc93LqMEhtF7R3OwN
F3KU/0fugBJPj98endn/O1oKFtY51MMP8wpRsIO5dtiHr6FxKQkxwJmU+3DKsPhI2x9/nsX52mZb
XHXU6BQ1JS2tWcKx4KjTmY8wpxLIViOZ+3IzwpGoRH0v6J1Jyj3Oy1n1UlimmFdW4EM1Q9u0nN9w
wmj1n3PTRJS3tfIL5Z17bdUQLRbQKoUb840Y31ioZVQaNHyqpQu0cVo0g/7ZH7HryuawMuW2Av+6
5V/5QYUEkHCjRITDnSJM/0IvWhJhC40r0pYriQuS3pSnTNbFIrOJwxBK7leKSUU12ewmwyKSIBD8
vl03Bjd2klfihgt4vBXetIMdn1D+v9lpIM+Px1AtebgFEqikI6Bwp1t3i6m6ByR1PP6ioA7yEquk
O31WfjcckwvbEfyhgbOG2oZfKtpfeJRqc3FwXGFsxhJ0XWm+h/F+YmYE+OsDR+xdraxKvCtCE8n8
d1GS1skesJzd+VG3fn2EHx51wLYejEyqy4HwU0CEs552OmHftVAQfXDZESZ/YdnDGiIYr6+X+g1S
mRD0I3ZQuHofr5nkhfvMmImc2aiSRV1/SVruZ6rmhSLgcbiZkHia9T4iy1YCNk8nqiLsIWkPXWtW
j74NvRdTft57FQUtXZ1J4g944qU7+JnsYRmD+zfLthtblBtBMfYkZNEWcM/gT/Hp2qSHYvh+AlRY
B2guouBxP1yjR+SME3fdm/lEr3tSpYof/xlEVvBYF/69MfIykl8VNadXSYF/wPIo40EdcBdeZRhv
2POdwnLDtMa2NRwAEKKqzS92FQH5b+WeEMubY8Rra+HDr8nwFXcqlBAhgpbYQrp533RpenCs7m24
WGekpfyiCJBrGkBg57DY8LGqxYhCwMWRn1S+aXMGuUnmwLL94YxKxevuiHQPTP3fXTIo1B0E3aU/
GJ92cm5XiKosMlO2M6tpt6zGRBuvAURe7PQy8nPioy8/ik6sQPif4p8ias/kIPFF20B0PXXwtvBx
oaj48Cep4z7uJ1i+MBT5UP5OwG/wuBGQ6CzTkja+9SgdDUBoI2KOM7/SQa9+chGJwP4E5pViLw1t
UoSF6bXOr9En3PRND1BCKd9moi6QoH8dqwOGVNlLfKM7oGhwOLRMT3fHtwLngi7PpoQeXYfdEnn/
IpE8I215M+aAmGdbgqLqSMjdi9Cxnj/8Fwk+gDisPxOlDaIYDmZ95avJsd4QWgJ5euQRQ/MuqmA+
tFSUpw2j4ucxzzOyk5bsm/BwCKOQ/4tieyNsRl0bNOp7AKlKtY22jTINCZSfgXY0QzhAkXO5K0u9
9V7lYCwBLebM534mL/qNhzO+xBit20ZM+vlcVdlHo26+3TuARMcUDW4lbB3kR9k+Bf8UL0A51Z6n
EKAz2FzXjY0PgggDDfheyKm0PiqnDpV2b3yz2aZBG0pCRoaJS30llvs+K/txo13TBzBDDzkkzuEt
A7bAfbtZu06B5HMmge3mtRes9DzI0t77q0N6OulbyU0B7Bwck3z1Fx+Xnvu0mU3NA1EktdI9y+2i
ppF/u7l8hOXF9LzLiWgtrFvQ+f8htaSvzuYe0AS3xuG5nKc3/xLdtaP8zH7Ke/g442Y4gcBpfwmG
VxRbMjfdvJUv0pGuGSRKrdyQjZqy6ZLkY7zM7z8xCnLI46YCtqKnpbrwePHI2IxY7yJJ5mQRvPMI
/Q30EiwUJtyjigFkVAj/wHKiwiZoO269XAD1SR6JNR049dfCRn8wY4VsvjHJXWgybSfAJpArokzf
/zlmwFgSiosH4PYXEw3qtkQAJeQKuS/likrKMP+V3yiUTxqX83D2RnBQgVSxI8VnSMO1/JpnVWDE
PLc2RSDpOl4KqSwQaGHPKnCpeRkuVBH30rjokqlhZ/EX7E1PU7X3NbAE2rU9aSrVPIz8HmOPcozw
7OJJSFKvKUJ5OhmJtKj+/0pK8zxiRlyvUxmfDGdzjB0T7m+0OFf1eA3fMgKMAam9lJgeAbjgP14H
fr4thqeniX5rYbIDZaR2Q+AeSlBHc3vt9zT+VdNn1GSA7Xhi7d16DvD9HQHZqhnZrodOzSfdxJzl
Uo8/OpIJs19RoZ93R5YgAnAhJurlHAXsR763Nhkb7hIeGcHKKaE+3Ge9I2Abh4dxiVaRg/Msiicc
ypqQBJdks/NsnBQeveMyVdKtXagRtujUp+f+mmeziGqbqgzVArKbc9JWYPyT+C9dFa1+w5Vfd/m8
Awucf1L6FoRUHrDjAKOZu8HZ7tNcA3fXXrQl7MN4ImyFeB2z61bgkB5mmwo/VvNmz16YeIUQQGL/
+6wUoAojTTxAmqZW+PZnbIT9JyHbhZf/suwDi2eRXQSkv5201ooglU7qaRMJEUbczYOhtkQIdmIA
p46Gsg40/Sz9gfqUknQAJTW9c3EtIOzCXwiMNSN2tUFvXwJ4cdYKuFJ4lo8+z/ExHq9es2Shrx4r
/+LkFyX+dBf90+wm9dsc/Izy7CTDH9a7lTIDRSCslRPQeumkipkv5e1pj0/xURDjaTGj8N91nDtm
1Q57F5xZ/V8eKatEAbMdxhLp1+h6/HeK/ly/UFxI8r5HmdhUVNV5ODszYV01E6UUW8Gx3TOxOBw2
CoxcIR0oSb8siUG0Wn1LkOhQdqCF1OGCnpnYwKrX88X1EKKA2a1E/PQVNeXWQJ3EanYeUICnLZU/
48eLiYJ7Q10mpO+6j1xWGORyBNfiL8tvcAY94z14a/SVOEAtxxoQtbErTbdGER/cxWHrKKJjPn0J
6JRHHp7m2Qbzh942Rbd0NmKW24YAr5R/ilMGNXU8qB5F/0ieuLkm30HskZZe4iFr1EIB0VuRiX7P
+VqI2jvGBkRKC7G2Qian5s+EuNn0j1d6H0Rhtlzj8Z/csYWp2B0pgAoNo4ZYR5gSU+Tkx4Y99GaF
4vgFFqWbCC5/9T/mPSZuTfJqiV8L8uqrDmy/Cvl7IELpMQkGgyOyCpJogGos1p3B6GGtqeVprLuY
bGwLbsxPRTBHmezQ1vrKBAnLfnxtxc8dAkZBQOG8JviMLiT7m/0Sjtk0LBpA9uW3SXScQpVO1zKO
saezuER4SOwXIqQkvhXJgPwxbHvU2T+Ph5ICxuODg568Zv6Eh5elwc+4zhVU8q3F23lLMAcK3fTp
WnUGXom4NBPm0+s2N3eTXcAKB4CXSrd4MPfGpTJFWzDlqHJr7nL20mEVnoPE8utJJ0GNPaMKFuYO
SzodxNpVZDZ25xDAcXPq4Ooa38l8M9PQ2J2sIQ0t6O56xh+KAdReZJVjVAwvIa7R/fPh6zPlRY6b
8uuEvqBQeAeZTW6KiXmukwU9maX0EBW7qk141+oJkXVuS1nHuEFpJlEst2ryKOPwbrQrQ4qCl0II
8/igUVfYmqHh483G2PlAUkROrEAkU4WhKsFYgSca+X1to6m0Po3uLnxaHiH0A0m5yRcMAPkuRYWo
SU/qulTKhGsl23YobqTE5744zWIH5PQ1M/0BFK9F3gJK/5Ft8bZIZYtq+g16QaNNx0qbm4+Fpv/w
ZyJvK66s956qLwgMnsiaOjRBu1WAewGb0X0BQd/qlsXzMMUP436G7Z8GY0oEsmhugqcq6QbmMj49
6IfU26NTKT4WTKb4B2AvfIycVf8qp+Nc38U+ur6700dmi0U61tTask588jydILfStb2VVW4p4ONq
7Th9UJJwiwRvbR9xvBxq9IwOg24sKRGB99ghC4V6/VE9I5hf5dfYx/GWL/rdvwz/3fPi9qt+/3sg
MvIcx8LUL10glN4ZNnicfibCgxjw0aqYzLnB6nFJZw72GO9JQXyVUg2aZOcHrwfUQL2kP6aIfmEG
+8uxQIcZgDAI5k2D3XhuVHtF8/h/9SD0zplAtpqk2WsOKyKiSRTYFVLPJNQnZf+03iBweQ8fMdyP
eMKv4UJpbl/vt8hWGGpVWwNWzTjRTMHGvCsyGEDgk6DzY01bfvAhP+9s3p205kOUkQ+gkZIYeW4x
LhbleA7jioIKrVZ6TdZbPa0hhYIs6tntVGvsDajhEpDiMRK1CRkAluKovIZmNoT7S55CDmHrYVSs
oOH3SwUdAiFUk8DWWhM20DuHHlFEmfDa5S1koqC2pLio9sC4uLh7SFj42jdWjL7JYhJ7dbAppCHW
RLj7CWl7kIbUO4JdPDVuIKct0zlMLyUMUk2hjcKCM34dW8Dzq0p5xl3fZitiJlnOb39ib2XbnD02
DFYN6Qa59vA6OEm51M5W4DMz7HkQMaF1KH6a6t7Qq/ZYfgTDyhCe9zclzwHGeLcLQuX0Fo4lSz3u
eJW8hHmbrV/69yVXG2QbiJgez24bUU1NBFzFZq/FByTpGiuO671yGwx1t+LHkRSGBPMnKClvW0MI
ksMDzg9lHIzyRXwviNXLHjT67BotDVceMxHPS9bbBQ+0CJTx27engmwpAbsusTQxEZXQPHMbnKxl
CNts5LwYU84bmhIpSxZ1svdt7vpcmKY8m9fvpr9yc2PlwPMJ7Az2J6VwFJmxpVIC/x+xX8JQ9Rw4
JbPZb9aiDPwIE5DKTVM7zCXrTseNNCk8PWrnDJ2mz5ZNLQYnt6bGDMa2OcjDx8ZeGa26IdxWiTXW
QQNrvqF8q7rWwsO22Su5MuvbVZblnah5UK28vO9UEflBpk27NAUMNQWVbl9aq/yRTdWmjdhb+2O3
MGTxRu+wrza/KXTtrnNDn4sdVHc+RRYOtJSNwExDy5SV/l7Pbtr8MnqPZdmqGyRXUpDe6Fazh0yp
VqG/kwZaLNmaLFDUzq23rM8CFAa+DvqBe7TCzk3ZLBSYC/MJEPKP3AtcAj5zJFrCN4QSR5dSWqMp
VSbiLXq+SjQZ11S3WvJc+e9Fo0MY3QMA/feBR2n8OnTv+PSTDU2CGC2W1l+QdQ80kOx8sNqnSPq3
Nnf7USZSINO77BbQKWj4ncohQGHQIZHcHMwe9uRfT/JGyuv3zY0p5mQ1QUDfUzJ1p0DdnTDPvIgd
XNGFYKtwq1phhLvAqN/qt4oB2oeQmOveDBgmWszAHPR7WnK6k8d0rdBy0WizjJU1k4FF7E+UJQ8V
Bfyfm31h2R2uvLprtTY7hDCxOClKQAuhaAHImQ/lSebrZSP04CTmg238wqEIyiEZwx23JB0GONeq
8f/U5lgBRh1QUAjAZ1zCH8bXwMuevpieAGbqxE2nWc/bfgjsV340QLqXfcveAuJWJK43Wp+GbWAi
JJzEC/uuAZBdPs+avJ1k542IO5hyotZGJKfsPnr0xTA3aPl1/wYENiqQITulZ3gshhHiA/OfBWlA
kqFXtoWTTrqFAW9iNhVauals0Yrcjj/hDXGvcp3Ax2R7OB99RAZd4aGXvhK2TVrtbEg5eR+Jzz6K
Sz8miqs/KyDs+HlxNhgCoNUyvPhTkrNVGR2eL2CP1lxKEnU3Y3suD3nVg6O453VqI1a1eJoSzdMv
HiuKyOipPZ3RL1PvVc3TwQGBY+FbBGsRJAFOcy3w+Y5z+nMWOOpeERj3d50/XndzJARJD1jTSsaF
qDxpfKLDr1gcxjEFY/21W97HzVEqjQ==
`protect end_protected

