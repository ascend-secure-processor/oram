    parameter   LeafWidth = 32,         // in bits       
                PLBCapacity = 1024     // in bits