
	parameter					IVEntropyWidth =	64, // TODO rename either EnableIV or IVEntropyWidth
	           					AESWidth =			128;