

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kHwt7saYGlXQCYfx7zNBKQMcu0muyMYj7eYlnIZ9GFbMNFaUqoFVkIrE0/fh3/gbM4/erXE8aBW6
jzaqCqMmvA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n2YWwWK9C49w9QMtHshqJcoxnJaTNTSDk57vp69IKBB2GWZ4gVNLaOn81anVa61EciEKCD2ETXSD
GzN0gKoSRuSxLzOI0eZv89Q7NIDvDDaOkxWv4kPUID8wzNSzB9s3M+FHQEyvfgEYFnyhpTtitsZh
lpoRj0I2WbAsS2rNjoM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ytM7iD5kqXlqI/qvjYzN7uHRb9YBSzmp7l6skWH2C+QqE74mOAk6mH3I2ow8pv0uEW6RkQTmNWbf
z1zCKCwITn6aEt3IkRhXyW8e9R0ZVctF/n/kdk2DA2960gvVLwGLXpFQw7FJxC/THlhKj20J7nt7
ODTURZ/DfJqWVfJxvAJ9QeNXanMNqzJeRBzz/paI1N1dgmND98IX/TndpnhS//anxgsjk6tTr9f+
MQgyN4sfSUfx0qBaiKl8QUDE6bzb8/xrADB/m57eTxWIqraF1qk1f7SQGd9wrQQlZe0SZrpt/1O+
UMqnts2f5z9BirPqEVvG1tYeoleJ1353IxUxDg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zo1YvHa8zYjMINYzyzAWEmTbEVoPtdgaUCG2W8Tz8TpXLZlX8ohsA33aH3MPP3Ark+vsCoqP4t4k
ZiLHaa2falDym2bkB6X/TP7l3Ya6+U1fSRCBhJPASmoTOQe76ixGVzSiaCLAK+9/w/6t0/HlWdR4
tDVia2recFcVoPWMeb0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tH54zWiDPBSj3ILe+EfBHvu5HiG55r2ommN9wiuYSzRYk70tRtPT9cfgBQPrYMUEGO0MLCPYkOBR
47ck+MI0CvHn0Gqu6rFV6Pl/B1llp2v/BDD+zeUxNpcn5O1PHT+rOnkMuMk4a4/7MZ1F8lRCA4w9
fSuHabgZKyhjRpTP2qwAu7+6uH0XlwSH+hEssr26BvihMXdCfiYgh/XW6KQwuBx3MAGJreeLFYfk
4rZJG3i12m9plvrXrrAv7/UuZVdBNvWigwwDz7YP47iiBAHfWhyw6sFSNQ9JUk5SFzv6BQFvIEFt
zjHEfeJ/Km2jKCGwe37SxYGh3IDpJ5WW5Huuug==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
1O7k6p8Ve8WIqNFTgpqE1uy0r4g2nSAPEKaPWZzkAjiLKfUHKp52Mm0lzPEpJzKTFn56L7OryAds
gcN3HT54u/SPJCjS0+gIjUfBR9rMPO58zT1mrgmS5z2+376bTJlvjtR0nnyJba8bVqN75IljoF5J
h+qjg1GkZmjYHuEDq5v+I+zGN9xb9N24xSxoep7laguw7qCULzB8EQCUvDvNTOnOROUO4U7Hsan/
YffjOTjVbYkf3hO5HJjcqFT4nhdyHZxdVSs2oT5/3oA7P5CcBDmosMPGi4A8usmD2ZJtaaLlsyTc
RrrTTXr1uuCCIDKphQD9aPHlY/Ui9BBifCtoYAHGqxjnlkHMh84uhGLoDL6E4k7XbrnvJVudwsij
Dqb8g0mHuIhViGSclJnIPfQvw5T/2iXJD3lzuozP9zRxBWHpnmA9isrrrc2HiFwvFY7jfNYBBQ+J
3kOJjuzAtHl2gArw1s+qDPmeNqSLMdhPwwAP0PKSzFvJVEgPkK+3g+oxgwlDs7joql4/JyRkaU19
nZrYQUYRxG/XvkWclJcukxtqAzkzK+mBeZQZq3ueijcAAaz4ism/6XUxVP/iQf2XQmVFTQiD2+54
nvFnwltxyGuxgVAk84g/KKSHxxCNS9oxECRjNJFP9GHFayCbCPMuQTM/WpOT0+fDgPKzqyeRPNxb
ZHudLWiVWDFQnkWdFljAnQydtjfFudXnOE9XMo2oltzNu17AUMfvixjXe0339XU9i63fFgG9psox
1IyQ99rj5P3o7xw0MMPjfYKfZKe18YSDHXid8C7L9ExHQnf88uW+oYo+irFji93xMhGN2C9XP8XV
AA914popwkhPmsiSFnDIuAx92Qx3f1dI02w+DgMpvfRPLxOk9Z3zt2ZAbixI5x+0IKU8grV6gssk
gg54hmIb25Wj3HRVPjsY81D4LDT0rR0SlH1vhxVNleGHW4aqNKtS5YNkrIzH6ZEGHXe1ZHW4vXM/
4H/axqPNJ+E/DQwCOFrKblqgLQf/s686Jm9dqXJZV3apC8tRZ4G/LFtxd/3FaOuVsyULIVvW+XDq
czhD9tq0P2qEU53SbvLOP38nHxLr4TB760J5KSYjTcg0CMlYPoRTxLhtSYUYPyu+BxBwjCH82wYq
/BI+v577OuC94h7Ceh7D8Kl+uY6zJxV/V1qKSrWvd01Kh6zHMHPplCK3jqJt/eLfuK0ZaRUOGMf1
/T3TDzqjrmVhokKgB/LsAJIlMVWHanobt9TXT4BhhDKHSakR2cNnqKLE15VxgoSiEDcSQZ53DCVB
tvZioIcrsI/cDgTXqwBAGi2/BjRBx6jmRJjjEybbYVbXhjssq7ZIALRRZ3feeOQ7ZSgWwbt6prvp
87RQnnSygFsrAGj/52fr/4Vcn+s0kuDO4nzbPAioDvQXZKjW+F3hpIm8Pf/rZO9faVfnHQS11MsD
eCLVWO3ZvvS+0XC9sXD4oqQqgpF5ULltfBEGRUgk0eBqUY7W2mrQ6ZHgslSqF3pC8IrPXWxJqK3d
/IJdM49nPRrAfY0GuXZiAMLXISrfgb/boTcxdxHNuGb3Okst1a+kw/DFVVmMJcDZyep5IItcEWhI
vh1mL5gDkkvs37SShzY8uTzyDXzkYKGfmT+/gh3zlU//ZPBSpFWa8JIXnNaIp90DIWBcHjnRqosn
1ASBKXtdG4BPzfGIw+gNX7LDQGquu0yFi2SJv/jN3rAPJffKfypjXMXrFXKgD738odA5imRvXapK
XCwAlBk+PgR3faCMcq0lwlrSNh02dD0gF70LkDYw5jB2FDvcvHrrr7n5D3lwuEVo7nO7KcE4MDp+
17y0BCB8kJilx0bUyQ5bawJcDUbkw6msgR/6/s84uM2BWs+tlhZ9HyE/YYOFNd9SIsVoabmQXNN7
VPnon8mimiP/rP3xOuBmEGUi13uARlYTojjvO0gVxsphmK+t+UmAjTtr6B3H4MJ51Alsqp1k4p1f
iUoYs9qHhfpqRJTiSxBrhRjntu4dvlMa64GFtRMxOoQsJxqfvsYC/bkfH1NozmHdiX+ydt+aaN1k
lJXoNNPdqtF7AtTGyoZRqq2Jsqn7N06zCfFV0eWRTk6qUPq48L4UZqzKoYwlydXMN6795xGoCqWk
tkj3LZC5sJXoBddPBtE4xOhkrGiip06T5bmfsluBRAcgB651ZBoT5HIE3GS3qot8nA3az3fkdTk2
+G2viyHXC4TxtyVn3n/KUp8YDr14X52QUBP8A9l3nMNJUSvyxnXvOfV3bTdrXQvrT1+JsF8u1KYS
Qn994Q2MHIFG9V5sWXoBMiC/32RFyuZaA3lA2eOA0n+c0Us2TF8VmXTndequuR5DWX84Z6ldTf54
aFhqWGJF820m56X05PMXRC4SG2Ob1ie6e+sT1jFmGYqMigj1ZrDSkebP9PLoRk+dCYoahFOX01ut
Z6D1dkCowZyc5y/iYAz4APlDEwOFkBI3NGjtQiTaHKZungp4ES21SC6JJo1FS52dzhcBa41yYk9C
b8mVE59AUen5jyWUcvrAGxA6pMK2Sx7Zpd8mreIN9TTUtwUZ1h+OEMA9L+5Ywxfk1/6aq9Ttxubd
yXGuIvMzU5iN7jIkRo5DM6d0LCGatfkhizkUmRvkHC4gFLfdcl1WU3XKZNVibfmewyNlJUL8tqtZ
kFpZ6TO3WFIr1NGSrHl7LeUBc7jaqXoVOao/KnOpLpYjeT+3I0q0cY1lqdr8JgvGLmDDCsJRrL2U
/AW/ZzKgeKcfIMNjKuH9k8JbL17hlmfEmy6ZXeIW0aKQUOH9VJBzh1GCLrhS0+bj0tDapHjkEiZD
bsfFG4ygGp8VZwAtqN/Xz334/s3xljc1wAV+DabL6LQAShzM+4jXJanFGR7OrE1j+tsLtyqrY9/U
SlZdD/OGdMXZKfaLP7XpABenjRXMCsNE97sBCb5gTEF3wFokiXcEASJ1XCaqUjetgoqRmu0cJhDE
DgHJlEyy6TaX3dx/+yVaOcxE5ToGWfqmOXC80kseKUj4QL53TFhWP7Br4du0X3eWYe5KTV3L63HP
cXLzIWb2u2wGB2F/AbjlYTquzj1oGOjnlZvgnohvnDd23BJTDU0yZc3H1wOUpyKd+AVsJn3jYBDs
hKHzhb1cBU1rkCLY7Pjq4Vpj2lhO6INPmmKjtlVw6fxCC2gkscgF6BSkKOIwNW8fnhyaoCSEFx2v
lwUJniOOTBeoAXiB6qDGBV2i/uk4qowKXnDlfPMA7l9OC5XRTotMv24EJR8kSOeo5Yy0H4Uh1GAJ
16Ck5mkTBHgsfyiMYwmcqwM4HyUVgjTCN/0upFj3oq+MnAl33hJ6AvjxfQYTE89LGqp69cNn6AOb
15GEfTEm9vWxUV/oyF5u1myO4Za0bCfQ/Wj313Fa8P/FsjWuZ0zrfqWyzSDcJ8aGugHImHfl47eE
iLfIjWSq7PXs8dwsdf5WQe+BFgGh8zleQeh9XqtLIGJSoQSLJhM4DFYig3DbxU0wJgXYK1nxHPvc
Zk1i0Hxg+7zN9w+2aQR+qu9LbI+fv7rxvOPfpm45WIshfniaDHprtm+xbMjWMl0+mly81NeVtmGF
jswd22ZYnhx/3CBN16EcqEow9MyoBpbQYK0cl6QpA6U+/PNdNXgfsZTx8knH3jcDwj9Srh0HLQlg
/nFKVIhRmQr6Z7ns6120RaQxGRt96cN8QxgUMmbN8aJ08YiuH/KiVhb7mV6kTDR0TQAWjqXmaAIW
12jj+flUKFzJTDXjmPztkdGo1XpmL66kENM7dXHtbMVh1f8fV9BUY44Lqr8cgIx/v1l/dt3ixQJh
JwF8s8pOKJIQ5QvyB9eaP+dhuwwMv22BTHXACIq14/uznhx5u0Z3qRILpyxerSCFeVdLy/r4YiXY
mEGcJEs2MuoONaitpLMFqn1dVWkZrP7LyqU+a+4E8V5AUDMr1Dq4VZ8e+1TUTpQFxEluBvMXW7WL
hN7aYlnuUBkdnedIYkalhpkJOB0EpJb6wvHJs5DV/KlYGZJnowaMiyd5FBL2jzIgPK23d1FnSyL+
tl0iqjR4CiGBkEiO+xwFMMtEYV0bIFrEp9SuDR0EEG37nMudyye+T8Va7n+ACMQoWKcJReBmEFWm
57iB3bWiD/51QQ3llitu/z0W6CGE5MYgUiWA3sMBBglh9g9+1qGtqP3NDuKhWJHBLlVGdHcM4/k9
GPX02suc0BllF6ihOv7uX8ECJ3/eomikNupnTFhSq3SgWO7/6bgzfmFCBpAQnnKMOT6XUfrPl1h7
w+zIlrd7bYJYvtoUz9F2Oq+nJDO24Q58IDMIcvDYImeu+usY3QiA9aGNShSsZAsJwksMiRa+sUOn
PXpGs4n1nKvyGaNbmQqDSWQYIpdRTeswwWo5EPOZsV4C3YvBXCWF7V8qTdp9I9mphTflD9ZY7XSc
NIoAVU5zjwmFshJtAb4xqJ3dHqEza5CrF36oiP/dX0KAbz/wloTnL23CPG8phhxf1c+CSEgxq9l0
WZ4gZCHLmmqdVxBjK4yMWq3lBsBZ3S4kRXEXkQccj7lq8co66HCOtTqPyIXAnQhCcOEyoVPokglq
RIjPypG8fGHLxk4OlR0Zseg8z5d2OhNZ4bFrJHH2Y6Oi1PI+Cp5npJ4ZCe22D0F7Z711X7MS4GJL
PxXhPyjDsvNOStz9h5Qg1dp3oU/j5vymVNzOH5ftsYLqOMMrYCsXcEH/TZ2K1+iJIzA0BvPvE49G
vDi3qeKLjwR4MPJMGeDtxJ7Xn0U18nC2+yWr6DNLqWpxp1UntWmoMBAGpa42rdoy03nIQW/sZFXY
1p3VVERtYV0vAHT0ysVWGs/fer+UAsmEXcveoic9jQqP4FFkqibmRVVmvRFLAfoLShVRP+30T00J
hVZBUFyhLHAk94zdOpvRcUZsHX1HshLjW0+EHqd6BZ85bpBlLbexlGu896DOxjrrr7G9AKo7N1Nt
/OHZGgfBZNP8rF1Ot2rCvlkuCE8AwiDEl81W53LH6gKqni/JjYC3L3ynT5BYFXHRHlsoX+eYm9/y
GfZeW8zgaKQAM8gqBnICI6hW5bvl9DrPoHgWuH66t1tPkaGCxbjyoRJeGYXxj1rOCv/EBqGJf8Tt
UtfGpVL7XXv7w2BRLHoo1F28pqM5hc5Yj8NDczQ59PvVVLxlEd38SmjNhihIBaPAMokwOq3ECz3B
OxFhOUqL1R40gAk5AcvkFCVRX0sENxaWxZhYmFTuDIn6nU1CrxcvfugHH0TRsesaQmGzFAtDDZgW
u3i7ovtGz1H33cg9oAwMC2zbAOp6/32QKp8vbZ+ybSPyQVkNMVm28LPSEcyTR06tZHXhbujn5D98
Ho8uDFyPX/HGlr6FHmRcOMgjx4zXPf2YmZ/po00M7Syex7PAv2j1GHspBMR8aizR/yb3rO7wQRYd
/AV7bmxhgkjYOxUSA+twWMp20C2F6nebNPkHQhj27eeoJzIt4Pxd3zYNjECM6A+PgM/JIZ5ZAWbZ
IIZhfd9ybNp5aZeV2qfMRnj9H0+g0Y3bbHOsCUjNbu3ylJn1QPpuBxOr0x5yUN81kR7ewbgXgEj6
OgOhO1M18TDE8UFA65WjSUBiGQUbuUfm6SOquN5m2zgGO7xQJGsCn+lI9ZglLrgLiARytOXXM6lT
wEGWibvikCP3BvZzKByBTaYBFWpxA0Ge5fnmCGxNLQ35Tcvq94X0JeVwknCFmrTRs6MZFvfkAGJZ
tQhqEs82DaOoO9njmaI1V288Ulx+8UFIUjKd0AAfWaXaPUKGjmpMs2Q6EdFgyCrl8HmS6IdLURhF
8afTBFYHngWp3ETNLjoz9+/9SzvSDgqodbwvxeWG7otVj9c1Iw0I5ccpJonPPlln+uo+upLZDtLQ
p+B/60zJtQrD5w+SKwgbd7vSPP3fu5oXrg24t7vyZohLEAjqR9r6UTMqzOgZBc50EZZOWHu+dZH+
lPKOqd0w6p0dLigyg/5CFBHEvqPTDSNNE3fMPpjUBS4BmvMM129d8DbXkIZ5XbbrTo6gOPxAaCkv
sjPWJhRV7r9SiNoLEqdZ9TSUVtIIBA2Cn4x+JbO+FhVGNZtSUGIV/cCnKYR5fGeKitoLIJQrUkcQ
m554OuNowgQujA8lPgNsPmt6knyShj2MO0g3saL654mQ20frLXr245cZoNq/U7h+aN2p/z9ET4Ku
r4LR9R8EqwTQT//1/2TLmFo/X8pMbsZJHlzLIZmO5+qTsqWK/fFiDof/ot404/52jlwhi5J3ggZr
wkoLheqnkglUP2+NGdeZTZcK2Mw1V7RswM9b/KNY/rRzpk5gJZ93fkQyTkwyxD6MdvRUOtNxELdK
RIzmiNtw8deU7fGB/RaHrBSAy+BkAFKSKUZZVkS9mciExxOAp6U6SiAd/1fcK8uLfNwxIE1Rf8aU
PD32lOnFIm1XWyKi1gyCgF5uMmFDGOmzzkaLmvj5XTxMSGIyhlDVFLL22qhY0Gv8Hy8toyRjvbtM
HfvuQCe/D0YjRYuB6ZP6L/KBnljBH9hQuW7gW0BFkHEoEBZLgCEXdi5fSSUvsGOgdWS7tFB/jTHs
6N/IpxNDb6EZJ++iTRo+fRV5p+VpgJ9IbxQJKns5jBc21UQAI/i70+8yOW7lYvSHSm+f4MQM8Pg3
6ZLb3sI1pIuhgmYjJGmxSSqCEg/m3iadmRk46GhNG44x5Eg/p9BmRDFuxNDnHdUBNabrhl8tq699
iF4E1Q/2ZBLiIq9/7ZxhUGvo9dfhHnfSU+N4yy2gboYh5kp+0SOMuoe0nEUxfIzHnpfovBp6LVb6
+VzuIdZdIETwVDmmqJwFZ74rqRIPM+ycEyv0W4AYG7/JwsJTsuhYl9rMgROblbLbsIM8PfgNh5Fv
Q7w88AKOzsJaNvQ5zY5WzzvRXfnQ+tx3FrQy56raxAFvzPEM3IBznskD+thrSBehB6C6/pqTyp68
HrSzSz7UixjEbTSya3CMuCcE/sX5M0cwPmMyUHFng3l9M5EGGamg3PdvYLvhgDa8ngbasLYQIo2d
qcfHLQ==
`protect end_protected

