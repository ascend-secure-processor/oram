
	//--------------------------------------------------------------------------
	//	Data Mask Width
	//--------------------------------------------------------------------------

	localparam				DMWidth =				`divceil(ORAMB,8);