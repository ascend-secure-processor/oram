

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
I4rva/cuf4t8VxEsBqPu8efL40TgUMkDqF/Yo+sT1X03Oj4YCLT73IcHuEBecAB0Yk1189v5a5st
XG+Mr7PHKw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H7bdBneOz64Hq0fEibwIAzUnDzdzMnokctesc4WQ6LqHdwGx7+Tvd72mptonuIo+tHt4VMorxvNX
E4sey2qbkiCMVPvUwzQcgYpz6zg67jAFITs5zy+Cj9JczQE/k9WvDA6HHh7Ck1/zQ0P3ltwJzZGC
DTv4t0DJDMfi5J2olWo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oRLeBRLdTUZp1yLrMwbsUOF/pXeFH1d27D0aDIxZSDV6YvguOLzaLYZyTZrxvG5IB7SwrpBiiiTe
QMHB3zj+Rq1PIUKWdQN3J+YEGXLNXyYh6cF3FzhdUnJsxJPBYusxmlKtVZccmmDDAdVMM+8eBrnC
2fdqD7D4gRftGKSB7OO4hbfZEEA2blepsYpXd2aON9iW6qegOSqF45zSC5iirlAhcQWlUBYE5yAN
3B5dRRa8BpqruHnC4fBMMgU74YmXJOGVqtf/TRdxUuUh6tQbzVYfN5bDRDi6TdYYHZmoGqQAesjP
clNzvpNa49SD8benFeh8YVwu3vnFCRGfa71hbA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bvaNTGZ21ZG8Nb/2A1Zs+NmKg+RCqqnq6+lNXAHWKLXwRic7v6RA+LaB037GVhqVGQWO2/AtGEKc
bIKDBtZPKPVzkZHCa/Khzs9+YhYProEjTjFLQzW92mJh/J2A3oo5ZAvIyXPE/aYKD187Ap3XrgE3
TxiErtJCqjbn1Riy0BE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EVVLKsNrt41GWcAAD3vdBOANd28+fR00pHRU3ceOV66//xapj9fdQmeBSf24gMdvVFv9nQyZ7Sex
eh8VUE4O+mCkHAcEnL493jLg/U2qeo/QJxp/jsbtNMcj2xcHNqd6Pnhp4f2Lbb0Q55x1Hyyc7Up6
F5ejmN1lAdlq+/Xnmjq65LEoiWWRn0W5RL+AGCq6x3o1ELaGrJC8x1+D/MqhFJ4EaJ/3APdqabvX
XYWRQsWTYll0dGph2+N/C51EbqUd9m78XKevLIgue4dYBtxIgDefDDcktHqg5qg8QiXQeCzxdXCr
Mm7bJZpL15/3jRwlA36jZGBpMcyH7qbm6m66Lg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 88208)
`protect data_block
jFoGpHjn8W9aQnjrYvpzhbakYfQCBm0BPZflpWT4fYn8abWBeDfUXrXQ6XFCUEznIDgbt1lgfTCB
AhlrPh3xaztYxk9rtOnagFpNF2IDQ9VXA4ZZrJkTnAWCba6+ncB3V5v99u2velWehQvRE/J+MKwB
1aXny+EwsIXlL9S4HfM2V/d3zAaseiS01MD4Wa2Wn9i+3GodNk/KUgxImofqSsAv1JForjgNWCMD
O5vG9v1Jcyi5mD4SkEx8yNBSUZJW7ePkcF1Dq/6eVepILo/FfYkjPGf5DCrbuRPq/9h7FfXnHscj
KHkB4/ZXz++R7hCwc2wqDufmq4o5meCZSlnC6w0RZ6a7hsdDOl2hCCZ4qPTvojZDFlxjFLHsP0vZ
NsIxrj/kmlkuTiAbpqBAX+n49xpzTdHKWROVWhdXV40BrdZs1+82WQXY2RggW9VCMoqYBFmjfBV7
IIbAGcA0PVZc9lu+bt5I+M6jUzdKFeHrqij9BLbgsUmvlhYMjeSZG6SmcXEtDexeuJYyUIZZ3+Ns
FKcFBizWWBfnyZeolHl7NDoXRuzU63CsRA9V+eaTh2IfMV8xsIWO2FP8RNYURlVDGYyDHSRsJVHq
P+2DN5UQDFk3TdDDQr1HFYnTKIH14GoR29VJwyH1xYgTbryRIqo2sdszXLt8ina0GgDGHJJkWuhi
8uCi1fx2XgAPAChJ5Y8QEqn+lOTbpZ2kvZ58iei772Qq0Tx3/d5EHMaVQ0nzSnV9vEQYleT2shjM
Cgm19pnpSaUZlZHt201Gvwt6ymlB7Dy6Q7EBsz+F70LZKvR1gQmpppMpIjzXyT1nVAfm8RdaxPkS
O7aIPnbjry/8ufqQk4niyF5MRUDGbRwYBoqq7ojXnJVciQ0sbmCwmFK4ixsSQDR7igd2NuDc5Sr1
88pUaMvADYfR+N6kYUiaIgFy97smOd1vPExhCVEPc+JllZrI3xEDWxrAwTIUFMhWJQJiBNpYIHMO
FlrSpTL2PoZ4xtQnWdS9GbXQSh1mqrHUN3iVRAUUpf8JIcptCbf4Iyxcly0onVdzWISv2vGDUbpG
QTO3x1Eq1pfHrBpvkxxz6QRPJ34/3xX+PtljpPsRiNaqGsUhgEyw/JYauEUXENGhbdsYeC2ixQP+
7rQngbf/793OdiXsth4L11FHm4YTQI7R/et2yiL70bD4ssXYtAuzIM60/9AIdxlA8uF5QdktrmfJ
dF92x53NEeUlvrpj9UVRivWVK6oa7VReZ3WA+jlzWYwukdYY4FvWqsc3beXVc3WcIa9DdPYafXvB
tnakN3j85h0FKNljfqxczF6BLtdkq7G6OrffrKeT03ekp6s8mZx7soUX1o/Z7burf7UsLphbHgNL
bFBjbCdoDfvi3v+FPHvak3Vd7GwEMAhkbTSIdBtjfKZv8dFK8hpVM03YpzPZ8vOzPrkSj5DD6h6T
RSt+2vIrqNWY4A7MCWK7NfOVmChVtGKZR1j+NqNwozqnuzqI2Ohl9WyShMpMax4sUZ8K0iwgTAKz
Gi3QTG7k2zHfwfQ9k9aOHUlQlyQAAyi5WdbqV9v599W4FuAfiHpTnkCtbySUQ9hioqelmIJGl6a+
Po2f2ynEc09lSzS0nC49FP9z+2A4v00YmfzTuJLLVsEOej5KZMvR+VgI2zlP7F92DYvetVK9/1H8
abpLWzavjE+N7iGJkBKFqDgTiwm+00jCc8RMtzFdvZ8R2Y856s7kBAs4ZFo3A8kaiWzVTkDk5lHP
hhusbQgV8DTtRR3FDOux2i5/mNKg9AoqQ3GOSYTT8tDN1qJHk38AXIub0BaKHUWixy5I19YGKdmV
55ceKvm82x+HMilHO/VZhxFU8GPsWqKkOufWl4q/cZnDYL2cpFwome+JUQroeyhpsibotAeEzRZY
NDZqr5g3yrxGwZ0ltJtPULQj2mDuDxO13TMS5OqV0ewk0T7H2jWLRkJ9DjLXn2cCOVPRqVzeAgK2
cg9OLuC2IYdr+TsabXPVO+y2HexO5emDINk429qvXsf4Vis1ibhhbgh4ynOaS7BvZLePaZN8CSW3
x9xw+5epGWQUdQEMEmstcuovsEOtT5vrN75KiTxHSSiexlV+zfDRwiUJXKk89kFKCypiqhFwHFUo
NuvGT6kL2xA0PVImDoTNpFqsbW/7SBrlzCY8v0fAgDBFPy5MSJ98K2Ph9+jO6PiShuKR1dLasiGv
ymjuhHSL3Ab0gdGtoDZq6rP/BCJwLSmX9NXsUCWsKQFLSR7emJ0FvdxDFNSYLqUJyCFEBYEFiIX7
2ihcDL0/4kEFcTdgiYvI+zRljummSAkj9+pLmWCUfytZCExnio6PdEuFhHCsTR/ieobhvcugb29E
Bl+r78A5d5NxMFzmHcBBfYulm+fQAue0F5JhZC1eFqcGsKdI8tDreCwSNAqpc0LAqe2N0TDW/K1L
QmiZW61d+YZ0sCBW7Z6bwwnnr/6uGLbRrR9oq4b8JzFYLEkQFfkRZfgCUeek5tevsw9OvMeW7VB5
NHfILwhkUXmCfh1rvyfduALr4G/Di7Lq3/Pm19UZ8C5o2Trcjozl2uzEOm+WGYntYQhWZoKPAfty
DA+rio3+cAwEFLw592LAm2zvfHABnLYGCag8jx5y0y+wv4BYu9GvoiZbX9ecvXCD1js+lQnwN3x9
P1GACyxhUouFGU1FwfJxi8iDII//Hfy3WFu51k8nK2i7KDYQ/zaeubXFF5rjC0lQIIrFNbTaTij4
QkfE4HJHqPPjkQKFeOUWR8dsW9vT1OTgnanXkry+zkqfMSkOhgsEyG7sxTx78Oc2J1Q2AIgf0kkz
Y+mBx3AjzpR3kDPVDiahKkn9dSMsb8cEyQIxg2InvLNg6DMivaU2o1jUFwSWyGvU7uxBBwLcK9OT
pQMdEQKv30kwYtICdFM4mbHz9tx9FuQEpvwQoo1Ak0gCqMrcUuhe9tNQYd2f8cEFlf543PlpTNX/
b5EmVAHlZT7hW4qFYL3hNBXSutTbiqGbDJtOlZOpgoV1VTjyHtGHJsnohN6J4/0zNIzNrDA907fO
8EfHSl8G0RxiQqG20r2gMQ3vBeSmQjXDHRlHJrTSApZ2KxI9NRNWYrs2KFlrshuTPowaurvklBfw
wvBrQy8rq5h0n9gWQ6ha2CwQpLmFbABI9bTltUEPIYyP27e1OXN9szrk8qJrOv9cJzci/m0fyJCt
UWovsMHOh3t2g2wd7VVv0HEUUv8+cy7Udj/e9qCl5BPn81cZVL1R7TnkRa1TpHpL2qblrTQZ4af5
uOwpeOLbPHY5NtvMrTvR+mFXor42+0J34DipbZehS/+/4toTWv751Oq1gy6Q1a3E9yiJ2lb1RWpP
mMF3GXKY7MLvVGRzdasdUnZU7EmCN1m4G6SsCLcZtqUpr7XYidj9lThN1JFtM9x7Kpabcga3TWLT
JTGtQVd3SZ1dYrE2IOqtHbchLD/vteI5Eceffj71ien5SxJkbcRUSX9eMYJJ20pEt1RbNg3LhGoK
8XnLExo0e8/2VqzmpoK/H0YB4Ip57Djr+uFTqAkCZ7ZpyT4YlYD7aszKi//mZRbRhugAEnLX2VZy
LUnSo/HFug16pLDX1P4tP3HhnRxZ0aRCttj7wkXBe919EaC0IhNrD2KnV5HA/1vuSQndGuDYImPo
ZJzLhAoioONjOWu6+D/PFV6eKUG4mUmSxuUM/nw/pSZmmlo2KsWmUWaimd3Hv0V9sd3AWoqzpwnI
fu1fc220k153DJZKBRSRUlqO671FQCp/s4tibW2kyAZDwc/AXu+WfDHRW3A9fcNCx4oN7HT6ZLjD
C9xLHoAlDOjHLb0DbJ2LsJk0LYvDQZQIxydoSO2mB8mfl23xFmF6a7rIR3qZ0+YLrxWZvdTKV34a
k4uvPNFpUjw2xfMrxVmgBjhsitQf56+E0U0frYIB9kJgeWJeUvNMfDpt5/+GDxdFDFeoxiqlYh5P
3uc6l3nSBsXrHOWZoLbVuR3Pa8n2HnUhWqWvAWFPXS/cu0y5uoZ1mkZAgF+b7c8Zik3ViVG8Co3E
AA/dZrGV4KA1JrFPpOmumUTs7lomxYyoRPZEOzJmyNNFnQevaqGqkKqKTVE9NuBRQOokdZeJzjBD
zbaPXDYJyhWdKC0aM6CSl3OJE538cBiX2Lqi0BSPrnB+ITKRcztH1Ev8CBZTm6LE5aQwsb+4W2gK
2aswwGbdew16FyaxYfZjNdzYhH4rKo6T2tfKwTGr1mxC1NKYn3h2Fx09i32Gz4Tx8Q8yMh/2nR1G
edqIB6/vRLzQbWSX3u63bffmjQh0/H4Gewc30rde0WZfmPBRMp9UbteWEyynlAVgtki+5P2ZXawd
LqL0nG2EMSVhspgMzgtORjEg64u/+ruWYIQ117osNdXBTGmKVJOUkf0pj3rdH3riwizLWtgrNe6Q
S7wePEReLu1B44qB06RQnzgAu6xfW6kDrUgRKZpb9tXwHdraRiF1vF2y/7Vvxi4nVyOKAkyjnHaI
lxrpmrnRPWT71fFF/KRdPlOxTaOkofPSHAAWqPlxCAuwAwv0OpIYrdSCNLN+Gb4sZ/6ZA+4k4AQd
ObAMhprwb0LfGoRZ9MEmSkG3cjKILJW9sdERVfs5NePOfbOVldZ3ZzQ9uBiISnILA/j+qETbXAOy
YSmmE6wFDlGYBmDY+I3+apOQ9KrsHgf98gcdWQtrxyr2l6Ab50apvrxtMPoAFBccrF6MWRRwU/Mo
OYQuTi+4OESSHTKyx8uOIhsXYx6QCrmqy2djvnVQRs3j+DcfNIwfwjdRtFJzCONp+yiNz3rNVkGT
RurkkKbo5FF2a4ZGbEM5Fxjd3Tc3bXVMwewFNyDyvMMFAi1KlxFVlPFtzPJOSvwt8GBoj2qieC5X
D9lnjdu8wgPUQaafwmoFN4r6bs9UtDOt+N5PVVPHdNzqyCTiiBV21TGVBe5h+RmEvlpZUDOi7ea4
CQocFQrIgKmCOSSXQREfjgAMZVRzit7Ch4EVgoXCgb2TLzzJxs3u/oIVNywz3i5hdL48wp93U0FK
NXvhwfSfrQp7cXJE60lqu0RDF3FtX8EuXty6M4UpAGDnp3dHCHrNkinLzN1YSoBVN33VVy7nfJbe
vFXv0iEe1vXKLckjzZLhQj9Mn5DjqUtPK1Gdm8jISIa5ukpR/wX+uzfrttrxLjo/spLm2uQ1D+y/
fO9WHcE2Oag34hCuRTSJB8Fk4OFK46325wQGFdVADhN74lrIMIHmARmG3rdPW0Hdg8/ClqfBM4R9
UEZihw4pALvPaEDJ6NRN1kqR5nJPkMh1aN0JUGvXRgQLTYq+Bd9kEqkS15UXpWjwk3wx3GEvBNZN
HYhVcDZEmVvlZcxjljCn0xne1zuQLQAy7Ur/oV9PGUCka4BkpUzzmOE9DRvDU1vmmPG/JedizHQH
MEamdnuOquMhxEwFF376peVHU8glYuOUpaT1rutp0FvQRV7dradn8kaTDzwPYxzBhBdZrrsjWz4l
wf/ixI13NgL26O7TFY2GCas3g5hcdzbe63CrpLxfko0v3qiqk9yAvEpM79ucEOgYuD0OxLHg28NL
6TWERNu9yjDbuX3CImugCUX9Z3HYuPD6Wd2y9qG2HQqrUwhP/50eoU4SkQA+qcc1blFC1aieqsTC
jVbI0gFAJ/XJ2IMgEPO/sWgOu9lzphr3SfJg6+LaF12KjfQ3pY1/btb/nmfPsJa+GOw76OYjxzZN
GZFYHKx4EvRyJOpW/qEmdfWRhNCcgxdz4RyQs4pZBCmhkPFlG5B9s/+4WRkaOpFlNPDQ/OyjzSo5
qx47F6SGuDp8RUC+6sae9lF45ohuoy1CQ/sKt4WSWSEC79Xw7SwnWwZIQJWF2NPk2F64eCkThYoE
AG/l83PygHYp1OuFlCBDSBZc532PAgP6NGdm+icoBfkjM3gHgMLaiCQM+TsuTAv5rwTOA4mbfkZA
R1gnABuu4D0I46unEfUZmUPmbTLc7Ag2czpsYkwXFLiwmkqIbaCOFHmHDdUkns+zjj9UwdxWryME
ORGXquL+lIaSngHJbI8ripKMVtdhxntFN2SpQbf//nREk2XqB9KEKybUvoeverR/NH4wXbD2dnqO
Bv0moJnlpqRtHSDW/16Eca66QFWBaQ+9K1zCpzQH90V6zhxAJQALS8EX4PC36DwmQWK9vcKcX74m
jEFjoZndR2CnLCe/a/iMs8XKkc+bogTdZknJVmoXHy2TvBfC8WuezIM17qrdW3GSpKMJNWXXZUOP
4/+2NewTUJlhaz7q/2o0rz2/uzS++QUDemEZaTY2Jlbqzycb+lJ7fkrnSIlYoUThlPtMuRXvrMvC
Hem9Tgi3yeN7lDUFg5J76jSQ9bjsiv6zwkb4UhRRMvySD+w3mbYVQLbVjwNQkxkACo3Y09babMO7
y10n/53rKKwiFBLtIZv6Xd5/bQrVYcT/eAf2Zs5xkUDm44vb2t7cU4lKSR5uB3OOMUytMQwVyDwA
gnwkESwShKZEnxZ4bA4hszuqSX9HoymfebI+ofAG9aEAuRpaOgDr0ET4ZdA/FQIJwNh3jTsiuhdK
AzvEh7OGbRXyNyV8D6gm4o5h8mZ9vD6s6rU+d3+c4qkduqAoh6fm8wr6cmSb+6CG4RzVzFgxL6FX
5TFdP8lgArMriizhmLycSl+VeKQ64vadNmNyM022yzuPo7kvPN5IATQx5ZqYMAcef/lqyEhdzKCY
drMLvPJmznmtJW+3CeVD5AmAk5Ql/+10j2GpSdn3wBfwtvPLouJr7SE6hDHzJUvggKbcaxqVLVhr
j8ogfOd/qJFJS3oxEtUhDCISUegFvb55k/0VOL2rxQ2z9m8ZQq10Ys6wWGZaIyG/7FDT9DMDRkap
AYiJvZNTm5G4iDgoArGnLpBsRB8qc3VA3ISSPFOp9ATnxR8OEBNshYaki0mr3OOFTa7S53we0oPN
/mX9z/lqdEUdMucx9593LyWr/CXs6b8TK6/jDWSFv82LH3nR+/5I4R5DDElQIBA/EDlTOEwhq7Y7
q+8BJ2oa3xGO754/1W1dem4rG4Qyqp33EMSHISoEnrS0KJYvGM3ixTOx+uLjsCGHHEqmgSsJBFrq
LNP5jUckM0WFY28ooh0iTjjTYwcJHSMRAbmXhDMwR2A4OF7QVCC6sPCA7c2TuT8Ad8oTQ7pBB/9a
W271TwgRHoicNuQjqjYHvVerbfr6D4seJwJ0kXfAIKLJALQ8r4M1QgUYKrpYq2wNbnW71ksMMaFo
ZKlMJ+J+QvBw7RH8geMTFIuApat1wOP0CRm1BzSL0pGs7Q5fM5wH51NqZ2k+0zGQqfmQCQvoMxre
5xtIdW83FeDl5VKMIwXyW5wcYQKrE4bWJIPt6H7OogIUXIAyafjnFrtGHdi8lnU4IcoXQqSb2ksM
oZCbMFKs3mpvkHYpAmS838QOnyJh/UmJ9adZcplhaMFfXVSxbts9eqP2mfCqw2sRe5mosEogkxkl
rRXnDgip6dCpRV6yUa19UnE4OAFWgO4qGPtzS/mgEgivaTLsnf+eGrd4QUfH8Q06YwTGIF1GXhI9
0rnM4S/dsMoOEEpxMKN/Zw7q9hhTp+VkPTGrP2GFnbCM5Y8e9Imes/Eze1VTmH6vx5UA4lvRzXmp
gNoGRkgIFAoXcMolA74MfUHYQJxbcGmeNh0QBVxV0aaqb6nwgDoTFiBPd1pPYt1iEmvJUjibB0EX
nA3ZGL9hTDed5AyWDEGT1thSI0ZSpeIHErteDfL/KIT4g0FvQNaX4mlA06vxbI3ph2Hy1OoVUy2e
0wEa/UXygdpXrxEzpjSCjF1wKSNzMTWqw0VB4W21frMr0jafhGqO395A3bFwrYHWjg2hQHA8CWYN
V41uN/xm5g6wbwtp04ENk/tktoLAMc9LYa4odCt7dhTD7FHW1hmhdO90P3U+6EV2e96kKWsWOkJw
t0dWpXNk/MnzTtDHGvIpbNhgLl5X3bOTiQjPlrTgZCzT8jtnaq97miX7y3iQgljD3koAFA8dmfC2
J6rgtvHSwsoodJ4cd+ai+gB6N822hEulhMzpqhPZWD9uGlNqNsN4THxh+R2SJyhexSxUSgDIN7VB
xV04U8rUznJadKIqx/pCo5AEXUVLkyee79V8IXAcOY8UVLuI9LUrL3EauVM1VJO7Wf0TNKs2Pf8D
3Ua8qV3ac2DF4Fqjfvt+fqqPGcSbKE2KFJddJueaCaGMpAWn13OYiAxJfl4iYhrQ619RMX8LN6QY
ciMcU8n3BJjg45rrQ40oe3n1Zf72dwsn3cjm4NZyfi1whMx5qsY154ES/YI7zbiVFaY9zAlTjksd
MSlcXjF+GhL7nRP+YZEozqMdBJKmEjBt5LCW69nHVEcETp+qfSbYUyBbx6cN0zx0NBUa5g99fLQE
e7aDa6k3ojsdLDw2L29DLmiAAGN4zv54a1I4M1+iv0lAgoRaCoXV2qg9/APEv1c5suMguZ2HHaM/
hVUCpFzNX3WDiqnwiBgi1qIe9/wd3A7lGoZ+k20QRmXSCPjY9T5GialyfHtuMUHvPJJXKNBFxR3n
GUfc7ySKdwdpbQsX7yTHSm7hMzydcxl+nG7nVG1+qfsh8m2ejA09cBE5DvcWooKKwWm2GkT2X3/S
8FtERVqTn/wuoEJjT6WsHtGS5EOOpOoL9UQfIEqQFo0sxeEC52mVmmQOVve3rDpigBVFT9MpOreJ
3cbPktF+oybTZ/NT6c4z70fd4mlW+mJc/RMOdaR4bZ2+6WuZbqkuExD8uPBzpLCB2IOZpK6Hg4RJ
lwq+d6lRIEcugznGDwb0V8rFdSgue6HLHYyLPancjfkQ7RLmeibeIbKOrnVKpzk8cxuJ488vLC9J
fgIdKK9MDMGAnc5SkJf0SF53Q9X3Bx0OjBk1WMV01YgP4bedwPJ32cpvIPPGDEcHkyA4nZ5fIQSK
kw2wGy29Ydmu2KE4RP3odwkrf81SeFtl3vg48AIjI9D8kB1IZwcjol7xY+Dbbo1uKsVKI7BZNkzY
eWPGk0pMRArMtqpNPIAYtYIBgq437585UN5lwg+1I5pMw+t+fbWzVpye0gfbauCE7Fyg3Atqzatk
C0P4OZ5INuLsg1wc1CATgTS7yG04/1pl0BWg+L8b/26KLEGr0nNZQyo0XXRmOz8e1WcG9o1u/lxJ
GAbeNwLO9v9rPZeQLV3WsPdexH4Y84CROiw8BOt+qg9xv1/26yycmJvM9T/3TEDnOwz7sm0UNgfo
F8dli5kD8r2ZnF+MLU0lActa7RyMkCJnc2PvBdpy/AUWBh9n1+gCIr6k5hwI8tYZRULK2R30AFrV
AjYdvsVMaEkNjUqZa59ORpDcDqKaipF+kuOa1I+wXLEZid5JSTVQQHYM+RaOcm+aLoViUH8Y0SeZ
ap/isaV2v46SlSy3C9m/3+9iMUz8fHMJUFO7wGv3DKrejOFzFj7cpuXig0QNrA6Vlms/1J+ucsox
MYKJOfFytSL333/bC9YcEL0YnTeYAGUzlPNVnopGCxJoVwi7xJ6kKNg+3at0RCSkNZt3i4HMG0ZH
Bm0Esv5RrNvVYzhb8FH811ZBch2kyPboqARUGzELRoi3DO4qUUXRe+GC3O+V9h9dhou6z3DZ9y8b
/Hv8ziA9OBV5+JF4AXGxOIHY6t3fwxSd1tnQl2WhWCW0dRwquLUuNQw6gpedSufWVuP+8/nMVQ8K
VX4mXlWaZYTiX1bq8lpjM18M3QOSqHNEc1KL9nqzP0Ovqx9vonIm/uKRfQxhXBChXlCBloEsjg8o
xIQn2dOkCcWvt1+QFkSH6kmoFhF8DRiiIEaq0ZhZBSYWdyUUTjr6Jx5WBNKf1GhRrsZdDS10sshA
3VLXsNXcP3VlwDiDk+/18c39clhVmTFCZWStzbZdcMnKDaUIxOpIK0Qf/10AjvkZCd6a5W0sstzG
vYt1Ph2M6Mu0G2XljfUa2MA6shP/rqiLABwHt+j1ITWxO1bZOpnePz2K0izKbAsD0LU8z++muyvT
+Ke8o4CNOFYaWxYQGo0Vuql48nI6k3QMHcZvHiOolSlT46EJGgT6t07dmca4JnMrrM5u5KBl57f+
GQjuXwo10r4m/VuwSQbMLLMd5rWGuEqdn7QA61O4WEywKQtPCxjcjWbT07ab31od3jpIjsLMyZSc
GXMKS/jz2QhxFXdOSD8KL0VXyPmeQZRdHzQvngSCR0YDOs7X5a5iWEDqc5XyW8ANaHEpO/UN59l6
KjzRql/C6Sc6AwKQxsz0nDcBuQln3HHoSzsIG3r7HlK2YnDXrC/kld1tqD23MkaP1TF1mWNB3tKy
sui1qowhsVwurJ7SNxgoLr4T7lnK0IjdWkIaLUdpbc20DQsxGVgp67o07lwPUC52SSHVtnDmzdLc
2GyNfHZrY2AmaAH+tI3l2oJaimQy4TLn8fukWHtHcw1C6PScuLdsZfioVxmj37vYKe305xQ+++it
YMnit7Xe9BeKKZY8Eop7tMBpcrNvgL+qWEGvyiReIbgnzDzE/D8CWzCU8tOGVePMRNmuYp8EOHVm
jdmwGdgEezBwRvFFpduFEL1G2C+u4T+6xPDWsisTpVbrQE/qSYTL4AGE34qlsq3NRb4BeQN8wPme
Z1DMzhM/Mg1ncNEfOEssSI1Lxlu7Ute2QW2VfKy/Qm611jdIVziAEv7/2IEFWbYLn9dokG10AGJO
GiHcELIdNaeygLqZO4JtRovVX63PdgWLfMv5rxOG/m93bZ2+cruxSFPbeSJYNKnrAJxEwztexu7c
O5yXx3U+shJUgDRtKNTxJ5qj7f1BPm/Qwh+r9VoiQ5ybgz85h6zsF/PbZz8EKR699URHMZ5QujOJ
u1swZxs1QtDVf9/tgx15af0YgIehhn1AabWN5V2yPIlLdYTKR4IYa3JgCfTqddjJo/odeu2MIveU
pcPMeivtEg8RSUM1odbAOb/qPdWGajIKWtVJcTboWcELxfudQ9dFHXvPstiGbs9j5cCsh9x3E+56
bd06w/4Gu5Kzvpk6h/LU4j0oVm2Sjo2YaZDNcCkkvaN85tVYouLhvV1XmtBOVCbZkDTzVLRGyOaf
9UxAtJeHi2b3G4zQc8qXxlahl4b2RFiC86SAJoL5OLHOeAugPtVD+Tr4m5hw82iNjBECArUdV7iQ
0gunj2mSqm5eXD3WxoYQAO8H0CB4tN0aUFg4IwrdLmZmQGxmVlpBiac3DkGFMsuiVfAoX7euzOfu
RhFDBATSLIWLaCGV55pIy0cIs2JF1HSNbCHvtwf7Q2og7c4CLyTlm5aLbRSNGX5mtfK1kcQG/Nft
eqkAnj3BYGdeUN0hpdc8LkLDVGKhkvmG2RGFKkPUDJc6AGxMzXt82t9YmXHkgMZxEkf48MmNYyY+
INfinr0CyjN5EY684diRyDXo5PBwdB+hXJSxcWZT3+9xQLpLebCxBpM5zaq7RBrjEOwG2aI8EqSp
rhD9oDFQH9VYtznk4KRY+WVNEhgjAZmVLvQWR1gthFv4mAMF/ZHv13SX3TZAPWGlHyYUsx2O3dXr
s0nGvoGA3H/3qmNkeh/91hV2x5eepxJS+SqmLugZ2r1kz3AIda8yTWi4vvh/ZfUBePHnepgRcEoy
Hoz5sX4PXD+uwTcCKsxibSMh/tUU7OhEk3SRJhCUC19m0XoMWXdMOnXqWLGm8xezdBT7AL6TS9Sp
h6lTg4lzLJ0fOCNQnKgYL17o3TtgO6VSXxturitFbp5MtEPj3UkPD2gBICt5umqiysNJvkHoKWxJ
wIZZC6ZEl+cm/U3vHA5QRDHqSFiaVgm81tNV5yV+QGgv8F1qQtroVpXzywE7DlmiNLZbUVtMK/Np
OlcBVJFW5YaUUyg5w/Yn6szTSNtR0sTGeSwjm2pj8oReNsMV8aRXv3dd2gE2HwagpczRzTZPU6hR
csKxrrwxTaybaHNr+9TXH6N8xgePhs9zBO31bWwgTBunXfPTNPAuDqz1G69HNKKPPmbBUe8yRvFD
tS0zo/dSXFCKXnf8F9LPDpgVMJyJO7NgVYn+sYJZBZuS+0T49cTgQtoy6TjOdXNcVLjLUTzgZ92D
n0EBd0cHV5VxMWwGZso471Q4Jh57Bd9rmorPkL5UX4j58GuNnNJAF/CKFakTh9ypxswp0PWsSqOX
bNor7+YmgXwUK94apiH/eBvCd3FZoRf7xus7NegzmOvVvU5dM+0OeSmnorLObLzYhXokOixVGYUa
3YzD7Me6/J76WbNZgL9pHzeKu1mscArroL3RZ8wCRg5PynNgvxWBVmEeUNwQGybKxRR0g1qvHzsk
cnKPaSIcM8pidI2gsv8Nhk2hVjZCzmFOTrqQfsxy5c8g1jG/+oJRvGWVhRGW1IuD513kCSZQFuT0
fp+gWIMXqxmg+OWjk5cw5PuTqr9tVOv7huVXdEZl93NxF9Pe7tBZ+7cNRztmkmdSZa5PzXsrkf5f
lE9tvxu8KoL2ReI3CpVy7FCin/uAJchgYL+xa2B5EActq7FH6tT1AdE9GJojacVnUjFqqtUcJgm0
gqCyGbT4hrzSSTQF2Flf29ii1Ps3wVBQD2lrITjIqvQ9VhQCCyUYCAcnRzi3pL4l4BswMmIDUQ/r
H3LwQ6XsCAKF4wjTb/+HwyRTIWVOV3YwDlHy3ZMzqByKxaJlHUObVK6nu1/FGPRDR9QOxNLUuz36
pqCBF26bMuSGoD3RWTSt/9xyPE0jJVpNxvfvtx3KYCksGT8uF23rGcYlhhEfhd7H98dFS6gjAnSj
RAcFuOyXBmMx5DJ7g3kyC2q+A8FVh+Had1rOnGfELhre2GDSCVp+hKgvexNyQFAybdoPZ8dRA4Cv
HL5Lc7q7khPaDkfCt2P3ff4fpezbwyDWFxASeyL/6OnU5FtBlN0Bn67hOWtmHB2b+gJfVjAt8Gsi
oq1hNvQXm4Qh+jdU2g4xzemC7/K2kWOogigOILDLJYhcO+gLSzpPYp4yDkGGOc3G+N5URiRtDQYi
pGw+Po2xuIxNU+tjwTosDNzs9CmR5gduDlBjX9iJkPL4hh3Yj7twa4QsLwhGEdiWEzX4laCfn/Ky
Lv2/sm6slvi8TrCoEM7EeNRGzTzB+yWxe2icDDVIlODTgMpC7aQWF0GAgSyvPrNISt/YfU8vFwB0
r1TkAiRnyWt5BzKIxzfuvOi/4Sih5M8qvBKQQGLdYKdEHJqBZh3gBh9PPCa19Puj5jUfjyyKMREm
zRUMMKJ4WmhDUS2WL7I5almtW9mL5pFAwnNXfEvp1kCcrvN8ZlbHEL3QRZIkp9jk/PkgA4/QNF/r
7Mtz9552o1iJN1M5xVLPFnnpjEsd/REZZ2z3IgQSUY9OZSf87hFm/8dViMVQEnWr1gzS/VQgBete
q3qS/2uOWTYvxixw3lYR4XGUm92h6Qqvu/rtB832V7sKDiZO42pMkm2JuhUq2LUuPTX/bPZE1Aee
5O0YO8ny/PYR9/jnoVQX2WjQC3+ZK3OYJFSg3eCIWyd4s7acrgaNTeeLc5b5zFymBM0ej8EG+crX
ghv0IyY+CyYxVc+JvkKZZ8ualsfJ6dLkar7s+lMw6tVqDJlLXGylRpFmcp54B4oJ1fdASs4Iu1dZ
klo9PiU7cNIbqzIXrSfHX8mW4Kf5QM5lJGraN5zuEDLPHrHfaXBnsVTGgiIBcmYcF3YQ3SlRo34+
AHvogLTiW4E/I0C8cioNRkcS2yynhKN54av961JGPHkGnSK8Grvbb9zNFOaC3f/+YzIhwbAlc8fJ
enrKXaI/Bp189j4TdQxjRsjo/VQm2LvDOAMAP+f29aX11XQVa1VH3yq8acRV99M3CkDhaDXMccwY
vJQNfWcnKXyce42t2ujS45Hr9eqMl0OFyXh4bQ4XHaTYxJvg5wjS/iyPg2OZ5dni/DHjZLTLeZOA
xb2T26AlwV/QCc3EN/809hLiKHlMrpazvLUgNhVDlA+3plc1ydnFVIYpCFArseWtGtxWIAyTTN2r
ZA3iviNmlaRidRlItFloMkR+aeKG+ghQtIEIObTulgwSVxDQi4IX7yenQ+raU2n4Zr7T0kd6XxPg
sd+fNRIrSeUy4dje0OkEs1d5IsAtlMg7xmHcZ5rwbKikuhltJaUsOeBtczYrhjmSPlVXekX1N4Vh
McmMDX6pzldismKHZ1t7Jekt0ClCaSJgAINUErt1joFiz0qdCKXEd0uHYobT/W1vXZY0x8MKDavf
4yZJ+xRPueIC27xOY+A+z+VI4chHHhFLfdh0WSmaQku1Ab298lMm9cskXQpK6IHmgjqo6dhsCO+J
HwLACsXIRXtp5Jze+hSIKVxoCezq+wod4i+58iA/ZauDUaG4mMeiAEpZHUWRNTE8YzgoHxzLTOXZ
aTChNDq1K/SapP+eiS7V81H3KVIGGKaPyCLlhfoaEjDX0v8zrkKIsl+LlL1jP9m2KbeSRcZ0VO1W
iIG2W+vmF3QK65YRTzJl4eyOM0knorSgNAgLcMH1bJMH2T4WP6PyF/yhOg9QOKrSXEsc0VwxwkTc
5rL+R9xEPL1rDfxSjbwoU7pktFK9slMO0R2Ec1ivaA2D2KIC4PsfzkFLHfDU02TbnaTciDDM4gxY
SCwvyyEURGXCpfO0TX9JSolKERvW176VE1EVqJoEHzdQovDlo+0m6IsaOdzcIlIFqBax2yf6TUbH
Qc6R/sAjTCcpBVI0Dq4CZ/I/T8dLYIt92oMJZwxNiwl4Ukv9uhwokWbbSXBXxwNdxg70HNVAHaab
cRzWIp2ZCjsnf9ko6v7HPZN34Fx/piogjoqxQKS+SARzBISiDWmqG103OHKoXuPeCTh9rN6/MKYV
4YOvK39b3jKAJMchmhN2INUoDp5qGkD+RHymfxi6fPtVGgk6fReELfc8+fqhHkxB3F63kv/JWuav
bReFETyB24/AEP++VH9/wNWtCC37BLk8r07ci0ZtZtjqmiEic8ICyDxvBxzflF2iAe0XTVQiAhCl
5uNaOUW5ogxtQ9ptPZuuil7ofMgMMscv6o7SUTJvP8AA8qZzhYtOAL9fPvf5s8s2PqVNYShen7v/
LsTeZPTU3F23UwqS+ALz1U0GyXFS5/jIVFIVaON/2/A5AsZ7QNWihrmdGsDsJLMmuBcSE15gN2gH
3fOhrowCO++xkGybqE1+qlIu1Bz7cKHHhkEIhegD7ctDsxUM0eurgEntL4SwsqNcD9eXrtMw2tdI
mx8sSmxGxAn4KEf3m6kxgo8TW+ttAnys0w3WRVDusFRxXeG+HJjNywaeI2OxyUPryv1Gi9qSmgVI
OBOmUlyfoDPRDIPWnVjKTC3pt8QFtd1aftqnRvbu9msWUdVlD4awW7jXlpbJrjI9AJzR5zQR/43D
Xna3MpDeutvm4ALnEUKgP4Ttk0W5IFtyXpeaICRuF4u7IsTjuOEQpAMYD6KCwvcRjkq1oK/G0qZE
pkvDppeIKgkM2vEtH4KyecRpYatnsaVKcwOqKEPmPTvlrYfeq9AvFlAkpu6DGpZZLll9WxKENhro
dRJxH/jtleB93kWM/zqve7dFOAUFMEAnbNCGOq6Xtda0rHdIcKhqioVirG9HJdQXPcudEcuhpT/4
JaNbHM1TNDhNSaYYIaPFM5Jhp2ZGcpSUZxKKYaxvrttfbSCZabSA9xthoNm9K5DcBHlI0snNsM0F
mnHTJGCZtOdAZo7/45fu+paYBYG59JCNnYbceDBqPxJg8zFSPUbIQXh7aW4ft1OMmIXYnvVmKHZ2
hICyexj1ZqGXSDfmA85xqp5O0aHpsScn9zjMPEj2D9Q54Ic/rmEE21bV+tbhmBy3k6sblPibXtCO
mJX6PZS3LN1S/K+srmk4Rz16eHk7FN4Ld7yhRUNIFUbNRq92+Xn6vDLEChRJ4jEyxDt/7MHFEg+k
mGu25tIpFGnMUNU84ys6DRGrZOGJhqRCAvwKVaroujokWgI89vGwaDUE6ao4/UUGFDuzcE+UFalF
u5U+6HFZ1X/4dAaQSNqtEV/EQCY6jYPGE2m1Q5TeCpvJm4N9uQbMrVibKamsn/9Iptsgk+rJ6Kel
vcQP2+5XlSpHa++R1wSmtsHo2meUnAht2R5DHNIU7BJhoOetS9Ta9mOl8TAONErzKnu+B697c699
P6VgwtDU3sJpbQICzvRlkm4c6psUbaNO3FyROl7APuDy6BL0pcdaX+elNjrxLt4tqeydqPkaYkLC
rgnrnR41MZqI98e8Eap0Q7RJ0nQCg1ZtheQqhzfZhrRUAiaHpyUUCS0Df34OumRivykoxos4tNFY
mEuEz+s0N7GLr68b58f7YTqdSj4uDBpcEQxCT5FWF44V7siXNNKA0viiQDpNv8CF87RvqPMycSDT
0d385561HYkXEc8h0qLSi2YqfEeoTG1S/I+IDmKyz+FLFK8Uov7LVgR6M3f+AWwW/c4SdXlVUdSh
y2MGL1gpUzkpBRxhvOZrwmLqeCPMY1u9l4RsRJb1o8oo3HX8IQlvh92Vtj7zozMBzXdBQPTrIIom
DdVZ1jRfgN4ch3fCDcHuyvvpHuYXQvix57W1fG6JGDBNzFujygDAz1lmoPyNJl0gXkNi+r0dHo/d
LcViSvLgR/TYmq5E1hy7+M5cpUXnOuqbWvqCZAj371FJFugoQ+PIJzIWEd7DQ9dGPLGU896KDPKf
m5/PimgvaRRekFSphkJ9Rmpe0H9eIewcg0qYEu0luURm3qfNfzg2LdAF9gmD4NdcDe4qioVZuq50
R7CeJ1WwkW27PT2ycGPx+Xe4uvGvAQRv755gQp9FOOqmL+uASe5Ghzr1bXcgVu2rGOiqRNZx5k4L
JQk9ITvvmp072nGAuaBSWe1b3I3m5byE8vpb35ueKlZzLTag/Z0aWmOCm84RIniTBX/bMIRC11xd
DYPre1oZRIEB+4NxGz2ejJZVu44Qn9dHqQiSYrpiD1yqyIG9OPY9NO9/DenRHra9kCLt2j6gLQ8v
96g/zVl7IegNj7HpsO86ypvO9Zvog+ueWF3p1TwcEo/pO470ycdEI34mslUPTI7DBFRfXovW/IS3
5deFAAKYEUNzbu+T9U1k6zdMOUsBmRkSCZuJO0P0NYsvec9cJh2k4wTlQbIjibrBJ7jnp9rzKLEY
1bmEPNlOD9kriDU+AHEJM9YDWNcdnVGZoY8zLfZFoQk6xm/ajWI25jn28/KHyNdLeumBEwpKxasc
ZG0/nyO7GMbUT2m4tnY00b/wpACXIYtNf4UvvDeoYotCQjdLKMwrTpwiJbW3zgCVmDo1K321BlOA
AyL59eyKaOIl30VA90ADgA6FnPVYtqcdCV2ytCgRRYbD0ZEJ4YnCLud+9lyNateOGzC0EeVfhkbv
HvtDDeV8Jt0khenQ5KRjVYqVF8z92mhENwGXcbPetysUYejgD9/5VxifjPx7Xwt8YAoeIaYxiRCb
WP8GHWo6p3TA+r1u1dpv/uCjQMl93ULzTPWX9HNONvEi7CJnu5gBxL+z5ngjAQGoJYzcx1z6k2g4
zciwnQB0S/YgqymHaHVkzr7Oz711y1D56AqJfKpdO6aVg5TDQZ/5cBgv5X9Y87HyCNTUSnhSKvAl
/j8Fumc7692tYlwreKu4ZyH6MN0siXLbybrzxXYfovchDKriNLqwgfRuvRHqUUID0yNSe3hY7Tp2
c/FsA+CLXaNHJw5ABoK6/8561KdhTlqLwLni7P4s0oah9H20MJ3RDuCrdD43jLM+twikM98r/Is+
qpFqQ7WivLGYKhRzgPt4M4PhV53dkc4CITVNxfg3T7hOCfEsNQf+hhrDUiiewOFb/eyaUjSSP5n4
T9GOr/jIYUnNWIl+apwwtKzjiHIhTPI2xevBjefudFoiiagWJIvxoH0VJzWbT++PSrK+eh5kINuC
jWinhZ2FvPlZ2/SH2UgScmmkqyWt39Xw9kvrvxzUhESkDPiR7BALmwQmkYIQ5ZqEQplA3ePjG1IW
1Itr9fWJD/g8EO9PE8NHn7azaLidtHfty2VP9z6ZV0BMaKm4MJ4UMw7K9N+smIpHF7/TlFM8f5uf
iNMrkkWaTrpKPFhYWNBmsuf/jqFwt6lgKUsxlTwtFY2eJj0QLtmI+Cdi+vnUvVqNK48h3TMP/98l
+iIHugMJ8j5Zk26SfLk6/ISWIaOamU9hjF73h32g0eiW2QEKZyRpVdUZiZqxiqHrvefcPnCxVff3
EEtylsRYKNAbQNuSVCbS1oUbpcFdEJLYrthiA8IXPNU+z8YFVrcLKWHsI0VPxrkEinvKbhYi9jEg
7g3C0S0iDwU06aky/gDpWskK/vgdtsKZkM5EiImpphj3x0PYkwiP4iAlOyiIfwHSSMisa6FjQaZL
Z0WLxMYcmEuVsFGV5eJtkL51HZD2IiipzoADrLOJaGaqlCxd+psP1H/FlIMRX5f3byn/l1CNQlGt
OB/Gy0TEiHVa1gPa99qK02A1c/Sda0i7kN5GSveCqizvI8EOBlEdzZOjLg4VtH2o1ODQwwoWc+ZI
p9aSUop43MzdC+5lhPD89R4L2nMyGX4bktgUg85RaUBeLmkP+wbDAxJE1D6R9gHhUI0pyd4iV9eo
i/96X1S8cMjnJEzSV9Rp9ipDrJ56QTiyjcgZf0W6rWI1mJ9E4vQHPKYpiG6/Y27m9yd20T9sOmgL
WaHpWAF+/I8zLsaz8P3kl3BCC/CjWvCp9dj45SJG4Y8LmChcgSmL8a56A7QIdPLVbjrZjF6qAZ90
3doCM6Ctimj/1nKh9HQRg6rWRn7yLS2NkPckxxlluGxVhe+xOiBaezr2XN7S87VWs6d/KWaN+K3h
mgQpj+UkEA6pvhO/XtJuTfnl5AYMQANCrzWaA3pQ6FJ/kC/fObXJaaQ2e715n6EzKcGPHoyTprck
KSU7o6Y1KgNhSHeKCXtagKTiGj8O/UsAMPNFb0YpP0L3BqaRfK1oa1pi40zqkgXjlP3JW3kdvRxy
4lXRo+DqgAiPlmJQ94u/flo3xc78Eg8ym9hQ6ADvrpuGJukJgZwMIhj4trliADUXQdxZZelDK2Bc
ocmC65bAStyN5WJWeucM2pSJHLPaPqHig3YYnp1z0R3m5q522TDyv3cSYtpdcpbNrgU4WFicLEJw
wTJqOkbK4nG9bJN2C9IoqYps3ojyOHGQcQ/3UUvbgHQDwp1SyD9V1Z9gFBA7DaIpPqMh1VA+P+zg
dI8+BTt+qAINWo0tJDjhj5XLfCrSrM+5hBVm0C2U+vb1XclR8QmV9A6H8NHPUQ9l7bPeCGMtitfb
rJuaQ9vinXskWMStHa0LypigLsfjiJuJOk35UBkFCrD8y+PAXKnGOZuWTfb4pmd/1mIPA7Z4po92
BZtNN3eRVnk56Me3Q4RYJ8+0v1ZtnchP7fj79tyle1eXp+EEOWD/9vh4DVLiGM7JzJAnFMap9h9n
pXa7RRxEzmzxf3Kql/nS10FesUaNrJCW1BW3Y8vffmfhNGvAqQ+TS5+MyHA3uk+b6Sa3oI4YyLll
luIqtZw1P6cepFeEB7YQkvFAk+KBlo8xPk1WWWjGRwfFh3wbK3x7Byu0QjplEGuba4xa1Z2OJHGV
SWmuBA7J/oddvDPs5Gkz62pq6lHSEj66P+/nS0aj9hPljVy3fgDnYS/MUM6sUJWIKl2524nY6X60
F2ZX6tTm+IMv1kjLtUR7zSHSC3OTAJ0CWaXHuQ5scUPFYs8C4ord/RAihjwPt7X5PktmPahQP/eJ
lP+qnBMZdiGXWB/qFMuWicxBsimfOhN0C6VtvnvFo/g8+akHO/K7BmvVs57Bq17hWnUNT7jP2XJw
oyaMH+Mo+wmtj3cR7/I2tP4gK4RlMkpNQd6PIuEIuQ1atCmBz0ZewKQG0YexUFtSSEcj545yXsG6
dxFwVS1MxFYQP0ogyMRYCZGDNogeAj1jHi24hMOiH9jJkXhx+aHok7B3Aj/d8Jxf7thka8NiFul4
vqIVo7NPlPlR7QBsN3qX516kcuHI1Ci/TOqG5cWklQbJRYSVbAA/QRJCluV7xI8GpXzQbhuKxVPo
K7K/gNZmgSh/RNAgs1t2wxpa8KNY3/6R4cIEkNY3Drr5CJ8HPTXOCP2uGjhh/ZhqaEi9YH7Z85EJ
AIVRkF9ZwQm/tEOQyrM+5Pg+i1jpsom0HcqtY+zB/UYVq4Do4UWkLooq322boXm8wgoholYtGXDC
TbL6Ipqz428rsruZOmRYFsjl3URYmnpbXYVMKdI6dSkm9UA0iS3mfK1D1tB+t32Ie1J7AjSKgwNO
zcLyV1j+KABhIGzqNMiGPIy0mEQYzLbcl3kFA2w6uylFlxfqenrNuirDC9exMJSxjww1v6o+DUF4
dRdig0ExoantkYLFjb/8asQpjDczjPs2DO/6jqNgMqR9CPS4Aa3pWz14KfocqZ5BeRQ+xFm2oZ1E
w17MZe+DjfYLxXM6O5qJk4UEAgrz3ZhzDxCRj7S+K0ex7HK0/RZ5Z/efTW1ErWYKtq927Rv3FHyw
5qNXGwPqa1KscN55veUhUFql+FXhVygRdWI63i+5ijtAfqYVMvsmnVslf41KRur8/vKXcIdmfRE8
cjj0V/6zs4bfNJQnPG6sx+1dUQkkfr00tEB3jUBMYFgsdZoAJ2Pd8KDqUZ88Xg7+bZjlp0Z/ku7/
ScXg1JdwAgT+BP11kBwFtNAcrQ/AHUbIvkT+j6X4Hqs8lTw9KXuUFWWuK+BAS9ri0zHu+XlGnJ1+
D/qEzrECjOPHDqFlwuax4UcVtjpZzMul5alDgly7/6nXCt7sVoprcblyw8XYAuIyGaTjd4oe1bCe
WvGTERjyEWXEUlsIYC3QmRRbWAp6XcX+LF/YuhGNIERpIe3+3SvZYQslDd6Z2hdaCgYuqPBSYVVm
9Mx1lVd3lramEnOdw6i1NapCeQTssq9GT8wzOtWyBsUtQo9Qr1HxoG9YF1OHZCG4zALTGVaBXuxG
BMhmyhSNQkFyErJ1n1EmEOt0SobIVQpkRPBpGZaY9zi/Hnd9Y//qpuMOHmZ/KbQj9lwq4RO5JYxx
X/HsyEarUjbLPGiAFgmk6Q+IUbwAdSBgJ9jLlxgQoR0W6rOD0Uea+iE7mXFDTH5F0qt6bCqF9faD
kjqoXjLvfUpCTyueyMqeaEQ5tWg/WDW4TMQLmYpU+VpOYKC1ydEt9hE7QlMk91uiJ9mDir82YtBE
1hE4dkeezdAVfl/MH4sIrxcjxd1F/Mf2E/V4guPGzQ9mn1Dc5al4p7UeMdEYwMmD5y9U7TB3r3Jv
u7oBXwYdhaKvqu3DgwMs0p6c3Rw5eZBDUbC7COdFd6XLgwAauXqlYWk+Lhus+vuuM3yFeNMV4dZf
2KMJJaLhrmw7f4no1mtTtWnDdfI6BlmL8Ce7eBdiTpIjLwXA94OvRwvTbWBrB+mhRpU1vWjaiA82
lQHMPA3ZchFeWFE2sSLu6GO3yhOCyqxZCg/L1Z7GslEmRl7jFXw51q3FNyPdTVehbrfOBqI/dsAU
b20A7XC+hQFW7cF1ArX16A1agid81TSSASF5YQRDtf5+AZjhIZBgaps84RwgOhNENYLJStkWm3g8
BOTQXzLbGeo+bC0DpuIZwdIDOZH9o4H8ZKqDUBX0eiEGlHkp3nw3IxfKLAyrStJnh43cxS+g+i0V
KHNABNkwWiY4i06PSyTnWfleiVXY1HktBjW00oyG+/iUzSDz33tf/CC31C/KN0Fb5YJ0x4QNvoKi
rw79VAgZP+Y0Si2HXtqwQDQnU3JK7Q0tPi2U1XVsSDpMwPvYxTndY1Qf3jfx6RiWdwkjnUuy45K9
f122XeSznzHKHpvlYdWx0b1opXVhCo/31jebqtOS0Nozo0aPhz9+KzB8X5b4rhmE14XTVna+IB5s
QZMrY7OTpkcg6hLCns4CFRHRMGKc5gNqek3NnW76Xoe6rUQi1kUJ5E6vLoKZbxGgSfgYiuyHpfhc
u0HYWpfiJp2as9yGe4tk7U1ymdlgMyePGG/K4MeiIa675wm9OYy/FG4BD/MFjUsLlhZLO1A57SyQ
I4q3sa4OuM4aEL8uWecmFKCotalK6+ya/gBLC8lKlnit2ESXGi1bCNuTqQf0PRpXtczvv3WlF4ry
9G/VPAlTZh4WGBLUqgUdO5+cBdblHiXjI26yYLsofQzb/c644Is2ppCXv4m81nCwvVDzlWBoQ1gL
tha7HjP31tw1Fpj3TE4663w+erG5yw4NFY8oPyk2HmkhAK+XUUy7067yi6CWzE1csxyRoXegidal
qRf5Gg7emYhguoeDUVEwfoceRQ9YOpJYxY8gGwr21AH5Cuapnsrkk68+Yc8/bi6Jl4ajuDbyWnFi
9e8AxZmV/9vsl9ABAfCgvPj22Ac6+Rt/vZPiUiK0GhPn2O7XI0hAa0j+qxx5xaYF6NsR6HJLehFn
2GSqOs64w++4LYL1D/TdfHKnYFwM43U8nfBjifcsTVrF1cmPY6cmPZU4t5nd3yat9cv+Uvd3ArAa
Rm+SrzMqYlwJz0FdC46QcThCM0ebmV3O7uK2DZdgJMrTpG/TzC1UuBBUPCB+d4LBD1Fo2g8cbN5u
DB/uwk6Kng0hxNztgtpbIipvziWFts08DScJPNjanat3YFQp7YvBjT2vFEoPYIEQvOUY0T6RHOT2
J10VxUIPmdPVEiTFMj9x0CtLiWctgG4EWnYb6XpPZyXqva+eKYW3/phEvoVkryJf9PGQByJl9qFw
34FBuC2QlkViUuix1QY33f7Omf1B6JVYcP2xgaWn4gUD44oRQnnjfUTH8AENhs2QVx4yl99ZzwtH
pQIxiHRVI+p+yR1SYAr1XeXgDetX0ITSM5sbUb7t7JrK7vdFsvUGWsSilf5YpwR5V9En6nH9SqPi
8v3wTCR4TytyqcP9oM6wfp0pMIFgYy+HAVLRPdAhDKce+OpiNGr8zBybkn/rbsUaWNL6Y7rpVlCs
PfAhwmzuTXkq7NN2buUW9JEJYr9OnTTd++OzFbfs/s81G65Rvwx9ffUjlA9HOzHeU3waSL7B2F2U
2Uq8clDGwDf8/x6b6oMVDtGCkdr6Y3YpxmQoKRkCCDlaeXllsU9+PeKukYFPQ1To89yPxSLiRPJU
cFE3BVtkLCLKwwxYPX668/BeWPLVzgkzfpuju2ZW/BtpEZAHtqz5E/Rm0EWl2OCYd9DojT+N/tJE
5hTmiyAgVhdc9GcNnPQ5gGPCSH45fiRfuX3rpl+NSmgEgzxX4VBxM/hGRhLhWOyg+CxnYErn91D8
vZb3ZFmIaqjE/VcaedolPw4yUVaY22DwK0yOzYdbqSKnCOdEibmM5X9cHlgXq3waG/wqXLsxKD81
RifeBe49vRVGuaMTu8UO+XrnyabnCHu3ZLAQBGR+q33fqz8hJBLQindKzUXkrjUqWUWzwbYXmqpZ
L8wRaDafv+ma0wMATXB+l0oCpYmO+kbC8PHs13Gi53/gCmJMc+MIeFsJsDniDYtrhMGxYPtKJVy9
Juy/7oy0heX9QC5lmhCDOGi8a9rdYvVRHJbqkU8w8AfvUyvqkfAAxItX6+ciXODXwal9AktvFzRu
cy4LHwwq+bjAyTZRDPl8n/tLChjntsL3WfPAkB5Qq4BbXjduT1pzdVVZRvEdIwSMovB8oCovFhnQ
NZlqtUsCSa4Pga0zkrTkn/hqiC66WS5q9PH13oHxvfnIWVtGNzmsOu3x4/gf3emhy31lRYC00DjA
Td+67lF1+Mb4WJ/04qfUJbJYLX9b4fxzGkNzpq3/38/Q5yPN9lU/F2y01mVacGz2cND7ZK9Slsxl
GPXxrIr5RCXv67X8FknjyIU6hRQl8Kn85Fe8HW65cAqzla9iSOwQeod4czuZTaD/VJE49ZmJZGxP
JRg3FfozZJf042vgxkGejkrtxpTKLhEqLwdLa9E4I9yAV0RlOGqOf+b1eEojx93TtA+Qzfn1r7VP
V44ZNG2zeszinK8czOLScnRwCHo3G6TzKSQqsr7Rf0IXYegCWwUmrNrutqwji/Lc00QP61YFBHTK
LFGNcEmyrQSVnxTOxX40qbGz8sPIo7A+giNrgZT0jtj5ba8Rg0m5eZWkjkx7VORWEsO2WWat+DBH
aiA9kwyWY72Ingt2WDFcezawKFy2l/2MV+zonctwO1lkbuywUcdRktTZL75cfOC2sOWh0gzy8nsF
ymwkraBu8iXX3+vbpe43DTmx/9qO9OoSnal3gYN08vlKVeHZHdympi4SbSYH4uua9nhxmcUpZwux
Z/b4gEg/KmcqQmPTrzZ49lskJZ+x28llAnHDRvHUa1wJFiPG++rK8lM7IwViTjjDo5CXl8ymbXCd
g/3oOnCX+6E+7JMhMSNrrDHLAdS7alerW1xn1o/0P1l0OrVUsA+R5a1n5mLIz6o+9cZN0knQqx39
kwEUBiohgIHdBc6gsAZg/k2IQ2hxXg2nlIOx9/swViV/YRP+s1ztolOjCufK9FaCvs79IeH/cILi
ZvE7GY/uyggcgnAzF/mguoRZdNsYUnPY6Gge4zRfrS+MvqLrXDWeWAXMXkXYGGUHlMhWc07FsNrE
IkLBd6/RB/QcWh6jiIxXTy8EzhA9GjCN1IqXHTSEmT2572dX0bttaygkV3Z0Hvx37qqxM5HKLg1e
sIesW8jLyoQYAS03rbFzuS4W92c52xa8N/GKYf57OMHCeBkC2RnFmk2WKBPIm2lL26gU7dCj1A9f
tS8rN42I9BVgJHuI/BlJWbcdqt66Vrm9S5Gsio9BjoagqdXybML0R2Vb89KHTdNivRf0XS59+Cp8
7jvbSg+WKoTeYegk4DjbVAXO0o8M8RW+Z2WN4ShuX7O4Q9w8aOx3aDzYwz9rjCRus8dppzfT386O
0rVYX7uaZEmfMcTbKtXsAM0A29sI95kTpg2NlQJg+0cR2/o0jL/py8EPa/Co07dsyUTt5VoqXULS
tMdPGP5zLA7UjTQHqCf/iA6AcOPPMA/UdmqphzqjsWgsOm31Spt0//2r69wN4OsvWeGyKuVnWbUL
bz60PcQ136O2VkvqypdwXUiLq//LHBAs/GYqZus9Aldu8I027nEg7yZWTF4RODnFxi0QNVnnIiNn
saRrERosSlKhdrDw7Lg/lZwe+nmZ9H9B0yUgqiwGWsnml8qyF5W/fxIvdl8BzpH02GT0pE+8HD+3
9a0Lj4H5VSMstj9R3nbP7cxdgXeTk0ZnBDJQRIHOJN8yDt6zHPmuR5aN6ZNsFpcB2eoKA9pM9w45
D9+bn6CXi1zBQPzivb877rg4sliXF7zAYwzvDIhR+Pi/iSKw7LQH82abNXqgCc3Q7rl9wOGDwvg4
dXqDqW+ETNy7XisgheSUgBKLeCqcr7pAWHMoI89gBaSRAUZQlBS73r1ZDrHU6GVeoX7yigsYN6ch
TPPRmJYPLKLLJXFiVmhBvk4v1891C57ZcX1a4pM2ZqJGpbZp5UEbhndCMkAUEA/zxeFRTVR9mDm2
BuHeYJC/YH4wpzKnGs8cly7rcul3j1X5IbN/jwfOcEELooCGxP4VhEwqm6ii9EM6iQPbCN3lVaUh
71q2cOYNjut5n5tHHNL4hhI3zt1TUKHomwgJpAAnsyaUR4u3mWlUmJ4PRuyW/WvJUexdvAbpkPii
TJvY0YaDySmv4HcYvouQcwQxXIO4Vnzts54ThnTVRXh6/nB1fpWvP1pz8RRpma7n3RMEsZ5wi3tP
LX7yD7sziXCvsg9/DqpzNYfkwUCxsZ4BNqiOqO8yV3QUzzyuN3qe5TXHMxelDextlqxbHSG9s9Ng
P+RRj+0f4det8v0H8qXc508TNs4StKuYl83kuWdj80JBeq+kThiFUEPmkB7T7p8iCb4zWRlOW10t
XznPzmZOlnN54rf0CltMf2jtmrTg9QtE3pUl5erNb27Xqb+htUaNxxKFxDzJu7SUTsOuLDNuL+wU
clqNKrTA6y8cI/J09PNzWQKxxkqsn3i1qqkYhRZ21Gm/f3S1UN2GOdriSnkMDC40djTJMs/IFAtz
KriXU6jNY2uVRxfWCOcMr2aQir1xeGDoZU2MFdndn+2YTiK+VHqXhvAhlPKhbDY4Gq12XOR6Bibl
Mj8egxa1J1IUjM5nuQdW+m3dZHXcV5+1iKia83ZeMRrXDu7syIIC5Ale2OGWQPNu0Wb5iobAE18e
/PdHXc8PwsnfVguEhK2Ja1qVD7K7BHObdu3E1e9oitblrWJolllRsZ8J/H+ok3hPjSJZna3hNAmu
RQUKyYLhvZrEHYtTOmgXRC16HbDLXUyArYmywplARi36uq0l+UVuqLOuYhHol8DVDIWbQM7Sfamr
JYGcl13Lk+s7zhs83MM49iQPHltAJSe+ntjrX5LmZwHuaicha0Azlrh19rgG7XFn6YCYVQ4BX+QE
XDghe6Km3L6UgNHYda4vNEk4b1pDJOxaliwJK/rNMKq5LL/M4+rPdWMLiTASfg7i6+CHTaDAQagA
EUWiTnLiZ2YjBjf1d/Xk8Z2afs2l+PW+EsCZuWa0uVHRw3nhmW+b11fXhKQv7rujadskHMR+ULOp
SeUHvIP0V7zlIpGYOD+Hn7WWe6j7napp1dcExdzAimMoGW7Jdx4a8UgYff+1Q88yt0XPZCdDA/6I
O0JtvR+QSfMwrfPDDmDZyh9JgOEB9Nujbzo8z2duQ/+xNeSSk/ZEOymMgdD6+WKUVLxU2vhrFg36
C26H0sHcJMNVj2A4wHgeAD5uuU5ZC+oCxClHOpF2OGNdqazKWDA6MQXHe8/jwV+NeOYVhpGrHAxW
Vi5ILooT00mnia1hMpM46+h0QlPdIEjz4f04n8BXMHSUt5wjSQwPVgoe3YvCgfFIrGZ6t5OQyeI7
y41k3APYOxzItohWa5t1VcQniY/tIHZknlZ3yApKS+UJ0IYx9bZSeTJTXS0RUNEKG92Ob0z/QIuD
Fta7Vzygdm8ml4xRWwLvFBMeMf/+HqXL5pWnp8HFpr5JBKIijE6JnXVdVcacoqd3LrZpDfGWmSjP
q0n23Mh1xlR94azfrL/eKi4j0gW1mka1kOq9jJp2AswN1UAWhoOhHsx3a2fx7ApX5KgXqN92BZO6
+Shnu8Fz7uZ5VoVHvY6sJkROFMmoCfzhM5rLKtErqYshhED2wcwGEWSN25+J+Or1BQcw2spyuVz3
PQswDb5pz5w4D/KrZ8rh0fP5atd0jBszBI2bBW/IF1qWNFC6+3J44putyVX5O9Rc+mkCGNYmUrI6
g1MFFVQehfCa6KT9k78zZeauCy7DbehXTehPfNUpbLZ5uF+wb3SRcXIsWNJi6OLKtxaq8QIq2yk+
fvgIvhOrHG1H2MkX9wWvn770rHHRE/7FnXv6at7Dz1v0WEkfg2ymSfQaNw6k3nfzfmE4bNO8eQPF
D46l5l32Mm3KjJoo817cTWozHwVsiUoS2hTngR+slHg8yq/tkZGvX5u6WpBvj6cHyo6RJ5mXaDKS
ymhCL0NPcy6PH/nPppQuYJN0XTK2V1mZRvdNXrn0cVAoexyplhKwHw2CnZicJy+oGwQituquOUxl
d+4RhDp+/o+8Ql2dDv+AVZEFYrSg3hoUt2FGPd7hAI00q11yHxUiAqwZmCXTM++ampo1bI3xHORw
7wAwmIsgiSlYJ1LIFAhsU0RIVCblIXL3yYU0ntRXoZJ3MP2BK/ZqcPlI6i1z0Yq3E6DdIYPNIr7Z
Rd6FrxDvXtGwAo/AqKe5xNwtgoV9WoLaT5/jEyvYOAkBpr7RkLyefjzrz4EQtm+OcIMg0jalpagU
YKo3dvm0NnBsAvD92q8tWXioMkE7XcPf/uWgojnCetFO/nvMkQCHd6CKwsdEpgJal7x+0sGt5heV
0fchkqd6FcBN/MIyVD+Qtf+svRYkkoAqxp+Phoq9wSuG9ncxxB8JgvGEpxNIekYi/WvOQL4MmcCS
AmKh7rX/zzoaGT4AwY5CJS8yXEgz3QQ3FVaLzNFbhfA/UjnfSirVWyujOuz4Qh3oux7FSUauKOk2
Y7XoRYTzDL7o10Pcm0ZcmIXHfE6JsbRgRp2mAGOwdTu7IfjsCE55IBDcQB1tQCK7nCSV7ipIKITL
AQBLW4ljSH7lsNY/co8+KtDMcbcZRKyCQfgZC1/CFBMQpCjLyu88E6gg+uGLjjlABNiwbeky5K6r
FTYMYlM2Yx2Ruqy7JwtiHN6kVnOWBabNjdaQZGtQOxhliSv/iUwPpq4SEiASdFP6hDUhYx6OYZpn
4wQov+qewh0FH8NtcEVw4+Ld/wvzVqXSrnHS6yK280Wb6vRiFTCT61lNnurxfFES6A2GH1EaEtD4
2/QbCZXrqD2oZ8whg3Q/TpWJGir9YQO0e21ThY++sOkguTO6JTV3WMUxhpf+RF1MNMlW9vFZNXtZ
TWNyGZ2vO8vt16Qkk5iacXnj90RanNsqLUN/XS9d3T4n0OrPy2pAcnwUxv11/pZZC5iMT2MGrnzs
nwUpVoy+itiGIK2RAsTlcAEyCIVlGozr385CtLO4kj2naLVC03XQgcr57y4hxwyWzEW3vzsV/K/P
W8XdiJxO0nbO7dlqr+PeSgLWZmbtNRdppWBmNB0fm78PawEmDooTTefybh+u6xKW2In7ayJHVid6
q4J0FwT4C6AeT/yEIb5ofhJH8AZ7IdjX9L55rlhxOUsVZChBTECp9KOlgkxrijxeVGvYvFPDDj3D
o7ASOIbFQZG7Bnv7BpEW06glOMfy+na90vJUuO2EMPg9GAMgkegf61Igt9IcsuW4/LUx+n0yVTnE
uyDt5zyP1JgdVNUlEUMGSTnP040/ZF7hOLHJROFgUV8btLlu2SajIhvr3UNjM8Ngr1MiJsCtPSnL
YU7+9qUIRvtFLDsVpUzIENg4FSxVCpDJ6rfn2pnAlgplodVsNvzHTbOOTfJ+gBQqNU7zOJ+vmm9G
F6Rb9odP8eJSvvix+7lVzbDpQu98AB2RLXg9dyPLUf0FnshWIRtr63SM1V01orKbS3nnMZikOTzo
Gu218sCPFvlt1xwtFgVzLyMZ9zFcImKofRghWAcJp3m18Tt6bB5UHsK0oaU7uIBTZUfPu8ghO5sg
kUjnaw3KcRrdFlr2KnY6V02y4cKlSvxt4nzuP4J2aqejK+KA0CFhLJ8mUKvtJlOdRV0gNWD/lgFB
gbT7UslMtVP/Y+EAtSnp+rZiI2Khh01lhfBd+HzcW1bqiFRebB5J0ws6f5HlFiQfSRU+5b1BQu+1
XmBaIy53zqUg8OA+sKFikcOv0ikjayo6AqoA74B1bexPtkqLSS56X6DzhOSIUftmaK34sJOUFXOB
6sa4z2PLjf42frjnDBEwZ4Yydvp8mRIE2EW7EJNvDXBiJj29cmv8RKCH5mn4UcveVhVhP55lGI7K
in2SJqcmQ0UmUeXrP2zn+Wssyujm+lJ7eM8KCLxR0qIp5gajpqGCh7+OUsT3VOq6N0MD/cod9Coy
h5bzYeFhr7ptjaYjORMGCy4rvRO9IRiGKw8kZigAYJkceziTau3r+CBTK7LPePoDv2bXl01VudXa
F5sVdYCytDsbzW/ox8want7smz7SR1jkovsgaVcp73KFfHQ17gnTdfwC2HI2ax+P+xNW/lZvC7aI
0jgEP0IFu0b4tx+esWPEoij2m/pAbUnpe/mNktPnDY0h2Uds1pFiZAOLqETLfl9pKtfVYYkpNo+J
6ZleM2mb9F8C5BoUTMvLrlC4ZsP4UFgxbpwUKa31vPH19PwuK4FeZmcQBj8wqlU130lHnnE3pjwY
xnp+0tX+VTZX516bvrVTcKeosp+8Z9RFzJV1jS8HAbY74eFhlIqgWLkva7oWrDT1fGvZBt6aM2to
OACNQB2xYgPfiHTguimQAHSIr8qJb+6aSJp/oZgUsdaBdXrkOW0eSQAZoyOvW8aVKDZmIbgM0VPl
6+wPyxMeW5BRRpqPnjrzWknEa4mMQ+iystZ9HtMQglyDV7th1qr6vGjyw1U7sQlu46hJOe2ziwPA
0TuY4H6fil19KpVPN8/x5jPBF3rTb53NvfhEgSp5nzwst8c1PaUP1y7ECxLBNKu5QjD6vUH8M26n
3BBMb9wBKareIdf0X4X+0PObnbCIU5nG/XTKuaQxJ93Vy7+ENwwh1/4C3maGl7OBouiO7N1RQwEl
Jw9MQfI+TETlt5ocG3mLbIcCRCeRAgYjCHHRryaAA3CqCqStb49EyGAEu3ZBSYKmo1hNpFvU7z79
dNCpfE/aOUSY8k7LStWiiQS0OfK29yA9gVzLkwlwPb6SDx+HTyt34kJdydFzQQJhYY3RMWIMYuJ7
MxozdJ4mmSHKEkeimWdB2B6sW/qcDU4C1cMmVL+0I+/dDtFEwnIZuqhdueGipl8PokDtLKlriUKl
CK4kecOvsl45Sq69SKS5knV2aifAvE0BpmIz09s4sMcZDYuEYp5EONs+U6XPjPigJymcxhs5Erxh
HHgPjTL7ApRmI3Bkr2ts1yBKR4Y6BRnZ6xCjo23TjnakYpvxQc0DoX4rq/Uel6oy8h2UwL1P5IQU
4uxi330rmW8eQ96X1Gx27W1tuW8JRpPselJ5rdjD0FyHIs7nkHgpZVwhhmUG7vdHh5Am5mVIB0Ud
zmAyjtUG3AXoor4La4ddC7E2p4zHJGdQ0knFZzG/odnoU723+WORqqyLi663+bL7pq7kNSSE2MB4
PSjLpzkGJa0wlUpri1qZqag+cxOta4L2FbUxsEJWnQPSshsjTdwXl8bwJLYEurDM63SVkD6+D8nO
DiAD0qObMqRDzu9zstndScmkajZG0J/hs3F3LQDbVKRM8oQsK/ZpJWPVD8wBQBByJXiKkFulgFt6
OF2dW3d2/EBF61AtO7onIeil7tB1GCjszlICbWQ0rw6lgJjrLShg5zdVo2p1Pngt3HyILR3Fgpul
+1IcGUgt1vf5HjbzPlgpG2ZE9GWPQKedcO2k6VDWL1AUR7agieWL/HkYnBcG+8LSj/Hh5GdJem5y
g8odjX+VOmCUL3MFtFC82em9OJkjJgp1BjEJfVAxJ1OdpgV0u+aRdQjjO0DkIbftvhLxKtzbahgJ
NcPZH5HnWaJ5vyPC3Ilf2ZaYB2C+8WoqISKzBpoehYZ5Nm4ooBzMOk/wQRD2Ff2oEOe1DtDLn/Oy
KwBV8yfqQuGXHA4dztwt807kdzxb9LFDd0sIcm+yPmBwQzE/FXjlaqJOQ6FDzjO65MrYSbqw6oFZ
sPacmv2MTFwpnmepRI2lvEVuUyMJmzNzyE+6jzmKLjbvfUubyEj7aGnd4X5eFXgob0DwTJ26/AJn
qWwYnxhpeASkPJozAOWgU3k/7uTbg4/61m7x23/H/WkksiOA64sOUsJE48CE3ZxM8VsPADtfr6J4
cBPKDDhi7BxZc7ziKZj4af1dhlHdWSiD2SeQNkQZ/dgUK0vRmGpat34053XT3bkbL/4TNvZdB5Pl
hJVDsW0qaK6qyACjcAgXACYadcH9by4OGRtAD8cyD25Nsk5nwkBc0+jma6dT+2jL8JvxxPoDOoSE
rNFJzn1sixaODUVjBYWp+No690Bfu/qdq0ntTW4DHRAtwOiC0qyOO20+NDUh3TsPLnZUtiTmQLL/
dHu9W4k3Y/P5YDobIwunnHcu3yNtAAzd/+DpSm1KcBPELdt8Qz1XBUup85PvRaIdizlb3F0PeAVG
C9x0IzAbVV0xssuwkNkqT9GZUxrTPNRlhx4emOllSVoAftZ1F5dqBznPnJfzTKIxJIGP9148wRkA
Jq/yati5Wh8t3+pc3fyVVTNjpSEn53ZvoW8+Digzbpa+JMCW5VeQ/l7X2hrIwYrGQGN+10L/3RfO
v4EZpeXpXmk6640CAK2X1rRjimcZrupnbSmTSNQ6a+oFZxrhLzmg/qIQc5TfGQ02luLZ9nBWJOxf
tDb/WmSvfGd1IK5EOvqBUmi66HSXP9wEfAciTbTbjB5gDx7arAGNW3xHcQL+ZFWlq2nulkHUmubU
0zm4Y5oK4HSxJ6cIPW2KVyu1doGtKYR5sZSt9qB8Tz2+tEk8PYclZ5hzwGCEISGzRFxFED67SVvW
ZnybPEXNhKI90DO2NgaKjN0oBppf700az3jtpAxKVcBqoHzJahD5af1iAAbggMNxHBslMg3OUyN0
cX9skvFZPMnyH8lijMM69RKuNd30t2fR8yyh62S2spKmKqFPEHkIGQ32WPlTT8ZoXLswPdqiNrZK
Hi3rQfUfOYJ5FDOTAn3BXbyYAG6n4gf60pTXywUH4505cdYab7kDbkV+/krF9Kr2qWU0JhmrFSFd
IWXmenz3BRBB6nP96otrHLwGVL39OAE1BsI47H3D0NJ9ftK60GgjVykmkEINjJklGRBFQ9i4K/9Z
6m7Z+bEaH6Fh9jQiSMdIWBUflQ9pvkgqN4qrEs0cxxu9sXwqi+0UnC++7np2Olk5RsJizHAIM/Mf
HOYWKPKburZrNPuS/0E+evng5dZziwJ+9nwZXdZzvf1ZVlNG3ru9pytMJBoKo/IqMz1Gkd8mJAzP
rSkKsbGg/inxSTLOVl8D7SaXQh5/fuKqEoilcu1Y7zFyiyfwtQRnxFo5S3pHKkq+FxWiKBKJg+8k
scsGyOswda6P+jRg3Tp9NvA1YXVNB5KOaWUvFc1BVhx0WtoGmDFrdMozIIp+EigUOx2UElXSQAI3
XwPPd34dzWAinUygLzxF2jBlrtXP+a9mSb8kYqTFaDKYDNWn0vA6zjhCZLbMntSEn2nIqrAMJOBY
13NmDrvVslj8wfhC+duqo0VYk73J0YKiq3krN/qktN6vOASjYhTKYVpRXMY2yb48GfXT9PlEduHr
Z+HPTpEmol5Y+pcuI/vhzRdccb1NRWqHtFWXgnE4oSIiiAitQTktIKmk1YhxRVNVazTexb9bSHf6
nlSceThIwRUjnrPFC1Ac2+ry88K4JZMej8+fYX5yypP5y7TKCEiCVrB72zlvhx2kY3M2+rad+it7
jT6H/I90GAS4ybJiTcQCHrQ5GOWomL8yCpD47+rsNRldzmyKtgdJqgoiRBHoi+OHDvxaC945avlC
Su0g/Tx0Hszb9LKr+BO9DufgE1V4rgKiAz7mJuQdMSxpghMbvpJLuLufQd1TSdBRaBIpMQsEG4gj
xv5wfJ/wDVcTpg+ttMSksZ7ltx3dMOLZGl3RdzPMJraSUc3rj6UXzdQNrnHZip1xUWcnbqbJXfKs
VnWdJoJhBTtsx/9pWL1NdARTkxyqtPjQkhRMdJ8bcvGX1GJzWgw9pLhKvt53nk3EORJkchTQHbj6
90juRJK/wrUNeUsuNsSiGwUIryxvvG6/ClqMvhjtXFO2t2jTPX5MwRWHVL1hJxPIM0cFhDX8KtDH
FYZGPRD8B0ERpfwzOojtaGgVV0N9vyz+ttt7gFisGp/MULpm4BcjpGgmuwPoNoJZ/Qtttu+ksSfK
sm2E6sPyI/nydRJKyWDtgMIH4nGJchVJp5oms+rVm8KyDGbxHp1rMJsDiBm9AEggoMcmmzQo3vs+
US9u22gsRSGUcGebURtRsARySSdY7e1HUJZAN+wffPtrD9jIkb/nJDSuWYgR2LGWbc9xFi8/GawY
dMQVLwqo0AVDacAYZZfWeoNqT4Oc8cjODLZF4KPA8g7HoLUChxEnSKIv9pXuS/Qwk8h1s04psfLu
1Z+HjwNc0TTV/K4eZKQCcDgcccJcCVZa22thc0d0uhOYOPevu8s2lTSFDSQS5PI7EBagfQMVsdFJ
0w37/MzHBf2aIlwyo54zZGthROPyCwexUzPzv+1RuuNyxTWVyKLRaZbk+S/XCg6bZwgSydi78pVl
toqkKkp4GWAfRZv5ajrbMdLUq+xWgntxUw5qn8k4hVwrNSRUwsNRLjvP2ed1F3Y/ksOWNTtcQofZ
Uq2HjBGeOR+UHXqdKx4yTP6qmr9mxVxARiAvUOGUhDPrDabvsy3FVAFdy6G43zJ1d7otTRytBnaI
kbcBk4KekhS3x+kN6KvPMbT+dc7ALVvk3RJGkYqrputfgiPHHSeEaSJxm6q5s+8ZKoUm9Wp53Du0
3LcL+aU18k2J9oJG9pGLnqo4Yl6aaMR+dV4hRboYgIHm0hePCZ9PJEwx72XKsey/yW2GorXPicDg
CELfcRyx3i/+6wA53wJRBUIZYAXKahuS1YU02BW64iCAc4Qqq/mn2wtMk6n5BDoa9PJ4deMPCtEz
R4pd90xH0FdWgPuanuLNpYnkKQCJ9WqGtY774wXEqJqwCWF3VpdOrAnYDioxiQzQwgAroYboZQXF
O+oH5g3yl53K+DMZlmKD/yRvmyUIiMgz0lXtqJ1/O0QAp4LVN6PdStdyzSm9DkGzq8l6AakRGVPv
P+VZW/Ds5JSWG0JASPH7h9GoizdCP+k65vR5yfY0RBYcTaPQTCTqvEcAUsFL9IRQRZb7jYNRIzE8
dhePDYOKzSZJ8Ewbg+kwbkArPgGNNIZxo0l9esnTXCJvOCs2fItLAL1tCBanBfVI8+8w56Rimo9x
+lWlX0/Rv4L2kxh8y5YgeylPiwtPoykBhmuYGAZLo7Yn/T2OPnxEyJhDXF4xg1xp3YFCvaxkw22g
3i6kZpAqbh3cV4Z90qTqP3sB4TtFfbnlmh3zkxESEhDVeJNZbjrrjCYJnkiJkO2wcY/fBZkmcOZH
F0LjXQ05n4g9X2VZgjRrF0ngiXSDgFAImJDTb7bY4O9ef3HZOq+B5KebybSq7I+fkusuCpcJL/eB
4xJgGpDO1gMgVnCW65JKJAKrouPBNUQoUHk4uxrAMzYOnpnVnS7vkjdhWBksvuBtav0PC/yLvN5N
JBW9DVjV6YfLk05QNgM/vvsV9ZkcZbQqQr8ZeipepkPoLDsaBDZMdzARZs6AFuWsDywEhLvmVuBR
jaCPjbpSCVjVtd0qxOsKffVhNQKLFoOHvcAMX0XXgdnagZb3xJGvOXuHf/GyIVoQYQu+Mo0GcpOw
weMPw8c1UNdGVQjfk5kbwBsp8PnBryxP9ooOffATwOkZEiaPGsJQAOSLCWZ0zdM69oOauEPOZwz0
rbKSD4CGQP6tjC2Jxw97HyZ2DxTB4KhO1Y4rl8UavGBzLN+NrV/MLfVDInuuushoAwsrSw4UW8fT
j9/BTLmK6VFSxd6J10u+BQC7Santt0ZQTzrfsy90JspGDR8L1ioF4X+jGyLnMzgndluauWJlyYiB
+DMrMXh+//73mEAbHAkkpZv1ZzWsG7pyvW/24vuORgthjv9v4SnCC1EIbdquEvTvMrXXB12rNQxX
SRWg89CsNp9WYtcY6hHfWMeX04yBA83hT55AE9l+91n5TW9UlF59T53+nCQNYHYBVQH1bKRrzRQ4
FVL8eRRapC47p49XsBsXq972PzPN3A6CztWwt8XbacPMwaEE33g7goHWK3Ijf0gYnC47+0XYnIhn
dFK5lDjrJmmgeDUrChpJkP6/uYcgLduYmT3JdZPmubcQgnSy5kmtuRfAiiiIQvNbF83FbqcjsmRJ
nVxGg8RibdeoDGpSgmdGwpsj1E9/bvubwxztlL1Jg2S4BJgH0DLvxTb/9v6/j1lCfjtAvacByFVz
LeNvtzY1ooJOM8YbjJoXPoVBz50BNhRtNraam1oRaXsstgNqt5yGwFyKL4mDtXwpp5yYUcBZ4RhK
+pTkOCwKqAV+9Pst/jJhBWi3VfwaagXBTA7oB+FVEiadiT8GVNf1l5E+7YevWCXoPCVEd/d8tjE1
7WLkTNdhSErVeHDPMZNhD/XQKBn9NnxmrZENBeEcu6Hx8YldWtSKsD0WpGh+vmfUjQQu6lCYFHX0
RdndpIz5RT7o9IkYHn2vljKesdMWQp/1Sd9TD30dsQg1BGd58WRwbdTbc5pvo4+NoxAb7VqTXbe2
g0N00WrGDmseQYrKseB0DhJyUC5W613b37VqoaG1JNTGvlHCPVXjMifK7D0Cj4a/3MvVNyNl9Exe
3hws+4ln3StnyOHBxJbZWg2Zx06bco2XgrWmko4dsy0M+gx2e13np+WuuMm8a4HWIWGfSF+8spy9
xTOsCCHX4jp5M1sK7fAL1wlYn4jLj54m/8HK7l9+psF+EuaE/dtix3ZK0MlhQJGxG8fEfNHoxpbw
tLyM+9ECfu2FwB3Qb5QzBtaXOIZa2df6+jl0oTf2KTlm9hlPrkpwWtaKneHCZOMYSHtemcWYzD5U
NpIrx1R+bGymENO6ClNIVfqehA3941jTlMYGKZLPPucYR55Pw19Naam2lPcPT1+/dpDUqy13KmWh
WnObxCDsfOBt3D97OzRswsyVf3TRQnOmanFe2C3lMIjrBVi2xvecTKVM4ouVgkLNE+QddoCC0Qhi
bxWBKEdn98eUL3XM04i+vUW2KO4lENNG37szq+5v6lN2BKTJgNyaHZotmKzMeoEuTvYK4Q/jZTHW
bg096fuWQOXjfo4310kyyv5dU02z/a2vrRkvV3F5xIIZVS6DSSpPFgNTSzkU71sDcpvsK8FV0dgI
RsHZ4RAToVR4TvG89vLEokXW4Q+irtjq4utpF4B0XFVEvlotSLjfNlPBywwEYZeUIiDWSTHrUtD3
dMc1I30lzJ7IisXXSay6Ttw5yHRAkbKlHORUkxh8XHZW0dbwx53FSwAQUTQcW5yW6kXUu109XDYe
prxanFnX5uLZaHLYxeIu3Aa4lt0ELSdIdKcEV2M2MyBJAC1Sy0HAxfMIubqqUe26YLCgLBC79Klr
+eDcUJ3qHAVcEK/N9ijaiR9qT37Yu7jcrzt1YSoqy+PRyb8fAm3SaF2KW8gBpsXwUw4QY+9TsBlj
a/pHMP8jOmi5RYrINqICMNG7oHlptL+px2TWd7IhHGwaU2noE/j7HmoB9MF0LWAFww7rcR/sp94M
smKRSqB88/zGwwG9n8jCIh2HW3W4b0fYe7eKJxzxfCq0bDs1exnG9bncWhZdYlvoKc1K4k7afL6C
rqLUl6SmIeQwX07G2ImE6qNt+gXcfdAcbxaC4+2AUaSvYqdRGgDQa7VM6ld0S1KVREGIS9MrmTlT
ity939+Jlt4VBOm0/NIJElnJ7a5bPzWO6MGmRIlPPtzk16wZeqjRM3L+p5eBuG7tHNgnfzLIej9c
jqqgsxLxHJ5/2C3eXA0wl9KyHdosZJcOviBZWDS9F/RAf1bt3WifNPqKbuhmiwUoiUSlvHoNB1al
zDQFaylwm5PZzqC7MjpCWdl/5wz0+meQUpAWXm+RAG5S5Ijd6eR1csPUP1LAW15LA+UMxxvCWYKV
r2gl1wXwzP8DJel4wVZB5+SBQyfnZxStO+DxcubGN2FjbJ1Fy7/ak5gOw7hImD48Shq8uXOey+cz
1xc9sZ4v1ALb32+D10Ammz+lGrfBcaPgSQ721zIL/D0HdPVixjMI87VRr+A4FZDg8s2zMNEe0U8I
wi4GsBlYRQY/zFjhAv6m7s2TOcctiKSzyP3WoOSV61cID+Vg2UN0aSIkdQwIfrKTF8uCq2mq1wjq
t72kgkdTXFGNBTivgnoO+9NV4TtY5+YqXMAf1p1hZdNfhEXrBy9hmLkbSGv40z6knNr9XNES7trx
qH3cM5zTA8ZsmU3g839pocsRspLmqsyy2bJ3dj1c81HdCNkVoHQ/LZJ7Zil/DTue8rwN51p74qyS
CcojoC2ejigoi4RZQA5/RUP8JsigvRsOJAusTblgX2ldAw0jZXS6bfBysB7f8GxWywViuyW8NLqf
FqvGkRpjUZfXhZxl4pKJsX99Zwf1lMEAwC5WkHML9t/5ZXMEMX7B8FoPbYl4T4GC95DNI6LzL8Sb
fxxhog4as28oaL0TTNWRfnDSZk0tUBCiAk+l8FqvwfFOIE6X/poi58bKgAUJLm5E3HUtgxY5r3yB
mEoBnyz0TxiLtSx5o1tP6nhwFcI7C+DFs3FHIUDJ+ET9f+NhTg/Kk0jDamdxY09yDHQu9zJ2sizR
T9d69vnhkZ9iOrl5kr57j/BAj+I5tZaIRSp+cg8i9HFH2gzC6U1fAFRgak9hjWau5uqrGbXFo2/x
Oc81nTGfO3H7qJxMA25OcREi3HYQKn6iIZT8xYRRaGH5IVD0b4Qz6T05i3hQgWcLSFmLUj7oHO6Z
ERXV7MhECKuQGkRUve3Te1E7JlWPTwLesa43QhXSdcVaD3hvYHXS2yb74Vfblg2FdQZz8E6nIGQP
mRK5UMSm/OvwlTPG4d88hQbTb9YWE6EmSR5vda+mmNVRwYZm3xKmPA7wZVOJG3MP0qkKTeA6iuH+
7+7MEfPoEnLYkS/aKZ8UMoDym9U/atgbzTbV6yb+dWpaWlqYqJQOPmhqZCtceu1Y7ZF876oH4PJ3
KqdvN8QxPrCGcXlVHQrUIVRth+qo5O7bg59a68UrRIucLOuMa2u1QEhEZmtdoJEknVZMaagI677F
0XY2FeRYEcVXi6cm53/aHCOkb0lZCALGA1PB//547EDW4WITztb8reBnSBUqY8MqLCYMG6rpSqAq
cCfAivZC5KyctoRNVqUpq/BTsK1NDJnNtI/23Xl0UiDEv2bgTfoSEUhDJdX0Lqvc8JYtZgOwbG/N
BRncwoTPFTP6blLJtdsCdkgWIW1cgXQHFpN3q1qJb9st/rMpzPrFTQLe2d8iOCpD1ZCwojTsPYrd
MNN3KWKfF8UAXinggeHDfEMouSjG0W53w5VE0SY56+9lbgat3Um6zsH8WLB86LlFuvlziDnDoET5
hcgQRu8ZorShLiSKNcZLv/fFN01Yvi0qD8JJwu1F6X1GP9f4IEXzf/O+bfunSAm3zLrfx3ExfpVL
tEzrhR+YnnS7frodJNbSwEM1UndcqTNrChoyGHk0fxCUJiP6B1X1SS49FqjWssPp34cMwWk0gRCt
KrS5UQscDOmG76ipMQc8yHVLUvdWfGPeQCBc00Zy0amSb8mdnnfAw9P5LH8iT38tJxHNfu59XMgb
bHFVLNnGBUepGrrnpKuGTfPUjHphpvFDFKVgST7RVKzPzQ1UHXPBQb4sSRLGiJJkmepFCq5g0lKj
BIIEHlQs9GRQzXzM/W8KRUUFMKod8mxSRpkVc9gw1clQSYqiw88AtLFgDmMu2q5/mYpK0mzl8cod
PWPf8uM/uWrB3CEySh/g1W+DHAuDMtX05hlrLiSaUINfdEp5OcNLX/tYvqPHCkRPONMFY4gfac5W
hJvI0DuEd23qwPBhk8uE/8tjZYvpXpzWQlLOatOA8IIa+V4DXIVN7TCAXrM4ysFLoUOPOWiqT2wv
nX20pyfbOCOKuUgWy49Ggdu1V3D7oo+gWfbDWmJljQDxgLuGyhctzO2kksO9Y/Ty4jiiN+yWqOVG
O5peyi70g/vJ5wA8rlQxljC3mbBxHWHb/EKcwjhwLrGgbVt+M8MoyZomaLbXhH0VVOuzZOd8uSl+
X8zzMxNZv3oKJnAJ9EMsN+37A5oVL17yfQ8UiicyW6aKydX+BY0l8HC+j2s0AJ5QdanzaCrRhPkU
OX95lFaAmb6URdrfZCDL5Jpyaq1IKshtrqAkiEJn8CQ59+u3DNMvtkZeDTCuWSJOAkzIsCSvXdpy
7NkBRKpPTA8CAKN6wmTL1FlxZPGIg2dhp9Ov5ANAi3nTMEeppWgozqo0d6uz1N3GLfrrcYmCngec
akJZb3f5g//ScWRwuHdxbi0yniT0qqnPuqkswvNeay5zUHNm9iQbtxm76JPA9Il175PlrCBJUpTv
8UeeTVTjRGHt4KYQDXe5OukbqgUIBwvQbKUPj+iBCUg267U+R3FqQgJEoZzCR2PMsK8/oBruxQLR
aikje7n6vCc6g+OQw2Kl9oA1ptr7QqXpPPzKAE4iCxlpBNcZqP2Ye0yzuCEs/a06JIojEmbGBwah
CFnSYBkx4zVc0WeXhH+UINANWZUXEA0f4T2gPDKmZ2hWvUpfvinDrp2ucCqfO3VYWQWW5elB71gg
mlXh8DGkypr0JsHgxd+MsnMIK1K8ZlP+L6JOjR93X04kTUGbfOrYmVGhX4+LI93kkHp+9Y8tU8/f
7CCMomUq0K+bgyttHe94Qo9dQZNwa0LR3QSdiIpK9IaOfJWd7huxVa6+PHWRvt4ZOzuBJyH1PLbN
aw0XpgdDXZ8OCV58xlCHa3s4uxi5PwXFi3VgJrO1BvcrrmNM1QZPIphSSnWp+O+1hzImJaKSS0Mx
pWeYGnOtIu0lcA9Cini/pr4/u9UHEC3apYbwDBMLyXkslaQPZE9GIhvIqvaaTJRfCHcpfTdbb3hC
biDN40f9gTkDhaGAkuLUEi6oS/UK4T/Rp+a7huWOHpMAyuWf/C2ptvcI1DHAP6KbcG+szWDl5GRv
ovDsnxBRl+sSuYsTS1djkwJRrRqaOy2XiecNzdjzulk+9WIrheghJLuf31j1eQ37fvT1+SHKW0zK
9qTbbte/4qhBInFa0/I5t/D/kcX9Yd6xGZ4lLX3I3C6lK2kzCysOsAMeZWB5C4jEu5jjRiHUFgCa
goIOpJBbHPST8mtLXCI0oodAg9S6SaJrKsrNHs0b2LVGw+C6KT7orCCW74tnLxJ2ADKLGW0Ows0T
MhpvXVjEnH6HyWB0HwvAiEc71v04fgNqlenhEE50PmUknJ3CHFu7pZPTO6eE4l5Ed9PKIuuJqXKa
/2CoIoNf39WuL0pAL+pkA56O9Kl+m0W5cJCNCuAx+U0PLqSsGCodDyUtHk8KkRJmOHcRtJ+J8q5V
4TwPeoCizp3od1EsDj09M3eUW+T8g9fcN1t6g5jTuHjwMk68jUsmUGO5FpZY3smwkgRM2HIBOUFl
nf/ZoUTwNAALvd9W2bTLf5Az2ERVH59tnXtfh1qNzWi747KejHuMXtdmnj58KGKsn7qMP9PK5tV6
1TIeTSa37dQ7vT/pA9lQBk8unIDZMfEia4X0PMbNejkS3E07BvG6yv+kiKbqYckdG5qKfhONvHxa
tDpayIFNsaJ9JFzbR1ii43DgIrWJI1yOqHR6lZM6GUzlNuMSz1kIFBo9IpG17R2tuj6cK2y7DlJK
GDvKMtqtfVA+4ffXKlFVLv/u2DIyT7OWWWoMFqkOG+o8nmNDdqalSwnxuXwKjhmOzy4uhmE8iAVq
MW+CD7pawIQhOIRqAYeaauRxpfDU7DopspKnKM0099MeCn9n6hFQaoCwXsj0xmiuSBdRVI2b+JhH
aoDJ11Rxeh3vxT0756loHK8v+BBDBrLGcDkyG+RLtWpl0+Yo9iZS7fAaxIvl5VMkmeNChHiFWSRW
J5AyLsKJF03ZhSBaxU4z0y5EFVs+o4lWsylhFJOiIAxKDfXQrqFnM7gxDwZBD8+GD9WPA2Ies9mc
qKVeZnAiMoqrkpm3OFxwNCFspbCUbE5UK/ozGbtadjZmd3DpkKVMsx6PbG+BOqrvpDY0QDXGVwaP
lEF2xIPFf9w8rgwuTX4AsR88pNnrjWilUJgWwWs8+TxiMyB5KrzxbES7xMtRRp8Zq+FKy/2hc1pb
2OTSGzA73z/+1PITeD+V0zioI6vwPQiTf9hoVnu66cxHlw5jKX17lqAlUE9s3xEJc2tuBzJPE+LI
vHvUcbJ1UzYKE0XgPJ9yAWCzLEEGzCz6pTLXa/1+7FqrwwCOL0TNxAZ5x1ZPK7W+oT2mMNjhndSt
cn2Ji4vEgtKHbj3EgQXWOeC5cFD6iuG7W63ZMKpLH5OGBnbe2w/DnVn1tqQUuzQMgzU9WEcuUXjg
UD1dQ8isesERczeOyqU8sJuErZH0NzVQf0w294hus41/Gw2y+fMtVWAtHfoNGGM5m0S2k4gnsUT4
MmSPn2+DYOjPJ4oQGp7Y/2yoaqMiogdFf6aibU1XUlSOzE34W1WfgQLtaSZrL8S8nw2iQ7rfOEwj
wbQjN9xAcJawKal5yOKRYFA04a22hs08tKwwMXL+fq2MjO6fGNWt30SmmLhQUhG7ml8iJcme+835
nlHUMuMvxcO94XZu5bO4kXGYEEfC7WMc61o9Cl9NY3kx8U9POcq2qJ1V+G4OsWJ+md+mWkua3962
W7RnxJMCHI45M3F/kGWGyxVf6kPZuNjI+nLsHNe0b2XnOEgDfuC3LGbcFbyTYMluh3313MeY4UIH
XC48uEjxmQz60iS2UBHANHgA2R0tx0Fqu8lVb61SwZOLVFuNRCokH/tIzldnAPK6hJSPLfaumV8L
ojWUecfQivJW7pv2x00pWq6Szv03B9oDr75beU1NDzfAj7wsk2EiWeH6C8cZKEqIO6wnAiUyWUY4
/7lCuftHxSapzqgfmL14i2nvrlv9Cshed3S51BqtjpNOCJms8cj2RAgdnWEERkXUVndUvm/Rc0dd
P3YpnizTgO7707ik2ifGXzYlEkFaf1vmuXn7Ef5Xq+Hw2+BuOEOl9xOwDYgG+OUgslKrY55fnw0n
S+Eqdkuvy/UXr0XIZbqIWerEM3f7xMHKLAiXKFF2QvleWnaEpq1AWw4YIBjE5D6NwzosoiUYQAWQ
4DQU3nDRVDCpW3rpEWmz2Taaxo8g/6q7d1es5Vy/pNL8+CsXP8l3/sfUYm7jFwYNfzugeQnl3PVA
vic+qXnrcpaXBsBqGwx8VjmjbLEVCoKVyEye4xdxLGg5RGAGF7c+bbzzYG5zkZFNmHfag3IZ2R6o
FEUcvKandO7x/tERgY/kaQSklt7p5gsSqo8SWG6Rx5Acu2tiKtjp5MyawVDqdzK6VOwC46YY4EDR
eOCpAP9z6sJ6zyfQgPDWVFzvKeyEzPWkzPdG6/P3mDSbMHbT+UrNmwannIQoynxe9R/IAwZ1lYqt
tWKoti8XV+psFtdNF20xiz/ACzSTruoW58AkYneR9UXciCAdtWgS4ecoK74OwzdF3RBVHfiMfQzW
F37QQALP6bNwyHGEXLwJY0La5qjIosD6WBu5Ue3yHArvK/WemoSmzaLMJLO1iry4VJkWrRS71uDs
mVCnLJ5mJCWH5ZZc4zk7LAikEy/OVbAT1EfsZDVwkYM60ox2w4FBTdeBknZ4w1FjE/sZPxliQCT/
aCDDtuD131Zqn/5MabsQ3YyQoimSzhzOiwIO6cb4r3yDBjLiJ3YoCgRGBWUa3IwnaRJZw2jCD7np
JkeXWqsisAf+2+gRKYYPeXKzeEcGfa0sbMlRBRLKPa7ipjfgFtuVnygzENGSMCC90JUHoo4wfH5h
SvAHSSI6clpcAP8Gw4leLwckVX2ERJo4BOjpKwcEuyNiee9m11dIVsO6MQBuoMXspY1tbNcE2cMU
e18zZMk1/kgpP7uthL8EDk9oxD9n5uqvT7SIYkAF6d+hY6MzOt5gR4KoLbAkKQFldLlzbWn84O28
eAvR/tC05bJRgatvSlCMnKX+7DkaY8Arx15ExSEPs9Oeo/2MbbcPtRZ4nvEvVfVKnQBml0jan/YR
W3YIe68Ly6Z23AIaklGCkcGv2Rn4Wyxh75pPv3weta6AzhWaPVNo41Dx65Lz3LIyW6/y8UIsHMQo
t/HNQR+TsxhbEcX0hnPkh6PqfvIkT6VsH84hPK76PHznGmmw7SbWhd9y/li5N4clZ3xsxrQ8vb0U
ktslWEQgz84dtvPnbGGYssBHot3h5Kxqa91ScPZu78bDCBs/8oZcTzr5yAxIDMGzSPeSTyx9pJWm
2X/zSrPtAnTUk9K0PqBM4Fh6PhdEL1UYblKALH6Hi+t5H1TAOHswsHvrs2RAsOqET5pmlL9mfq8N
tbYIurJCG+XUtKSAnaXlli7hPGVYftWrWZtU785eQleGZZJjB+kqxy1oDSO6f4PpurikAQN+1fHl
5RZmvEhFQwr70qmTGPMW/KYBtLLbEV535MrjYQupbAYvHv28dZ7KXPilXMwAmwZo0zCOzhpLm6v+
KZfs0in9C//0F3g/uDCsij/nzv6CftJB8vF7iRokCIHGIVVFPgAV1vfVTCVKtrX4GjEDDoCbg0Rd
PRFyEk6u0QHJTDp4ZnOGSL90RJwdZWJkX7W9cyMIclkVZ7xKPrwBQjjaAFkGQXHn+Y7poiDgJ0tX
5oZEcQ8aCB/fadF+DUKr8mXg0sqg/tdtk4Eh3jycjFI3IsEQTaSpAIyBVW8RcF6LIvRcGsgMfbPi
2HBuIvrzGAfcavxnU7FaO0i7bwImv06PVgGsdON1mfZ+Ef85kfHGxefdpjRXKAdDEReBcRtu8SZ7
Wy8I7cqjYgqgyNLy1hxuc9httI3zo4jrRjg8m9YrTYLnobrhi/+o+eH8OZqunRh0urmIhmigi+CV
U6vek18aGuyuEakWz7tey4spyO9PieOC4Poo3lTMduAqYMccMACjrOdeugNTdRi5RP2M5E4oRaHF
a2IkGqHXLVG+eEjyO7YUW5m739mNqTEf3D0wXKHqr3F4OGP1SIY3+eYn/m4Q+mxauUmNkixgKI6L
sIneLkQwI43zY1NJJ88J9/g//Zjl+llBuJw8D/VMTkpBOeylcGfBeWczkbeFWVd5irO8s2XFo9LY
2N7XUvWYSzLT9V8N6Tz72ibjewDu9A9dvOURtXlH7edJPjfk8G44e23H740WLU8ogMUatKsgYqUX
709lOYn7m86mQklC5TfrKZft3FRYZ8YGbpI6L+hIdbO8Xfyre77GLu7Ix6/bFndfAjxkBVLalL7d
IPHa9KX7ScvqlPHgy6yq/tUiMDq8Lf9uMg2j2jPI+ab4YjCCggtM3gSdC5iU8kNjzNVo/cUNPVL3
ydQY3WJqn21Yq5fc5JmbwwlfhA77cwt3O5VO/faQK+uBuZYYxeaXICXTQd9y3VxbldKpqcwqRkDF
2/+UM59PPnRsim9RTJAtzOt4oTMNgO/8G8XzYQnll4yZ+lal5uNjscmvXesc2E38iZn2+sdgkgvw
YsK/QwmxDv1O5/pFDl4zuRugGYf1PjsAavANdLWIQOqDSsiKz8QSYViBb6yaUoM1/449TDLWZRYB
pJMtMUEOeWRzCAMlQDD4NQfAq1sQIXkprhgDxM9w+dtcwEdAlWbcXnJVKIVS/WoSA6WVTkTIccQk
wrARsg8QQhseHja1ivfHr8i0uHttYxvw+DdcZnMnG79FG6ZauOz14U6mXH44/ZgDRZYJMX0r/NfX
wqJ2B2P771knvUjXW9JFAkUJchDouSXsn3vTs05f3J37Ir/aVMrb7MZnfMsiXXppY0KqBcv2SXOC
16cEShYpGQWHHEUXeZULtgJAkBIPTSQTFFGZXE6iouKyrhXg9DAq3regsE6uLUoxfr8IT//exCN6
syqHU3OkOB6xuxsUeAJERBVcW1cKEs9Q8ajPxy0npto6PGiAj1jlkli9IWZM7PsqOBPmENPli8g6
EujJ/Gqscg6lF8q3dqIqoa8cWhFDppWFIf1kAwh4kcX/ZuOEcTsJFdYppaXSJtgYas+IoqWLNIpT
xZHWt8ZWtyTGV+0VWtb6fyhA89wU9g4tW78hhTkiCxgLX4w4exZmuecQVf3E/oa8vqqUw1Nz9EuV
6jwepWjqP01DmvKc0F3Of4cSm6bmrbkDl9RWutyltaiY+kfmLH0XbbQF0oWYzw0Hv+QoqfQ2hTml
CleLzl2qEzVHtL9SmjxhMNwRdT75lavVcuI3NDpX3NMn0kksDZgzIX7T4yITX9q02nHFdVJMOOva
z+Bf6YnB3+Uu0HxcSEPI1+dQSVx3JmLR4iGTwbTxFaFmXhsVEwoSG9kxcMELFgPJfm8GaCiBk72B
KAoumUnZ+nGeoJiLeuwId02NytPlJAGTN0fd8T77QWtENpqRjapGqstWzsyIzs+DXUeozW9vps7c
vViEC9Io8dxew8MvbFvHYr5aWcG6lizseisvDy7vbT6llBDq4XQpsXktC2Vp82QrdR7Uf8QruTmd
irn3+3/dy/6mCqew0jO/XVsoTxbX/XmoD5yQtEVqqHZ7Knmddqk1weQWONWBC9fDN6Lj1bPhQdyi
cFN46AXLxXsPFbDi+qS2ja931ilSgCsCnppnf9cmwKOx7LyVBbD1718OPrzVM/dpDhCPf3wuRbcA
UHNVzpKV5KSfxlCkyYMMF1VAnV8UKYuI8E0W5/dADBoKZVXyTD7qaKJ+f5PiPvYI/BuYskRLYb/H
W3+m/cycmzDJW7ME5PKfhqWwU8BE+AAHYjWchw0x+WU0t9+4xCcH7RWExf5R7q57cD5T646Kq6vf
vItrsko0eJQyjK0hmNf+j2JvC87Zc82zdJN71wyMPQcTU0q+brFhGilGZvXcfBti/dI2W2ehTZzR
1lhH29PiLDoUa/opp03oIn4ZLpa6zjVw9eBb5Sbm2RdyBmJb13uNTgicphXRNXkGYojeA8TiB+Md
9HZy6wprk+7w2niiSiBau0k2jZot+/esyPm+YK3H/nARJ30v/V4EqkGD6zr/qwHpDv/Ab+ctXs4h
6qVHAlSiKnsHzH5HWys1tH7Red4KK4uNPNu6eQxrmrTDCJhGZgihfE3+XKdNj9IsmjycU/tWjqAG
qFFu929aDLLnRON0a7bwR+LOBg5A0aH/lwABLQU5T75LS2Jvye2yGCPg4AsIFQhF/tthmhJCcB4B
h2WhCrATp5zb2qPHCAx+km8D/Lai0x7+3OZZCcdp2CjsncX74YNNJCGMHBIYa7aKWJg56CVLaDHG
bsak+IlXbkyYKKU97BwSlekCLtTdwVTdjUphv/+8GAtrHM3a4n2ibGO9deMJD1Py8tnRTNKuSuKX
DrVa2LufWaJKVGpds3ABr1iDhH0g5RDLOXHXuMAfbo1MkKgfcDfSlkguokFqQmP5iPwScJTrE1Rn
gYFNEmP36yRLOReDJLA7jTTNk9Q8NWgMhsS7BTXdXnNhjhrxOLZtsjMp8Dh5Jzce597bC1mVBccF
DTS0WnNpl3nXK52/l0Ea4+ET81NZrCfGLOh9WpvJNEc49nuujzR/D7BpEIzqO5O0TkcT0LPgAj3O
jKwkVqJl9Xh2eM/dzMIdUsLNIG9VXOd2unbSv7eYwqXf1BnFa15+/7VvFyU3/R1zHnqJeBq23cWg
FmjpXFaP47asBTAONxY9HfIpW54K90RDrbhMicv6I6Z+cIpNzNRFWrUZRN2GxQuuDzG9dXNqtwoN
70J1DTY6KGwmlwFI1dU154SokDM5RkodPf1tVEfvLRMq6AVeREwgpegCISUTsOcVpAIDx0xiTLui
stH76NQsETOrxeKEPdM0vGNWJ7N6ai6b/Vzr3hkvzUcHbCPc4YQJPLPkpbyrbkD5qVSXtCHDzmOQ
/J+eNS5204KF695ni3UAEV8wTxKUa7ZKx1iWI+AkwFzTGYKkWt77Pj4doNk0x42GbyX0enwTBrYn
Uh9jf9Y9h9bs0lwkzHhx5BPDd5AzHkXh7l6mr7j5bBl+IzeGJOXsCt3EfIXZ7Iuz64i1Qwb94lRI
XMwOGqeQ9d87eMBVpKyLvZdkCSWSqAveMjuXfeADMI5oI0m6xLi1+j8WhqMR2Z5iuazKLVyeUThW
w2KWSmPiGz0gvmAtH745Hs6UFcqtyPocFWlonJQBTWNqlmebJiNe/VnHnktNgk5GHHeH4nSIb3yt
BFO4ZKh+6Z/mwRltC0ajRhsD4DosMx3w3UQ7LbZEmvOJdsHsGoaIOtff21+aMDRW64FG3/A0STUP
7Bu4yGmp0XBLBbgJnCPnypK4wLvCtPfQWiGVhUBAXD+6GnneJh8MfKG2wRo8rNmz5A57g8pHXgae
3FqcBZK8N3t3ZmDKpzsyAOl+lZiCR43xrOImiH2XrMYtRKwfTZXDPT0aFXrYm6TC/M5B+ffE8Ke4
9uuPFsAqAEOWouaCBrPA6HrTAiomyve7uXfTVn2q5NUDzDQCwcF4Xrn92DnBq7bE5CB5WLCr0aCk
8MKvQ31PT2MIxlPynANP+75WG9iNP7TKYnJb8+McPiCb9kLCEhu3Ma5FszrnXGrjY2VIitqm/zx/
6LfnFQof8QbpCOArD0uXcyyNqmWq/RVz79jazyaTvOmhY7UWWWW8kOBi2OvuS7buMCl4yUUGDhei
ARlEQmI+fND5sUQ83RSXDtss0m0NZgQniGmedmZ/AP5TyfDM5NE4MwEb92mq/qE2OYRTd0gXw7DI
fhh5IvVOLIOK5LtL/8xkwCa16LG8LNlPQs3UUxAi8vbASOYjU2i/WRCjMKFCzQJMv18g67EoxrxY
O/pBlisxD7VxwhFf3JuCiWm07ujZglOCBgqb2VxxX7rInTRMlEIxi8N7Qt+8/DHzeb9561+mtqGM
SNgMPAcuHhwBEToQ63lvUdbKdnbqaOqMABE8IVxShkj4gyGwfxG+GbPeKtu1bVp81tEuxRqkgakG
PaAlbrFvnnrBwS3w1aEBvucRG4KhfmYZGSsoIsj1/fla2AkpDLLjW7YpBMI4V74dWc45+YTXLcGV
bDCNWeb+o/9gYa3HTGH5eoI4mTBuS4oHvFnl4kUmqDGfOxBvFhDy2iHyta3aeVy/bKf4X8wLZwJf
zp/g/Z17R3IntUV66ENxGvZKM8CqOlP3nNkYneDjka1JIIshPGBRvprjhydoAnAdR7ArLALhKjsm
UxVDaphYR+8LQxS8Jmp7M5rUHnfWXSCX64zM1Id9NmAiNG3Dkep3Wgo8Y3mXqVjbtuSRLdu7fKv3
+0TclImRggtNMPkA94jI1WRM2b9SjU0EYR34jutPK/FIjmZCeOyPQHFueSNfg9nlnq+nV18ql2JZ
j2F8d55+Q5mUXdd5gwRzT0p0o+v1JMcdWBA+hxS+lRunIMugrMFUDiT77wl1mSd3hZyNaO7quRmj
UbEH7ac9cGBXT3LoWZqRgH4cGbYDG76SGyS9RtzAKTqzN+Iv54vZdCnWV3JC6vVnACs+jdfo0DNg
MO5VUzJu1AT/417MpFGe9Y4UK3c6ICsDgQdwj6pBma0wSqic+uPbWRdguLVrGw3VnHfmJl8WTl7G
A/RRDRi3/Kf3SiTWTfKZgaKqk2Uemo3MOWwOSGAgtUXpRTsBx6TH42FB/zX97HkS6totB7R5I21m
XEhgpF5RXEzfG8TESV7G9PHUwflJUG6Fv6ds+3PNXHsBPlzQCVzn9onioODWTVOzFwWKEb83NlPG
w4GaAAQYg9N08Jk/tzs9GuJrNYHglODupOZEfxs4AQhn1advcfKS2sluunTmcj1lxXyYdlQl2ISu
E93/dcIYnBENjxsZ7pLn5tQWbs/rROHC3tdvps37Tb3fqO/lSoPZuH1sWJ496nlrIpexeIUQ2mBJ
BXm08l/vzgraCR7DnDvKmp3hwCLyXxcpf53hdoJ/1dWlsXhL8p5oc5QrCw5K+MKf/K9FRO/jTWM9
PWmlFRMEyqOGSlFSjiKXHH7qB3p/D0iAF/VhE8+bBnWi4PvxarCKb79jiBLMaRbCKpOEAZXc1kjM
66awEg1aShyjyQib0KlMdxJpMKudpnLsp/AV5zfFoQ+ANZ7LQfo2Ve36409kuHyJrR3kXUxIU8/k
hWVTU8plcaKv1kdaS8hinpPOkqqjotZojE/mkfq6ddHIk676wATDaZeeIoY6edU0symFqbBaSRWp
GPtUHBUJoNTJlINN/Reqp5fT+3tEQ/KcA7Z4oUrdTdKemchDzo24F8Vylpro0wtkvFd7c5f9/1xc
LbnbGT8zFVeN6vsGIcUXjz91kgq6iiZmkJArCuUCMVE3XLW+pxBFg1uElNOTkdhKIXEBSDliKFdC
tw3ydS4grgJHaE+CwHe0Dg2ceJWU439CHhCO+dc35QCVdhew0tYPLYG+TIr1s+D7CHUiyy7ZQ50i
1YhgxM3e4HNIgqD+XVa9Eui7ELEWcNkHhR10iIiC0ta0JZVDMjpwDCgpLbaJHCl1gBziD+Rjmt+Q
zPHgqXSR736QNPrUz1snUQW1LxnD0GrA8iMYl1+ZnpdLEXk92oStCNG5IVLAt7UbeC5Da/MdUKFY
EcniwbyZfuzaBHWmtb/NwzCYfqyQCgJ8htpKI+xt1nIVh+FIjm9ILdvbjYOyhX7K26blAUAMVQGA
a+KGcOFv569K86qRDxmH5J/VAnhcZXLlCl4Y1J8S+ir3rFif1K58thRwHqWmqqskjijNuPQCrOjl
rWDBmwfkiaPKcU9spi/AWoCvIqSmRu1ZBCLkrPMzfcz1W17I9DNuzEFF6AK/VGFQhA+xT6uL0Ate
KxWVZswFyq/4M+I/DrjBT4DNssrpOF95RlQd46O8HastcfDi1rtmxFvp/cvpng6RsEjcMFGqUAno
RJBt9y6UcE41TUY67x4G+Q81H15RFZm6aowWbhKkpHRZ6b9JeS1jWFmz0e6Cj8lnAZLO1CGGGeAN
Iuf+obtGBv/DRqT88tdEm2qWtFTZNzz33RsvrLn/nTTwU87PPTHQtORmfUKJMG/5X2dM8yjWmp/N
BPyj3C3Y5CEpQm2GP3962BbgRUA2jSX7EWzr53DXc9RWkxa13ef0L5R1nY8XHmWpJ+9mecPoN2F2
ZskJbxnYzIEfeTUCXxKzjsuVrb1/JjkSU2K/+BQqCNamKWx2XuNvEh4cdVz2ypnsuaPthWxnNV2q
SECtW8kDxZh/R1X6fe8E5kC6zg5eN9R4OK9XokaMOnXzkEcwfESe0YVhH7p7tsk7iKDZNxu82Bum
wLyPKtEqL+A4ZFnWv8c5YS2TSkaXnrYr3zbu4zOogvuuFp7GPkB/R0G/fH/Yh3dRunvf+h6qukFs
yXlqMG8rn293/N8J2cke/BULsLIvqWqFN1Jfhym1d76nOWRNDp9gbVKGHQ9OvdVJIDMPZJs3/Oj1
vZOEk6aT+zuafp2HRSBMVG5nzBxNjnaHvIs2P+fNm9xGHUJC9MsQlvMpDWmHNLT8gLc/dTTs3E2g
bnia+qNzVysecM7ruJo/53myfD9gSL13t2i4aho4z/U281qUMblYYQloOzcKX9yvqqMooJu+Gxjr
CQP+ko8dazR/yVQ41d4xruKs9wbdDSX9KOdnk1qhQKjLqBeyLL42wU9AfsA3Y4CmKzUZ64ieQMAm
uMruJX7+MNIjjVU7NHBxEw/NgoqS/SOSTb0a+D4SC6KBUUF70fn68iNoojFG+dyBdRKWJA+n0hCI
d0bEYCQN9uuUZKzdh823YLPfXg2NPILM7ooXYe7/NRiW80KKxstgvVGL1YS4MWJGfEfI780n+pB/
nxXT91ktTC0rVjJyAlgDSw+GuRSooqISveuL3BgpdJZx5ObRarsxcDlJFMeL/1kNkOp61DEiMzIS
p16E0x+eBrsx47VYAmYYf/oWNcsUs4qFhKC3TtM+MzUGLKZyhlLeSHVvXoSbKSCMXWsya/0K8bn1
iHdsETGl9w6LHuGWl1cdOloymzHQaRhcwc/NMWCjoDFE40y1e7ODufPt1EdfkUvCrhfo6MCUlkYi
uh65E6+Ue8xnL3kJXYWAENbHpFRHKGCNk19oTqGbkeHxeT8IEAanCNKx32afoVgwWO8OsF9qANmJ
zkFBQ9Ya/qGYT/mhx9ccoWWrgA1yixjKj+HIbuxW6SdX6sg9rfw+/oZqO6KwQI6trq/C2gWlJ7qL
oJJMsLd6swS61xnuejg66IppNHHFZDYNP5VP4qDiOjTd99/t0Bd5h7pR6JcSFI/6EBcdN7xPgOyg
da8DPfyWeKjfumzvh97Ay43UdE5NvcoR7YofoId/9GbfGI+79QUH1UFMPcMMk00Uu5zwc0LZ283N
XeFha4XzQ99U2zrmcMVgwwZJ4SUnsoH54K98mcSQXOTgV+JfqV06UHOts5yJXidGNdtxbHsgLT1R
qt35VYqxW+7hI7kjSBrqcc6hTl43IuHVrazQbZgCR8u+KugqrSkONVogsPWq+y+4i/2eEJ1S+pIE
iBho+dpbCRqhZKVDu5y5iwWgNZcpQQ9FkYKB6SH4lkE/M4UXanom2pX0ydPGkMLnMXnmPcEhHn0P
jrPQzH561i4MC1/D8uFyU0mRjWDkuiNNC60pbexpW732UO/oBlf/ey5jWjQxaMZ/kj/jrbMt5k7C
B1MfZqJoX5fLRp8Zj5GOzsPyeOK6vJ/HDspScLoXFjHyyCPE/tl6lPo82UoVW2YWEB10elIbc51A
BRP/F4U75VYaIm9sWrZ65l5idFuOR7+Wt3vCGp/rRxqXuTBoTmg6PV+9Ee/kcFDxEgFhjQAFB5Q2
mRjX4yhA6+xe7p0x5M6xNDVdsTshpIkYFYBSxqzW0HpgDMKI+7uWw0RHyr0iRjx0niyzKc2vWuoD
G88VBGMrhnnoZElhu0we2+xTUe3seBT2kFJYfIXxUtd4W1hwOJN5hlZIh/e44mLK2ez958GPGSrI
S2qzcXaY008OOIEGBh1TcEyGVjAB38xw2lGC/mlFvm8MlmGMo0dz4TfrItqEjc3gfEoes5ZbWH9c
s5YaO1XqtmqScNZSRVbnWc7U7xCKhgctHzF0Kj3ogcbv9aJEnYkrcI1xJJBxHVVfEtKU7X0MtLHe
7ImU78JEpnG/jQayMmoJ8ZIUYTFJCZmMCo32iGu7sTVJMF9Xpv/N00kXyZ8q62SLEsmY98qnXt+b
mKHqIWsr/o/4KzYXplVjf8zhhT6wxKzfwud0qXTuvatSikaDqLPdK4o5fyN+ZnYoj0px1Yn8vGxv
lD3ROTZz3CdNIpEGVic5jKCvVj4RRobBA1mG/6yG8nmtlgPpS0lM+wGG536BJ2ktNht9/bqL0+/Q
fLFxUM0YFYTpa6FL6yt4jByo+HIvCQtEJnww50/s9Z+5EQL9ZI1OYXfXIA+aHnB5TzMIpkT5O5ZW
VFpbooml5vVfV1FIjo3TAp9Qa9VwWmh5KvqN1Gd8ss1VSSP0jzWYlE1bboxfJ+FBkjkpvsHxQGyB
SMThvy38+uXOcFPjRXxRU17/JAq+509YrHvUq7JnatPbTBFdhn7jVlK9O7MzMwB2s9rk/hgta7sG
AU83fGLuuHBDS8djwTZCh8K9ue+GG+ocLJsvdDclaqVBeo0cI/J82g/+Lnk8wvEyxwpm6/1dX2bS
lC2o9obu+f68QLEWesm8MfCt79y7h7/T6PkZHh1zPJ77P60uRd7EgP4gUZFakQN+oI+xl2boEB3O
1Kpv17lCWbdZXTmcvqxHlB6ssiXlMMhpHxrbJGh/gh8YO1pxQfoR2pCz6pxKLWKRRBgctVJZn32Q
niBYj/XptwLfHpJQeyuhvNdCQl1dQFRtCwVgnePXTDshcoIgy9sNT7yZqc73Kv/WS9JtUA7XDdMy
ZscF4WV2nEdvwH/xTZgPEKgAGZ6EIbThwQ7dsC2osYv3ediEMuiMPbUh4AX1SopQvNm9PdLueiMr
SkUqIC7H57qVS7pd9FvyBisMonMvw4Nmdc+V+b1yWIwxxfXjKMh6uSd3CS6P9sZu2ZvR1wZCrtej
AXeYRl9PutnNMmDqzB/kvfsx9UzjHOHLMyPVljN5RW5sbFiP918cU3Rw6VkekEvhdUiVFimvT1bx
Ee9zy/UgONlB+yqo715P4tdcD90YZIxOfTQ+V+JXZfZWNtvxNfVmuOfDI0GoUuT5fgNIp8EWXzrG
YfNAyisb+ZW6JOnj7ok15NFYw/Us98KKhsiCN02BVtmOjiKS467SLCyMINKcoIH7Pg8gMgTrRA7Q
x2Adsm5HhXRjtzg3aUJKLwGA/CLR1oIYfuyT+ZKyqMrxsRqgQYGw0fWuE1cbDnmjJvx8Q4KgN+zW
1EjY18FNGjHyxLZ0cZtO9HZ99Sdd52bkNoacfX+QW5mxXrT6pKzK5e9hTA2KQqr9Glhb/jLPa8ce
evd9t4YWlQQH2B2GCdshgRtsdb9kMX1hbjCOstZxTXsQlHjNCDJspyZWMTnga48Ih5ObfLFacQgK
KC4TUI5irNzcsR5ijlNgeW0XRld5B3gcxNAefDBayTSyK5k6x0ggjjyV0InVKeVvKGAjoNB4X7RO
DeWab7k0ANPhXDmlWDPbzZBjAxd3qW19mNY8e9TYfMNRNk72EXZim/RSU7CODP1ZBnZt2EdKyozP
dBxwGBUP9d2U8pbZeKaB5tDhGcaT9RIAvWHUujnpqARaK5sCGPb4EtCX7ICJplJgql1A3xnnmdnC
uaSVrG4imLOACUczFqrKA1ejeqFE7A3swtAEfO5WSRxhSoS5Cml88D7cCXtGlKLMysb8cxwNzDZV
xq01pDGClRM8wGPUWRaN9XY4NbpZK0/SlHA8scT88qikuTQytw5QOdLsiB1vul/gR3s2VztOclOt
VMXXpH2ftAg3zWd4zyxVNACAOFE1YVyKBjeLg0NXiXjJmUPfdpW4E7g936XSPMfAOWBL2GYG240W
j5bBgCS14WxOi7Q76HpgK28Dh1bAsSLrIVPkj15W/y3P7Fo8ACxo/9fClrYAum0aTnLTYPbmCQ02
22qWJhINVq1zRdqe4J8pjMm8gA/4h4vc2ByNLJdEjwIYe5qHQg2cjZhLtK4P7FzW4Rs3cwmAotwN
p3bUUkAAzCYOUUo9AEFjwLyob7CR2UWr0/bMpBd9UjfueDx1+mbKEIqUfWezUilRC3+WaiL74Z5k
3ACeo7bRhcCLKsk9q8LqrlSZ3cq334SGYbKAxkKVwML4JLRiVBkJOruBanvXaKDBIz70czJw7EWO
7ane/gGbcuNmLAGPaAy+gtU6AXXLZ2IIEotyMad2EccKElC+8Kl+eW92ueFk3gOB2nl8UYvhHL8q
upyBCGvw95BYGwujewI/axxC11h1hZr0v4ftj0NSr95XPtObhsWSFdzwxJlNAqZSnGATmEzdkJYW
7Q73LRbQi/odpV46VFUgrYGMY32KkCT9oLjJvhW8FI1j94JPMlilF91x7SqOO2yegvVdHNf991bX
vcAgmZ92vydn0wyhhj/rievWTZUWk/NLP6agYPZeY/VvLbYHsOjIQSgGPJHBqiY4gTpAGb+xdrFM
YZozWhI32V0aHXTbp+MIAfZroNgJ6ugYCxaUPvf0nALLORM3oAcrCzT/AQVvechyQosaDyJTLjBb
tKAAFX5/LgJvRVbrwpbhTKI6EaEsV2NnQG2TUCI+DQxzFVcHSGIGyMjvdPZOgA2pa/7hTp69+b8q
46KYhKpnoDVmteGrwetkJkf1FtERfWJ+vtEJ0CVg6RH14S4yMwbQfcXRe3yUQzu+x5dl5lgE+AuZ
ko7EKLkVJldmk5O7w0ZhGkgHaT64zMAq5PP/1pfj/p2MsuKYVkjPCYxjrNrX8iipXi8WVDyuDt0q
Kq4QmSCduuglAVSwxyKnmSy0tTe/HjYP6tjpMK5pENwOF9f1khqPT9iXoh6M/sGHzsEHYLwtFYUu
eCt3fKNZ8cO7aRTJYSTs90qza7LnbEfaZms0nXC+mtPd0q4RcJbMoX0MVXxnz1HG7UioUs9XeuBw
ES14dTNCAnhVEQOncqSmKybOK79UTQPt0PMJ2LVePaDfzLnR2LehmySy0J+6aEpJaPpo90QMzrWG
nbWfyu4MUUN+1VM7PmXwceHTWmpYBo4hwpUGS59kR46o4vcZy/I8aIzOx2/nhAljjGgLD3RspLLS
8UWMJ9Ng+ldzpAqTgCyHm7IHVowErZq6+2014o7uXjj8/cGOQTc8oTNqngS2N0KhrUREMUih+U3z
77lx4eNNief3dZWBATZbiss/RSDO499eeaiQ2bzbR61IxtAEZBdQ97orRDmNFZax7svO2G7I080E
FbWmTXrTZMMUzTXLoXP9YyraLZ9Og63ngSAIA/6wJ6avWj/0wc1+9hkPDnA+jD11JixrSJM3ZrLt
8XWxJ5Wv1AgHcmo8ELNTDiMDBWxHtrbj4z1Ovw6LDMPo2uXa6avp++IqMHs3Jb7t+XsRNZ7UcWSL
lR4vFNoNAkI4xpWiPd6AcEJayftf5E/RHKkfG8tEmvY91LYNmiepBY8S7BaxSrM2z8GTEEaqbkkO
FiJGR4TlM8ONtHZIhN5xnA7DWjZDHJId3hNOu+xj5ptUJeb3e0Yr2GK41KSlzLvETLCyovCe+PAG
jAmiWRvKhayWovM4i6nRjwUgDtnT8/VzAGp1dUuJX69DA94ROlr0GXMaxxSx/Yysbe5N73SjLCrd
UEGMtibCramS3PbzLd0jvp0PDtpZ+n8pc6esXiAfGRVKnxNKU6xWd1c+l8zjen0qSsKo4ib0Pj71
M4LJQFMJTxfi/ZfUnpek7uFlVkdvbPuwjPvE3hOiw7qpwKL6KsenErZrH2mRMxrEXtVFsHg4y1Tz
gvaUrauKkKzvLMmJQfw2f+YveOdpZI7XWQzpBB4qxweTjaOkLJvT0AJU6YSZShjIBYPUayHqkz3I
DTsxBVQBgWjz221Pzs2DSHRLZ4AHF6jSJGddJ5UZShLhvA1sWMs3wJXwb0MjGW1UCxEhmTGmSqP3
NHBonmAiWXHMdGVKxz3ciuT0z/GH4TAoByCRgFwg5t9CSxEKK2zlzE/w0rdLSNsBDB+eLlMRIEND
o2ZjHJtDqkw/oshNTB5ulr5pBGmLKZe84DzDY7GwuJz7Jk5J99SXnAC/zM15NI9VR6+EYHTdRT2y
7A+BE0st7YTICY/qr6z+cyt1fcvRcPCHGkT5wvOTe4XRhYSVCPs7XBeXcPB6TtE71AodjI2/ky8W
ge8/PTW48kYiAJIUmZkrGdq/QgkC9IKknw2t8G33QeWfzwzPD0cHzPrG9QENB7j6Rne8OGhglWdA
XUEujJEQIfqE2SUlVvPdF8MqWBJNYkshFt3cBs6ZODeQx9qn6ShEHMsO5GLhvNP1yXvGIUggafsU
COggFwb066zinTnjX/zNCjaS5xYALrm6mC4wc6uDiMRY5d2+kBSCE5mLClZxj9vI11Rge6RExWB1
gsSoxOGCZyStTMcZal5cPrj6lRG9QakqCY9SuTg3KR6+2FlXytVYxAOFlcz6wg46iW/EjEQ6pVt0
mIlBc7L9UKypYSXkrYe67n+q1sM1o7bcuhNbylfgglfiadKCPzXKHpFxf/wQFDtglg7/Ux9pNj7E
6l/ewihKVdTkx/ZCqhLLOnC5nN4cufvHFZHxmqqyoi0f57FoAdGpnal24+ap+HmepZEvWma7ZaNR
FDCFBdkImVmyqoLGu5CG/cPBWV7VFexeEQVsmfmb6LR/AAWAIIKstD5I67bakKct0/kwqHaC3XEA
aUdugRkz+yKETzmDMDEKIpNj1JGoMmJGNDWj91pagJ8/HEenrsL1/F/SWBO+5gvx/eB8lKGhzyVp
FvtM6aOffCEVuz0RYPAZ2LVQK8EMcc4zlQSoB04WKj1qWjvFq0XShC8h+TYcycbdOxqK6c5kN7ZW
NGUaeXitMAtY1yfsCFk5j01Qk7sQtyFUY8NScOrvIEN9RlyXtOF5fl2Vh7a/L/G+jv0hq3gUocni
rOkgRgN8JaeCultfmxXxCaQkWyCE+O0t9a2fcKrXLRFHMB70whLhJY2Fu/tWvjzLMCsZYBzUxYk+
Lq6iXKiuvcr+QaXhTELJLO7PJ16OSjMTHiUi6XPOBudhhaSvP//5WAnHX5fOlMMXQGPrk+kUPJ5y
FOfrSjYknPz96qQi/prVqA0QdPfHmmW0Opw/p7zky4uzpS2km9osUpUHaAn9u0iWYBBc2nTwr+t8
iO7MoFKFtHXXhBVy6cPukcshLg2QR4UwK4o+Xs2vQik1ZEbxyVI4zYYtgSo21xWYbAD/bXdb2Q1X
RJCPpvchuDpE4o0GKEMtKcV3KgGPmNjMHDbv8fEF74DR6ieqG69GLoySfpZQTYz7O/3RJcYoTK4i
g3yhcMrU3o9z0QadOyOdVhK6v5UmjKH3LDO3Gnp1NV+AjbdkYOOB1BV8rbPYYxY68wQ1tENtSSqE
AgoIikMsrT7eGEFwRCMiOd716vP1dDtpCjR+hb3cE8NgG4HFDYvoL1aA6pKOY/Ioy2I7h8vDNXn5
Eavy3jkFPby3tVjcR8ULi+BWXeSqLOv4+iWfVvcvNJzC8Ab7E3AaSdF+JKX0VIsbDhPKgYGKufPj
eJL+Lc7D3fpBjuALKGeAbdiGBbTTvSRX5IaOXnNxc96M0iAeW92KpAp7vxG0ByWNhctdBXXaZ4CT
Vt7fwbZJyMF4XkMkwUQEgX8z8yYVUbTJSaLnNfdUwugME8VFNQ4ZsZ9iYgsZlHM7pAUf8mPZdV8Q
uKycrtOoKJFD6dgV6pEFCBcl9nKUezhluh3z3K1ztS6XuG+TTqgk3x7sFFW5O6htiUpMcKw/7V0h
9iVFegyZUac1AVu/Gzxgx9Qk+l0PKBI/IGL7ZEluNfKFNYJUo6S3afJ2FupIKFw2Ele3cJhnIJY5
Lw/6zbw3sl54WPNhu3mCcb4o5aAlZb6kdTvju/So2lGvy0xsumD0HwCIYILd+8D9V0AADwMckeNU
hkIoxGdlrGrdEn0x0zyp3VUpsJcZ6eF8lMTzJ50ztKMcDW5d7tubjwEL2OGdZNYIWsXyUJS1w4LV
9Jf0rNPdsqliSSLtYq/3ChyHNh1T7F+2r2G6kXA+Mvz6x01iOAuxNZHCRVwlyDCnZY0LHn/NSB/k
2HVQUzQaq6X7Q+dJFeIgRRizk42Z/OUWKAb2VM2iybJp4+YWIB2tAhO5D+5+5WG34iK7WEtnnYZE
kmOjJ93nZWvnARFJi/PaZZCLOTa9cGaSao9BxnVCAL50jZFQsPVnAJXijTGpYET/SrkHQG0XYeW6
WcxqkXNV/JVps1yn0pjyptcQGOInCTcvTmqz78EfPC0wWa8PAr41lykhBJLCrhRn8Ie+NAXfMrwK
/yjcuC+z0cKYhwFsLLXlsMvbE5Nh3G5EtFXBrEYi69DGVF/FsM9SVUT+69Dakpjrtcaj1LDogw71
A57c2Btc1WRPjEb5ze5kpcojYCpOvg4KFVPb50eupqJ5fa9kW8kCjh4wi0JF2aFWAFbVGQL3S/ME
fV4h/eecAMg54LGQTS8WOJAf1Mh+bsAlmn6IhiOpVZqmuGjNo7JbL5eApCa3m5Jn7B/F/pDm0+iD
uKopk5aDimk1ek4T1QM8Ug2tRIBjK8+nImSNXBAPFHo4s8A1d9+m94C/Olisd8x587jTRqzol15a
vPstqIJwn5IxIGESTbvKTDiw1fcWM7MO2VKIEBiLbbD74itvTvV+oxQwcFb9o4hNKkAfmCWezceE
L1DHtE9vJQmD7rIAj5mV6o/w0Ut5LIZQtUaUyLXBXAvTzMe18rYJmrC/fR9YzxO0qkefqzeD0TWE
vKT3AFSecFLduLzntRkoxdgNxJeWqAAsPpR/wep8PL+/soqCTvf+HUXc2ypyZbmEPQOO8DhX3Gtt
syrhgbSJFgIz3UTjpIUGVk+W+/Q8/3oDZw5oUrazvu2mz7w0QI4/SmP7bFNfHmRfCSMWVNgdoykn
DvN5duHpq2Ow4i4inLAfDAiDg4eq5GWZ4en2J1nzaXduu5vhAfJqTKcCpyvdiCSxVo2qIu93AKuz
EpDvUHxgcFbe0YrNdRHVr0RxqZa8o8j8UTIpPPJnaA/WT14WQljr/eduocuedM5bOspNPdtYH2AT
vUCx3eewtYjkkPNLYzyRFW5wDcww3N0NEZEUiS63KpAL5bsTvsrd4gY62Ks+p9+RxlC2OiMBN/z8
poNePErvvJVKBLXlAAkrgSSyt04ES/CYrblUvph1J1kMWuhRhahNDFuugbCU8LCz0VkFoS4QF+o5
rp6uICOit9xYOs0Y+SNemWpR+kT8HUHkvtoRfX4pRsBOVH7GTf+iM+v54wOTbaxHD1LlOL9U4y4g
hZcAVk1VAW9BSqW9xL47r6MyCzW7iqErhAOMf5SVy/Fems5816JFCgWyrf3c+B0AuGZjZZmY/m8L
2ErbKEEDbJ+0Ii0M7G+l0Nq2496rfNVAo1z++EQOmuPQ++mBzQ9RK93oTkZ2u1DO33I5assSOtcB
+vIKXVAQ7ndjlfOI4y0BGGSuZZrj4c+JkMXHDuUe47Qb8eEVvnh6sWj4JOpMYEvuWeobidJ+muqe
GuEBRBQwn3WyqSRYcGKoVSaQI1+Zy9xKWObnT5bpEYxi990FobZOq8oEmY0BUabHutTG0VT06fVa
WUq9dOQSjDDLjbS3hAWhSq4O4yGzzn4Qt4alRotXcdug56nGUbuqsBXwJl7no+U/rNQTqZWgAwPl
xVGkxGE+GMUMLqiuMjl8xvgUHwX3+Z8KGLIYHT21Y6q7tl0SR3OVmb0wDs4/4C0/dAhpCSrjMzu1
SqLiuHRjJcRpBOpIBBtwAzJLVujkI+cgxd98ss4F/gVtUcPsdhzbVLPrHp/rTBqylph72FUNp52v
VodBeEyAjImZLnbfswuCvSuwGjyp+62JdHP9gpUdSTFO5fMJhhK4vyPKglp8d4m4usPtNaGnYEK9
mWGpgkGbUXEpH7WbFGVDJL7iqHgSbelAyoTfXAmWJVSsp9IEegdRJ3ptsW7XHUqw5eZJJ4J3WRWh
XAuVD9sZn/45b8y0j1CcZB3v0tAri7DoJzFIAraOFOs286BeMAq5CbgY7sVf1HWrSdxYHVQmdPcy
+qmk5LtGNHJKMLgfeeux3Eix7imXliI3TxJHs6EVLXTQ3J/zUvDEZLT56QcJ6inccAY32OozB8OR
jgoSFfUxJsKKk32nTQqFqCPU54c574zZwLabd4PjhAoUPd5khgCJw1ZJCzAtAZ69VTeFPKwon8ls
Eyo1bJ1lKQ7q2parzXimSuXtq1R1UGcPLfWPatIoamf+h9ykpH8+QWsdsdm6C6MrtKuE2Gx8LuBz
SRdmGhEdY2YDk6h9+U2EjkFncp/sz91qWVUJG0X8m+jrS1UfJ+XnyxpdPDAi17aukp3as1xa9617
bGXfo/luY2G3l8AB0eXZUeP07OulZ+6JibkLHzb8CQDmkrQLa4O7zfmzd08IW6dBjqudSgsLU5Hl
+4LwKu0/9HdkG+c1ZsS3UP/optErSpGoPkQ97L+YjWDqWiMTYgi3zKqkDsi5+Qs7g91lyRrAVPV+
Ixxxnb6rEO98h3OypmTPJodTeLLrhw7pdZBC08cNNxxBmKFxS1UqqEZIdCNmLc6k27eTr+DCu2/y
ECeLOFxDW7Q9JorpnJe3vHuLtDqn/HwCJ2NtSADnXQkngS12Q6YUBIDus03BRr30eyEc98jDcTdv
fy5evDsHt45Y12Q6/i+jQH5N+lYgAAYRXnWfGZPBG3/MjNE+QYF5NfeDtdQZf7GrrWzo3+96TCi6
LLMraUeEoQ4PxSKaxuYYeqgI+AOMhfxE9R7pLu0d9xCVeW6lGzVZXeJmdtyWl3+/QgGRNyhlrav3
w1POywH740AgA2+z2sWus6GR0Q8wrT7unDPiH2xWeVbmT/3NQ5wwC1E8AsEz0qqQRMtC/K0A9SHq
MGIyhHQtzlV2GD3NdQwGZJ1W6yIlc4RAu/A0wwWQBThKa2N159DT6jNAMD1PFJEtX5fuQiepKmkV
iJfR7Jk42Mshyf8lsC/nGZp0cX1OuvHmZXNjhY6YcyyKHz1K59CqLHrTTN6onoHDmDj6c4X4Etgx
UtVXGmafUe/FbJpLTzbUk3ehvku3uISL+9LQqJVxvKVV+U/Dnj/7U19Xwuwfrv60CUZdfRcr7tia
YO6UqBDVzSRrh5o1yYaWeHaywrGs593aczazZwGY7Bw4KKMGxRhgNu5MSPPG7C5LCnAHJFWVDdX6
ldLbgLped9Hh6Kggx00BMensAmrad4OXknB5jbZYU9/zFoAA1CBO/QAQsDt4dM55dA6wr4tffEDB
zSYfBQwLE3pDLq7S4i/b+qcXS0XM+Wznu7pTZRsCRhQpx4kyoKK4wsq0hz2Wn46dg72FTG1fsigi
lxPVHuKXvkw1MnMLS7eRc6LBFl+P2Of+bgWnOu2faLBK49fSO3+G81YRhej4LpGT6JBaqog+xa4l
ilcYXkw0aJ+EGoUCXgYD+0dELz4dLArt3LMwDVqHv3v8maLDqi711QEzHEpVQS7mYiZ7ZCkbPj8d
RL9MmEEDjyuw2fy8NvZ7MS2P008FYsVi0V/lUq0OHYoGEIa0dMNwKciQBuJgsNjpFL0sH9mib+zM
tP6//bH2OiHTsGtOrfRPJar+tIspL7SpUD2teKajO5Kyj8TesV+z6f65KE0gJ+shEOMxxo4hVt+h
++OcJG42AyxqtPwNOBsoywkk2/5c//fWmtwfuPsX2Nw1TxL6H2phDhZrmWPRQreXYcmFbZsULNV8
DYOOVbnJN0vhAP15ylIKpb+1VYclr2V5is14IwzlI8pbq7J3xHQSrIDPE8F4yYn/46/KMZE7fIpk
Jl3cZ/N2pt1XGJU/47tpHH4mGbIR7HIQL3hXl7wVpOeWLWg34FghrQQnivVa2O0xEaRx6MCEfMv7
RRaaCmdbBsW8IMKoc18PdcIA1jaEtZYU2xMuBIRHMeCc82h8ukzDe9y9QRin4/0jaQ3ALWYUAZ0w
MUNam2+/GT+dK5/Nkt4bhtFgyotvkq8UM3G+/2NSinX0WU31XbJ9Yjy+HvCMTOvLOvBX4cUrv+3Z
hZ1VCeOb2t7UDT31LiuyO67xoA9Ycru5lc8IrtktpnxbCpsfiwOCS/DOQh1VzRDkKS1OoAI6yanW
XIKAC15gZPNAelKy9Y3g959wnuPxnaL4ZHQNQP9dqVAcqr8qH3/hQQGx2cJ+6b0CSyQ8g9kcZo0W
s4u0bE+x5PXn8HKaVrZRFTBtpN2jo6bDxzzGk0tvole8/J0aa6+8csGFKmbW8yf4NlU/R3QnPqmU
+rTqZejWQJ0WVnMnf65i0q1Szzb0CDH63XjcEZ1FBUQapDa9X+u8irIph0ShH+aBUI5uoobW9Rnt
aNe6CZv7RhrQvZ2+yh73U3Pr2jkMVKD44ObH/1stOZ7ExeKbsl1suQsKV908Dcw0fCJfft1WzBeD
p30/DwtqsowkezKFw+gUcPDUiQasgYvfjoB8jXxekOFqZvJ2ytW4qIS6INDJ+tUqsbDwXjYosUky
gWXIurNJw6tkz3dEIAINfm1c82SZswwxGgxAiff3MN59wcafYn7CAuLJ92G6QQhJDWHTixpdV1iK
+8+8JDxZ5LSTBTgrBu0351WeLXBrUYk6jQs8KXtxt/fPeDN3HWJXx/nouais2oc2xg4uyzGpIHZ2
pBVRYiTFdeVP9nstMJkUh7vmeKQQk/fdTfQcMdfaIgahr33KmOaOw+K1ckInz+zoI57oghfV1NOn
0ewHnR1X9v5bD9SC43BSPrYqFqmLttmdZiTv6s5Wm81S8dRdtiERFVjaszJC3Bkw+eqx9mdsNlBt
JpSgG4ca5Bqjz0zXOwUoFRVYr0WywY+gCUYMo3k1hrttv6m0uK647MFHVg747ktzO2zCJd+y+Krj
FzxtD6byrl4KU3apDUEpGWRoNvrYycpWbO87SVMGtxDUV88bxjASaS+ahuXPSASKvuTY4Q1LKDjb
fq6IIi2ogaHkcjORjJtqMPhUMEw3tmc5Iuy5CuPCCFSwptpIjajLRyksZFOpOIGgDsqZXfQiaclV
vdY2j5O4pvhW12jMlgnzH+kpaDCvSKgkIgObrqdyCiL4L9slhDyhruF6JmBWBpCmEXKkXDDTW9mp
bmmCtnFQvFP3lvCqMe7Hk0RAhFKPXO7xCIYe2grUCVN0OyW/HZR5seJqQ3p72n6V5z7iqejNoi0i
u57fIxijqe4ABFyaxcrCvL/UCtfv+Zb5pqoUcbBDVi7wN5gxgWih9srWUkGdcCm+qfOwwHnm4ii8
mM9zXR5LIqZlTqR0qxbzNx5eU5hdf0Ppy3mGKhhwZN8HkM4Yt69gO2wzQbf5PdiqPQB8m1H1KB3W
XVlLWkY9vQqyVH3BcXY4lizCgvNU02NrBQkJ1gaSzhWhgyyrwZh6bUROxOR/nSEZjJ0wyB4oObzq
vznI5azbGBmCo+AKdXQc1ByC8jujsGsd3SKTx5+0a1SglRfpFvOxbJEdze2odkpdS5mrIxZnr0u6
HWF8JOCdH8wC9TXA5AwbOTRF75O6ObrR8yPyv8Zqi+unHNH0p3Gz/dZ7CSL5nGy3K1A7nnSUYBPp
SQzGmlAJ+dEC6p7X1e2W0YsyixKS028PkKCdPgN4IfISDHVPWbrTNZSpg+AYN2WoCNV874+qElxi
XFPJiJfW3eWxAjrlT1mj9Icyf8ok3Gu8Giwcn84GQHFU0QpN8lLbCJlaUk19UB6A8FHsWHO5NiI7
F8lanUKUpggMOxLCYlo0bO9KjZa0wbX8ZMoErhJgmdZ7Q2yKl9EXsZecBdwawVwMVuCkL8EEbgK0
6KOxtPPzJIVIP+3hSwD7SRgLVuPySpDGMzbbl+sUjAaCEwUVaN5nwtECblMHIeN381qTXCrreHMX
91QBzsI3PJqjwQ8wYITOZMNdYQOdEroXM5ThJ5UVkOtyoLcG66zrZZ5f1eQuHVuN15qShnpZZFzL
9vUprMivxVKPcymGUKpFpgixmzWyrrdQXc4W80zRYfWwSdM4y1B9pEkV39KVTtKSZBm+P8SOWewC
91P3qj51pf+Zdp55pqNWVdrd1ARVwo5I0uPeGMhRzNxGkwMUXTsdMkVVmrXK0lQQyIqSH553yOgl
gCIEHce6Z9Fe85ARzPABMfofTBq2CD4NRMYmxrcHIykqOmfjRGwblAT5VSVFTMJAEUYJYD+FiX4T
AAu+/pz2o+wBBHtoB1e5F5LRl6lgHSePDx3f53cEHnowFeAof4WF+9xL6uz5HC+rpXXdP4btZNI8
YqMMdyDqwt/AhU8EdavNFjy0IIVQNJqucYnuLuWfHt8pSliOJSn3APGk52BMeTv0rchg0sKWPpfg
zrb9MraLy0CwNTxOvhBebJcQMegsGYi+j7vDlKrvxx6L0iuD1rW+W6GTqzFuszLR30e5hYAb7Hr3
f74WSuAcDt0cAE/0mqeeS/fHcRi1PRE/h1FWh7eGTBhvxnMECXf0DAjXzUfeV+3ZvnBPSlzzelUJ
jeLM9fWulTSitad5zcnTMcsKtguPXqRw5TzPNlKk1gU34qrd88kGFRB1ZSFWKw5E1L1yYaZ7ko52
sCyxp5wudanTYA3K2Iy99HVtOZ5V2uzh2RexvZSd8UJwCgInHEZYn2uX9XGBtK3bjneooZ64jb+t
7xc49oJQJn40pzXngbqtK6ieKxKnHmuPV9O3WQ5m7S6aHnk0n1j3Zj6c4DLK+OcP5IrFxSlAasdc
AuOLPfaMjh25JrECzRAbjF6acW5yL99sD0YdJbl+kHJ0aQm32Ys0mnxYHKIYncN0AhuRwuEevX2w
LPDFGIAOSiyzM+zP3P2w9WBtAAciQ+ppmFFes6LceV0IWeBk0zFgIt7dlewj/OImgnE96/65xQVK
h5KLyr2TSF3cT098c6RqBzdFGT80uEF5Q6wcyM+Fj8lFRN/jcK+Ibyrlm1hypR4MRy9Gdj6ulYuN
m3p/h3BD9TscM2o4hILWssjfAzrwzPKWIhjy08JsoUSpF1AhAS2CAvEo4fIorLHDJOOl+hcv8mTT
EU67RhGO5u7QhwqhsuRYbOktpAlGjxWAUzpVnc2MdMeGazuI4OZHsMgtW7Xg6wttm2aJNeB8oZFC
RlLrejrFbnqJhJxa6HFbSsjqJJsj+M8w913x8uKeYvPJaxeKatS0nG0wBESBII7vPkp0sQ2uLUMX
SRL9nriw84/Fm7CmyDsOHQK+D+urG1DQe5KFxZbJ6IWHaiMgIULFJrU8/2MFRjAZ8v75AUeZoqgK
vIXkeCvkjUxxNVGSO/T1yhNDxosd6ujcDMIG90ajvb1BQA6vQfqzWkBAVfIESfcvegfg0D4UjfNG
9ItkakCq3PJSQ+DH+aSrjNrU8v9RqUynUS/lZivA/0y9QJjmWDfoCQg/pu9yelndZIhwBdgv/8TA
8I69cTi7obNLym5Rdr7Dhbx5frneh3pAQjsevB8aYhpvOt89z3dUA5oQjcf/IZcNxNcmWFJEr3Un
nYD/K39/dUC2YNF7KH0IMnUzpVxyyLHXfd/3uFt1EUCCY9ufKOp/v/yDhuqoPYQOba2Oh/QcSm4e
QH7/CTsNNI1iGM2HuipqfkYYaYfUN2TRZ41F++o+/7pOOjx09BFp8d3NO0fgZue85N+Nz6WWsY4x
u+qUayKTr2BIIkOPwMfZxal/hg6PdV5jfLF6OPHf26zU6mvBQ+gAHNRxu7GKScN1J8gzv6hDh9Ee
od7iryaTICCXX1IrLJ8r8jN9pxevS4V+vRNT8OfOd13JGOBdy0+kNN3SfIGcGxsoSrC8iVQjm9wr
OhQHwSFox6bgapy6PCrarkyYh4tzTc+1gqLlILvUMRuw/srAmPSdvPs2UBfC7sKZVne6r+TnD+v+
/YlCi56GKS5RAXtE8hpynasYjJE+EgmH+GzTMIiVK87y7aWdhE85ZIM/q+W90gf/L170x1yTKm34
2aMiLXiT/ViE7DPdgK5kBWVsJwpII31I8hhBTXu0JaqbR2qdX4FQjO8QZCJRXeTcxSmFjGUxwyWp
9zMzUOaWEBX3TUf/4JVwpd169ZOuNaCqq5gkr0Hy7Tw/CxeCB/26CTU+prEH/A2krbC+PpmS73hZ
gPe5OHiByWcg2MptVytXEddZ/3N3aUWFUMqIttAXlaEfke14z/vxhqujJgp3XTvLt8KKpH9UzTpH
dfJDfVSnPNZFlYLsZIHW5VuqZYPLEe3/2l98nzdXzRK2JDd8nyPrhwInGCLxCzARDUwlEgqyiAVU
7q/k6dZAWKJhCY+O2QRQsqUFWbTy8hQyWjqxKJZKaXYyK6M5IyJ0yg6dLiYg+jxYLMtwAXwan8KG
momcaIDGwiOphGYXvvFOuWbGTpnOBLCfzzHS8TmwyGCwkpno++Lffe+4o3S/VoUgsnaKOGZS0osF
z9amCImXEmafiLMoYjoT/muWDXWQxowbBg28xH9FpNUeonx3KEGNXEETmBAMxH+6PGpaBZhYPRdW
8av8BqHlwMeNHxaKWKjDj+TMcO8v8O7J7C2uqlNDNr6Jm8O8IEIe1HH5wvYtd5JQCfwtfi695BvK
YdFKi+QLQNpRg3Mz5SmMgupiWuV57KJhhcKgzKW2Gv1eh9sbpbR0f53MMmHK/djHGtgdBH6RbDdq
BtTWogatkIPV+nsAu+KZm+eyegaa17DWG0iP9Ov9jV0AqSf69o0pkVwIPsHTQsCH2dUmIXFvG/pX
57iT01GdIE0+uhfQ6/N2L2h7/zRbL//9ksfD/IO0LQjuVZ4YQDw/tL7Q4FeHWRPJu/67wmbd9uuA
BJDvOV6uR8TKcSXrrDggzfpLPN8J1vPCi5+/j1R/gluOYIKTREX5KbhSppSIRyWecu/xYj6pjEPz
Am+QYCnElxDV6J38xOXY5c6l25pu3mysYBsVhGxOLrdBD8u8iJgFyimaxIRxhQ+HboiLWaLf5So+
xnKm+FBv2ubT7w+i1HpxIMpr+W64vglvL2JjzMI1ocLbUsTM/kcV+hJHmKfR2r7LvJ/8l+j5nUJ8
Fam7kaNLyjxjimA8aouO2S5rUcqf/Pj867VsdGrkwk68pbv5eU72yHlS71D7AaEpSI8J/2C4u53T
P2opPKFV1fsXZYqJ60O8dEUYFsYmrQFuxNPmHd+NHCPjKyrLVmX/o7L/ZBh5dKg0dG5/5z4q4K2b
Ptp3mSoyQl+Ryhw5GE8QzxSmlZgVbPb0uqLF6YugSaUy5rDXaN5DAVUaAlyYx8yKukKOq8p0hOts
anGfugkzF8GeaUtxqRgSGwHsMAqoN0UZ0IuhPbkO5YUfKy9x0cqqF3ec7M/45LXCZriUu0AI424a
QxVxwe2vYqCQ59BnRrKso2ImOpGcbDHVRyU03rac/Hlor1khFZIZRBNwtFlN2yg+q7Hufcv06sFy
/TCB/VBj5fWmjQsS0mzQn+8O7swGLNp/lkXRTA+g6XYDgzwDe6vjMg7bM/luy67p1HGs4WjV+Qr6
aZbBcNuVLavdpZBv0MFNLNMNlr6Y9OQa1MbgMpQ4NmZSfLpi9vIFwLsaXZDBNnbESHAIMHn2I/wD
zHbm3TXBiwwx9SbdJFy6bJIEuKN1gwNk92rYZcRQOKpstl4QDUHGN/5Xp3vXyyn9Zd1Cd460mwAM
VR/97NUyQpvnABxsRAiJGXMk9ia7PbHDLKAqCmxB7pIwBkbg6W6gf/5Ya2sycEt1m3QFty6edqsy
bx6fByOSPOy5bV4VHC0sg1+16gApNrbGWyRHnfAx4I9DE4aIAzOxk/qWtJk/rbFrKaL7A4zaFcRR
+r6e31enU3SjiD6hJQzbmVjoDq0js0llzLdAkLMm7ViUdjNUHc7zcO+FxSur6B6UaQVNsDPs5Vab
tt/rMTBVuER04/j9dID22AkgbAZMbDOqTYT31YIN01wVhH1FiD5zSuvE8BYdUPpJ5T5My4tj6Zwp
+2KpLlfgyyrqjtoKGZWRKk9A5yVtSZfI3FR8y9LzlsUEAvXfRCMDSv8c76wXZLFGfpz4Ac5rqG1I
jbikaXzNHCiuPMwSo/jISM77N1rh0r8cilnqE2Ufhwob2dcSoGhIWnT8AK7NGCmD4bE6S7Poq72c
yrjmr8QY9p09WzduCaIlf681lEGDljwTGXNgjUNePz09/YPOkYdrnj40MrxWdBBFDBdRoBUsIhhL
dUdejBW4IyHd9dERKqppM75bnyMSwoFv6FDU5NWbdvkdvkvVyDfzz5T4dXbhPCl05GhhHxlVRAVi
TiAYQKdWwc3BF2wyVTU7Icj74XvEYadCP2xcttHvYjHdBbRUavWkgZ8LDOM8Ie0QcJxFqsm5IM8z
MnNYn/anEnaxryOjChJl8f7J79GN0zwCVQtl4coK3DjwzVBhBMltB40ebeCcUv7+Qo/AmCwBgg/A
2aD2cUSlmm/VrMScBWbo18SIeFYG4eLTKYdud3KhmyEB6khlFtd2dIeWB2D+8EwE7Aa+I9uGsWPj
Au8NmMc9G6uLdiwvgee9hRteT1oEKad1ESV2T5ybvUY23PeP4xjrkaBfKUftqb6t9oVjseU7oNPZ
PMIBjhcIJ8yXmP1G70s3f3E1wDf4U4kSitTPLbWwUVtePtwAMGgrY0F48GAXE19lEbkyQgIJkkwh
2eli6Az67fPaKUZKpMSa16v+gKdPfSP8WAYKFTTrrjb9DocAq0lVihGyDVjb7yZtHj6DPkLryygu
026MIeD4BmRIWpj5YgAj+ODKi4vgrh75mQMTcWi0Hpds5O4NFPmGUkNYtMADYsl7ylSwOBWFVKZL
T8hzJODOQmZtYdrsAD30UFkbdDUnFOsDm4m+lAY33Ofq5/wqec0+Ttgai4TbCxp7/QPTleFrNEpG
rLx6JaegPp5Sm2VId7Sk1rZwik5MH0AmDJxG+6Cd7p4qIGuHpwDvYno2Wgw5SzS4j5EvxluadYOv
DybDUku68XFXA3qa7UhbppIBH+BzDab+75nyuaOpYeu3EJRuzIaHzTQMQxOPvLWWTYx2c8Y0bQlP
QyFvxOFT87PNHnMXg2I5c/eofJdb61+NJtzpwJQJ17boNcUw9Ka7AHHV9yRL86Kwa5smfulzf0rc
Eq9i70C4UEZnyFZW7HqU6WutJQ8fsFuRLqqBrk4EAUP/tRoRUA+gWDyPpeJ0akG1iVz2cdqmLfnT
ZcTXsCkFD43hfXUwAthQRsda8CByC8fHPBsnSqOMW/fT9C3AZsc5BrZZ/HLC7NcDUJkyUDUTvX2r
AZQcZv3kzI10oBznR/rRM+2q9sdOp2sXIecvmTEkXkLLEXnl6uX1SI4+KZuT4WoPVgmCTFLAXDQ9
nBmgThE26hB8Qr4tjIaIx9SLDST0URdfPvapbBKGpg6F3I+A0sMAmY1TLfqr4Q4IngB6/1KiLnL6
wZDOE9GO7T2X1akDxeCvQXEIFPCJ7ixofGBlc/yo8LufARrgICDofEANJfhv2OlSZgOoQVd0EbkH
rXa1BjAEQQufWbV/GNdCth4OJShylYLFPM3/f3WlxYih8YbzPgaBeDfMePJsSX8wB+eWB9XdWrLH
+D0k/9WOHlReuHsK7TQCDZiarb/kciPkZIqZmugbB5Ormaq4oDWl9+rZVmuuOHQjogDV7nQz+TdF
sEnWlV4aWbna9Rvnz2FucGzLYKqsSZCoKUdoyJog5g1N7DJs+C4hbO5x/HvZWg/mOqSOp1MC1Cco
tR58lM9YU7fRoJMBx/DJ+xoTNbaw3tV+l6jM4qmu5GXW4mHrg/3fADHb+DJVo023p/VoIt7ySgTr
olg9QYP9zwsDpFWbgCdB5LH6sH5KhEYqfAUq/9WGmTJ2K3clLTpQY5kenLLoo/ypTAko85ae1UYN
9m82oTOQ6L3Jvu5r1VGZNXRvAHN5U/TOKFQqojDWUlgAKqPq5EKFlBGT3E0MAO7SAU6TeAXWAjoG
fPQ6HQLIoqW58EHCs/GOHrnLo/6w783zj++00NDcxLnP3MqtCKgKQgjbSTF+bYZHhfx1RKzsZSRU
QMAMsjZuVevFYfZ1un52sxvIRa+rF3W5ZoBru39aMqFH01RKKJUKNdMZ1NwaUqbZjsoL9Nm+zTW9
rgPkicwOmjG/4Y6akDQkp0Fnl7TH7WcGSdbv8fZxH2zW3E+ftiuIMtFtW6L1hc7hlCUCziIXy4UK
1nr/HIDB35rr1oNaudEBmX8DzBnqXokSc2pYv8+lPRKoxG8L/pQMkjyTQXpbU6sShnjmY2xYoKAI
s3EZwmUYQLp1Z2JlHHyUBQf0VrXDkW+fIX5HI/ejv0mVX+dEfvp1yfc2RDbrqsVXIjHNh2Q8wqpy
dAbuGvnC+E+SGBsGfFlKilB2didMLvaNDgNvXflTAhZLf3xerUls8gpbFdVPNCCca3ssbtogZ0XJ
rajUZERr1w7Vvrow6I+HNipcbUHrE8RSf2sZSqaDEITcWQ1UodBC8CO+H1URLsN6lYh07E0VQzvj
yvU+sV0gjApsbKCLl41rZWfZTw9OJYIAidDGhR8MuG5Fb/+EXpWnhsCnQQcA5a1+c0H6Kg/b6vy2
N2n7KCaIPsXBM/j/rvLS2/jqHdioXozzsHRmYPbeKaZKvg2IFI/ZEa1DSS6WlLyY88vVVlQ5p9Ah
8DtFdOLlSjPfesTqw50KsqHjWShGZxNX3TNEoZ93J8CVUWa7SHjr3BRQvH9YM+tbRUooKmDOfdeN
JSA/Z5i6D5IINCxAtETE6Tpbr4X1vJyX68AZWr0CIe6A6JV4oCWPTXmGAAmYJ0MBdJ/Fe7eTWp1z
NlkFP4cA874gzoa5zoF1yA9KEPC5VEXfV91ctrNFYqfTXC0thIBryo45crr20jNyWCBf+3+AKPXa
0wkRecpsXcDeAek3dxApSgsgwtp8YOsK8Au/fRQ3m/Pd8aaY98e8Jlk7DhdRKNz1+jAzpyiV2O9d
XlsSEV5Vo/H0ylFuE6euwnbxJvjI0Qk0HNOgOHr6uO2J7Qv4EAreFD2I4Yn3D0IUREbif3G7nGoZ
SPrFjD9APZNlXajOMvAZfgLHzKLCEJEqghNmoGWrVsIqrTrnGe1Az7nj2I3jgysc6YJi5WNKQzjL
R3EtHtdzt49rnQr7wHBYjslpHHUZmdaECLkx+w6uywiFUMibnHfa3jOA22vZSWS+QZqOQbXh231g
DxpFHIQ4v9suPfdB1WFPPRSmDFbHk9TvzP/2F12BzzP+PfMyA6RhAts58y7Tv+iqUjLBfkLq4t++
HOm9pkyIxv1olzaY5X3Nn9gxKBvrhgWRqmTKpsYvGTnT3tpKdq2Exn5hDUx5OwhrsOMByEZBsAKa
tSflWULyBp19a7Z6wvgFzHpHae+zZm/57GXvT+XPGGyekN+6KaVdeCNsTl4kylD7PfV5XkHlLE+9
2B3VI49OZngmGjfdwtv4/0JHn3IadTuTvgSe5sUl3HngA9+F6k52dxRgl2Tqk3MrCcwK+dw/mXGB
SBgXqhIIolHZcw36LBAfKZzkPyH9WYgm6Baf4+T5F27JkMkQlL6B4E3ox/RCr16bOJzvwY4u0+/v
cqibHv8KjUBOOskakH/CMZwuPZEm5DCS9f7byYK41PPI30iLWhrJ+Tn0ad5BXXwDJ33Lc70Rv1JY
9L6Cwe/KCtodT78k5jhdCRAW4A3ee4X7OeHopVVq6MrWZ6XY6T4shUrD52f//1+JEwqvcE9s0aJO
6H232HHtg7gE4Zn7MR4KTuInQk6fi+Dd6BKdPWol7u86JoLIKFkTe93JRi7ayrS2eAaWmnTkIztR
bi4aLlw5ref0jMjHclS4pVuo6NWJ5+r1ysYfH7TokbmeDzMGKD8KRB+brxtyFwFxKlq/dYxsuuXP
s1XvAo2VjBdJF0D6qncJGnBQLeZPKRdG2BjR0bThLYdQKDBzQVbZoE0n2cH2zDHhV9aM+N/Uz+9a
Pg4YDQK4esCrvF20B4bh6Qdjv/vfJ8Kc9X6BpMPuMtM/wIeDmxfWGrk89h2I2QDnDnHhXyeE3QMK
8p/PLkoddzrRfIq0NyxXl+Dqc91QTsLxjYUcEcUTa73l3E+pYnszygBFXpLX0rgUYmhIt1w3ICUv
E63l4qqJLnlmz8ZqQcPwpv522F0NPuEACXeOTebzr5BiFYtcz9Asv+RSiO4tXazZxGyUMw0U5t8W
IkH8ekmX3uhB7wesdM6NqYYLLcRO/2A2AHhmHU58Z7SNFAvc5SkuU2QXrSLxAoqRTXxqJohEVS9K
GPN5+RMKxCUoWuq2Q4RinDna38vsns7jPMlcFs6BrZJPcY6BKbpdA/fDvQAkwXo4nnb7TeW7ZsRy
25mrRtR/ceWABM0p/2HVu74+h6mPuzdjJPmE83u75f/ADT83kEzkL515PGh1IHllVk0NoG6tfTg9
Y4q8/H0apWKs/6FtOmzrQ2CWAUgPZ7O5E5Q/+eB8uacq9K5EXkofgPKFDtsafzMCihlsiu4xanU7
CjokUJxAGscCi9HAUDzss7vMSXcjwQHv/IUwoLRbnbKS6oRnDb/y0DLKpg2XFC84oJyplEOmTSEy
PaJEjJOAugfbLXSR6lWbOBOycSSymN+9Qhsrr3AraDjzV0gZVgg+q5Q5UAVySKA7fG1FAutjAeG0
6pLpIJtgbe5qQ9Vthwk6ssKI4Wj3Tacjql0JETcEGMRldOZYvmKKuTqfkAOgn496aRWa/v0xspSa
D11+xcCPK/KoXAKnaL5W6CxCVx474MnwMij+FEsoAdTBz4Q5SFhqdbxzLdJciZu4kGqv3fUj7zdn
9rk1yFaDXS98SFapg8yCOL2fMQj1HBV7IX5WXJGRycc+YULR3m7Axh2OQd0G6QKqrFWLfZZGcsQe
pdDLf3S1L0ty2kZhFeDp3NqOWtRsq3u1AEe+pH+Na1lqEsMpNZa5ra+cnJAWnWxsuwXHA6e/fAXv
i1X5ScBSFSWTIZCAPPQ5Np4p7aiA6iG80ODzXK6ui4wmMkcVP4vNLJ7h+3P4T6q3x3NbHG4RwpUB
8bcRDrz3IuwCNaT5XoaV5xzzFNsDC+7CAC92Hc6P+YiRpoi3FWzNOy0jPiDpJRlP5XPAm1SYc97Z
ONw8rjazDEIEOls02Jpbvezstr8uGJ932PWm1tRqkbHvnihi1JhSbyOLNMku4WvIchLQQZsdXRSL
/xIkW26Ki4HyLVxEpElDbrbkbE+9WL4ClWoclZ9+iOwv8hYwYscnW917Gb8nVd4mfRCxI8DECHag
Yw4CTq+IdOZ2ozaaXGGRxgpkHuxRAj4f7TWJLGKGx22IJk36xnmBH2Z8JD1Hxnl4cc74VWVQlvdd
Qo7WEJGLPTTykz9QPmudcsf24FcQr1rOI65mnVKs45wFCR2n++JFO/2ZFm70qN84vpIick9JR+6C
H+eqfkH3CiVMVYiE7l3r0LNwrT7FPG9eRo8QQ3K9u+q4IaoSMANYcTuE5zla/wSM9XpXLqZjctnY
NUkbnZvqRR57oBkMr1ufaso36V/dp73C/k/L64bag6nsmgbH18VG5sSxHOz6yGzdk6QYsdm5+cMe
uVdVbmQ9zKcL5G6kjQJoM1klFKCyutU3R2t0JPAejDdA2adRIWixGsuXO3+9OjOMrO8zjnQTHlXd
TlEKQ60jJN8ekarZb6yplqlLblHcEzhjD+jrSqn/+4AXOMWmilFlgCQXAyMrxuJrI82ukGgvWkRS
s2j/QB6VYeurhQejkvF3Yaz+tQtck5b5Vyz9UTWQUiQoAHiyBoTR4MH7IJZjId96tkxIGrarX7wF
JVr0aLxd+n7s60rFIJsepj2/Rv/NCyxbh3fphimwvrTtEEoeJ2KUd+9xg3+giZ2pes9NtPwqN73E
U2RE+urZbK/xgnFEUxO/0o1cSBDg5iVqNt4c0EQRhqnwtEO6T1N0Qn0YH9/OkTsX82ALTzw+ng3i
M5nBhdQUNDGtPu0pgJBNbIp8g8UW2kEBRDKN5rOVrlJU/l9BWTusk2yqSFGyPw0T55eHaT7R3ZXp
MoXPlzk3rPjeDajikxybuc13qePwWbICkUeW6fW4zBTSyKWQu7xZFxR1JKThYsfAYwkSMz8ME3OY
460NgnTbQBMXGhatEIK6jk9Ul2PrYI9vykXnxx1Na4DQlcXRgFEkK0uFSl5Il20LXMEoknLPktoJ
UjRDHjlb0VzkmuM8ygco0MotE4vhRO3uoB1knJrt7wHDckDdsY2zMFfUgJCiIUylxpB8Zuv+llVD
8kacAeVMDiuP4lnmS54gU/EH2FsPpx5E6rhobGURs8ZcrjtOF8ALGWfZq22dTm/Ec49xpxd0Gk6K
d+eFE2okEuDqz+XNNgo9fX87wqADfMac5Lt69uFZ+i4JJuOeWUcYtfNQ1QngKxWwR3jPbEqMpqoX
nXaQIl23iQ7bzTeLVGFS2CTo461csct/Mw0A8UgZzMjY8PWeDbKJuArOkgjhfwEUWry++QyuJxhc
GJW8DdmbkkAMoWTbG0FF7r1bJ3eq8ZkXwF7+/AAMkDA7IwF8nEucUohGEELnVHsvHYBlrJTR2vqd
Gp8XtJwAAH3rXT/xxvfCVLBUxZEN8UduG+fiJ/r1Cuaa1mDTBJyIgmc5d1hpdbWUWsHdgQrWhNmW
xVu76MJHsaIuYQRQpgE3QiD2NYhfvF0b0IV158NkpMzc11giCVRu9CqAvyHbJ6fRwKsBUqyN/n6Z
USsl8W2lqugGwYbqQ9/rQsmSTSgd/Uf9CpxZFmSMX7Po1d3dFxbcFM3IfAWvV8KWj3IruBcZrkF3
2Ru/XzXrmgZmJI0/xvEZzk75qWbZ5g9ePHEfaH+sxo2uPacufLmLed5ixVWsDxlFv+IUMCdktjlK
Q0M5Q+wWeNR7W/V9Nm7P+wWJgxJLtppLFDCq9Ek16YGqzq/jCe8dEGm9p0PT7HKH4XQuAVmZ7o4d
3le2u15qRtUX9r3yOAjMzTFtZgvC85I8J2cxQOKTtJVjvPhYjOvnXp/TcT9rH/s9Em7Sw1gYAVF7
8TG6vpdyY8eklsCaE0U0HPv83uDuRAiH+sOmtbfuijdgDEcTa0PEuSZlO6BVERDQUz+PLSQRQzf2
iOhvR4F0STRes7SmLuW2qcSh+7gdQH2HFRsnou3KzBX1LR7zXFWZVqDmqMiE+UxMKJobPz7JjiU1
kcqkqI8+7hrtGhlyZsQSWz0Lf/2QFre502e2osVqMzMs81tPbfIEEmjezsi7gEXrsMBB48q7UgiZ
Mdo7zaFBAVXIgfAVQI7ydT1bqXDj3uFwkTWTzeDZrmCGFi5z3Hd3F6rtaCHqHkm3YFLH35LuEw+h
1OfNn7Q8IZJmdBa0lsAjmeek1MZUKu9w7oVCcQBpI8mK9LrvCFb55CmRix4alxmdny/W24TWPLpU
hzJBovddvMxu0m7oJJcIMhwH3Gx0ntVJsWhbzwGfXHAw6j9R+n4rLImCe3pJNtZfJ8MtK2YKYKHe
L1jrCkwDb+8T8nPBe50Z+luAUY6PpYcDiKLlbG1Oa+MGapBYqSRPVNZlySPMWgWVsx0tYs7nuGc0
gNbJ5n3ihfWcHeNqEssYHEtDU0+CTaTs3AbnXZyhOI1r3bsBa0jpGoWowec9D4yw6DCzF6H6KfHh
l6pWVvzPPhyU8ADRUtTAwCjd9tOr2/3SxoHAdEIKfdlQLjyDvgFtvGkZ9np29U0+e543PI00vREQ
Txzlio/CnerHYpr1vQzY9djB9/IFHDMldN6rrzStUtMqpKlvMi7Z+yH8PIvraY2kpltTlUtaVH83
J3ti3MxlSd2veDc1wL8+vQfBJPIXyHxl9988vUKw2fIA2pL4iC/VYZTFl6lUxz3o+KPayh478VE9
rPRoqXH+SpejIotI0oq9aUoYjwyoJcFKgpoTWImefyvoUNUA4+MMSFS1gCXQ0KNUjk0XvOXBPQf8
Zl+HDVtdtPztHdAnx84as7F8MgdP48uAfj/gJXDsBw0X6HrNs16Athtkdiz63P+OXoID1pCY2z3M
12LK9LrU9eBGr99JOozg96dLS/Z9qhbN6IyjOzTImsAX/MhzkP4Ja52+qNDDcDErrrtx8MoRapKd
JEdquBMAnb4LuA+pSDuiKB3zU/dLpNk7lN1e3c7uhnxA1/PrEgnNrIb7WXnOT37qVJ01RmVupQ6z
rv5N/W3fCiYHzqt9KCNl00f/7BwiwZdtLLFX+e2nmkcQGgSjYnjgNzjHHoyFg6dsTMt/onr8YsGc
QVLDxDe0zkHbwB11R5u7iEyincaZUxiYvdI9SaQYbnmAnC/2ui+E2EwNsFPQN5/RN8pGBNRxs8FA
Cu1xaqPP4Gdx08zHFGo9r/SPrzIPRjpLBvUXPoD8niX5Eo5fcOxWzCD4r+YrPAPUVapGoH2FCywM
NnlJi1UlYfvPLB2/ZjlG6z6ln4QLkKi09zhsEYHKIkAyStDzg3+hu2EItU/cx7tkML5Vy6KMg9LC
lPiZruOtl23QEg76zPArJwUztknewPFTG/4r/ucHJ0g8aKkMbLfIQpvTwJjFILfFw/sebOQzll+1
GqdSnIT75MiYRSE/gI1DUNFf731uOcWaRxRNL8XwPklBCCdrFC/0dPnuUBsz/t+KVfEp8lW/N032
ugomjQo21yNNPXGQW054yCcAdrvzAJ9Rhb5VvCXfxOQoL6KGgJS1fN1kUidg4dtssQX0mU0QmWPl
qDnyOa10LaF57yZ+bmXeNwKoJYBTj5sow+hH5Qby3xLe5MRRhGwVRNPxaFgjKJMaVIdx2yVBa2KH
T6bBJnIfYjEHNXeh6NCPPYAYyNKyGH7ZSyTdxLbfT2fd/CoJIseZH8AQnZ6t+JipZ7Flwx0VweFJ
2rOpZ9twoNTA+OisJeKPU8RA7XGhkP3iMsmwKMVX2GCGG9QMjzVwh9cag6i7914K5J+PKf+HAvlC
cAfoRdYIJfacyVFI94kPzLA8sOIRGbudvgq+tSFTa0vu8vYLqO3i2WShgkI0rz8WTZ+uZ+STCHRt
QRL0gvcD3dnmWQ/K5vqALl6v+Sf7z3WNAHF8e5yaur94iVoqzt/FC7dB+JtOz/1NBdzLXxFMaos9
ppu+Rau517Oy6e1CUhk6wKbTDUBma+qZ1NdI92YRykx/j0xHyXRM+xcNGs0+sWkpjSy47/lvGx4z
6AlvqVdIod3oxAn4LqjvIqWwbsi08Yiof7eKxXAgZ4/1Aq9g4qV8Zw8rVVzuzqw7C0IST4tJH0Pk
0zNvyZRxSVok225kGIsIMcveAiKRsHQDfn25nBs9eXVbRzF7M9gmHGP1gGUEGHyctObUQgnpG4Zl
5IMUlwePgizh1K2KqN9RVQzn+BNrAnSgRqfjLPMJH8zBdxCMTdP+aXdoabkPnhB0qSdokJ1iWS1+
lqYw9yLjZ+9tQSzihR+6af3OwKyfApHsd1mcxX8D8RBUajPS0CBuXF2OJRvjRiDdYPl8oofQ9wfl
nOJS95vDjlA4pYcwYYY+UrZypGTfI7oecAo5SnfBgRdd/8DAqKx9KTtBy4C4NIaRqZlKikrunFaO
jfzvDrSPZTIeCXemqc/Ceew05L4dq/6JRULMODd6COENBdb6liOszFrAGMgfKHDV0mkIYb553htI
wQIhyEbTe8aqxE4+gzK7NGZQiqSUp3pbP2AcAtrmcoEHMhMKw+xX4XZIgaIEYUxFzi0uuu5vsXQI
4taJI5crwoxwh+dPC2wdGCFE/VfSEOoANue0kbzerfV+0lBD5cULmi+rkIw1Jppbnia07n0e7zKo
6bgFjsxt+PaTmG0tKBvuzSF48yEXzK0x4o0lqvF7+Bh5u1xr+pWGuyqx/NDpkJ+Jy0rRpvPg1M17
/2e4UbgGobvvpMN1OU5DhJ/jKpqEV8N6EMlyWbD3Pu6CHehWpmImsNpoJGxbhlxhPiLcfFAhthX2
NmLqJUOlsID3qZUk6J0qBbxw0Elozc8UHGpS86kqekuq+ScYiOXyTPTd2eyZe1NanFZ7UPVoxRAJ
YvGp40b/+Vmz5d59RP+DUbPDIVjNbWbXah7ubPx6Z459pRWBkS1zyHfahyLgJ0e+hURb5ZMDObkN
9bSXBmx7q5PUqRJhZFXr8FYtVj+6qjZte3RZPlHGr3nFHWkqhzAwSyb/9nOKzY4TfG6dTiJ3Qnn0
S+33uRDeTVrwxTA4fRiuahF9btiWtvEVPyye1AibvPGeK7hFDdUfi3m6kB8swPHImx1P23cYCHpS
90pdxvf/Oc1T5hZ/qw6kKIe2Boky2V7/3H0ev7lmcfQ3XRi+5fLQoH1r/gP3f+6VTLLGa7x9yKPm
D6kWDP2Ses2K1LAO8fSF+Ibim9Ou0fSqvgQJdtsO6tAFDVtPhZ6reQsiAeIg82WzHvVQ67xEFnBs
Y4HdzPHF0AfVAUaNsvyqoDht6qVkuUNy8njQDW0xFUiGTf0jenMytF1vlSVs7bmQXN7xzy5tAMZb
e64rTAe2TnFvldU3fv8WOMb/wVLXB4lYjz0FheHrenvFLoLQaTM1j+b7hoYAlC/hlhlYAQPQu6OU
4Nf7CQc1W2h1wOHEgGnGhKdhfhAXZN3Hs9qvlRVmnQ8prsu6n+alUvWZmnZprESxKXNfnXEbeWNv
PPHfykLQ58iHOUE1YiUPYc/rB5LcYsyQD0VW5/ksz06sYdvDN0nqa+9MYwO+tWPiVH1BrYqwck8u
KFTCGH1g5xsRnugBcISDbGwwxlKFss2GspB1hmbiWE+eSLY24pMGnMdA5zwCRyNcUDztLeh6ogfV
E+le208C43E82vrCiVj+rfuyiYgPy8WKwYABeXPOolt8gQeEPrNKO9CmQsevg5v/rc2K76NMSO0w
YCSmSpSX03n2aZrh4iMV26PcouDrWD2EBY/KGxAXaY3O0Jpikm6KIebbBDDs5EVnrACoIqUcyQMA
QdhfITY+dTLWry7ssqlkuxcLLEeUscfRBRYjxer5IxKxq4CEKR9yG8qDyCaoZzf0qbVD9y72cqoU
+gy572QsdTM8tlmXnY0b3GPDi/LtxoVdrikEAkedhWzs+ompAdSmACXHNL2+XfuzqylVUu6ajfi8
DxmMpkeRHxJT/r8KqFdDCmIbI+7TA9BPPLNXeJGWMN1YiCU9506x7Qq7sTXgDNGgkrmGFHxx+zFc
KLub9jWULZAePfSp9Y44zYEBsO0miYgEH72+K4YGK0lVJmq0ITNV3S/0YbQ9nBuH+xvTmgOWqErD
HchHG54UURtxjXYDOuut3N2dXoIhQH4cP0An2Nnfjce+4wd/uvABKc8abSMah+FNyNNnXlmZEKG5
77zfsK7LSg1j1wQitd5O2BMyYvLrV9kLZ+DX1+V0hskgQ49hxdEuRBCLYrj1U4leYjkuu5K1vkD4
6ZpBxVxt3ljbR5PPeiU3ykyDef9YmZFFLqmLIMzyZc8grpdAUzIvaSRGWyrWlyQ96UhaLrrf4UeQ
GWq4m6Ms4rd77yNzJz8xui+pTaAMq+ysbEjXUKjuz6I84zgAiN6Ey+3oM084bCGE4Wbv1ncaSzrn
AgJSs7VVYk5Kcas1tJsrln/CSxo7HS3v5P4mUuol5+byAnUKppIc1SjyZ5XseHi4BLXdYegYgke5
Z9x9Q2cjcyAnTYth+3uy8fsix8NSRN2jcs8PrO536Oy2sVcIBtPtyU8244RI3ynYAbP3I/Z1WErz
vMa0UbKgvsrBgzmsXv7JKsBHcF/d1ZqYf7DCB8ulKfIOXo3H5N/sCyBqT1cMVwbXJO+DpKpzUoJl
Qlf5pa5+hmL2KggYM3adC0yUMOovHeFJ9o/qYhZ9BJtmJ09JppyM01pXUyfnGIzotkhagUI6Drku
oVIG+5EdgigLzhs4Q2Vial0lGfxs0HUDghH/1LaOUGya3amr9kxNNmSn1aLhOUHU96mXOZZqp7pC
66YYn2eT/o14brHLuXK/NQwky36AVPep0DrNoFhePhb6rWb6jjfbC0EQ6lu2Ku24SJkN3NTWoON4
CB3jzIyvO79dlbS0wRSkBwh5Uvi88T6mgSpyki0lvlzXGdSwIgjsahK0EvEKttXlQEgNeg1Oxz6H
oBzT7LEfq0z9Ho0K0vOMp8t2/sqOiUhi0MPQAlxIbYWXBI9W+FA1WY09APUgi9q4QxGOYgnKw89U
MXY4eEc+Z0nLTsNWvyc0p0VkpqpIrbGthJFbVAc5CXLmvORbq6uInIbXyeW/CYF5gnYh2WFYSoCv
flkLvcV1khci5QZqeE504Mm5YVM/vP9dBvSpENupefUaamctuuJ03mlEAoGEOv6x1iN5pjKMdzLB
wOLolRVWfMghC5TlO5XWT6UVDwXYyDQdze1xhARWpT9ytQF31D+QlUOjlgoNHeY5Xd0LSjHIQcXN
A5br7RFrfBO7CSmyKI9LX6p3nEN7klhzrNIOUzbd04CKzHZt5hsQ5yOhQOWwFLL9KKLToiD+MpdN
RC6NL/Tj6uNqUGtCwMgmuHvEScI6+iOk3mu6790mYBAffv/g7AWzgOw23i0k6qhkqT6+lDbkayoJ
pZgEvK8bm9scXIlJ4Or55BwJBe/BLFZgCrANcaKvg4yXTdcdux9CBj01qYBRCIGdjt2W6ILd8mbh
iqRoPpdlFdy5wLcqnuhR6STlVYxG4sPQl92+Ad0Ljtn0qPZZrt8tpWInX6NoXsEgfCxuwjvB8px4
eSc55RSL+cZpZKes0YLE0Dkjg5CSek9fCMCRVtxHtg+Wvhb7XDMTWXNqvrksmu6OxLOTwMpVf5t+
TNdTq+EDP8O1GzMZ4nkzqlLeG3aYKUbqlASwhRRDgtcEMqwGGi6nP0hFI5aEzU/R7CY7bMcAsXDx
lwBrEybGtipwvl2nzQ8R3vzeK5paOBkZO0qdhmkEHpHQQ2a2q3W45b7N9+MzmmcjU078FB7nDilh
NaihnGJASqBEQoBtaSWAzU30saR1M1eVxsXdMeRfW388rivN6etcc/Ec3vY7nVJEtoEjcXhrNdIc
19DC2/lbWfGV3N8HcvXzLwKn8rPS4iYDPIsJwiTNNXEZgn/VIN+txk1j38M662Z/PINUsWF5BmIo
acfElivo3b3+UkUZ01PbhhPXCruO28aahHKqRgwFFS9zwNd+O0UhMYAULIYYfxKYXDFFvnsHrWqU
ARlS/B7ixAh/diZMaTncG49pWGXGFXMzCSx2v0MDbrnzDmLMfQgaE7Ib8ccpkIbPdw0p0tKmZHLG
otQzv77B5buMr3L0Gh1Q2Pwv0sU8HSqaizUV3nbvxyTa1c8KN3LN5sI81oMFMMuV7VJcwDnkx7Rd
01NfdxEeMUnfeyeU0I7Ut+Aly3Q1u0Yztem0igvgS15Eki5da1D701Q5DxgcfJRBwjkL0LMdivFl
hRnKV6RIgazPTxGpMQBex0vg1ISDh/M3Lh23kKmxjEPQPHs58Am0s1Pum8GEfpgxFJk5PykSEm9R
131wYioliDGe4i+MArGfRURjCxx6qxH64EqoPDjs/g0WR4B0abCZMbBcUl9pKVAxdQQz7gFW/3Zq
viO9oH8myMwofHbI3G6/dAcEkwOW7wzuwwZrPuYNr6A3mUoJSDdGcI3T6kC7N8gb3zn8687GNNId
7rYOsp22QTRBKVei3vYKy9hA2qq8xH1mv8unq2vjf35p0z4jV5eNrTbslNFNIhFgggs86D+5KIBi
BRWwXSUMuItFB0sHQnYutG9j9lAg4/lXWyp5He7KNcu3IwY7hlGxMMmCYaMACL1NEn3ON7MxuSnd
KYVeEHfCWYlODuV0SvdEOCothMgAN4KSgPeyxxKTwHcTbQjVVdopgLJfL7byRZLTVyBQ+fCcuPxn
JsO4DFseGMyOQZKHpk2ElXFDCvkbaaLFFXsUJjFic0GOXm/bvHP9ohNpl6QcnbEjDTPjB9FW/BSL
kZmpTvPFNJZw8zwB3N+lLXr7GGihIkZnimLrVWoepECI77F6iE8VcXCgVv01LbrIwGa1QbJX0ztL
oStzQ9DucWWg4UOhGkwut9aJguj9tuo/ZIL5D86t9U7TVPLJdyLZMiAntIFw2HcyM7jv11rACkWU
fySsBHFMcboBfpd+gl4i0J/TqQX+7JlBzv4u3ZvkqXJJ6grdZoV9pn38T0VK3D6dHHgzqp5hlMi8
bgcDsueVTQYDar+p7NU1UZzCarUeWly+QOjhRCptqNgXNlHZSrEJNVuclp0Leo+/Taukrrn90G5A
TJYEShhv1tocuCCXpfov8sLA5ziSp2ndfAxoCIJC8GuKCzSplEKB/+ycN27CTcmCD4zymx5Lp8EN
2vB4Yfp1DlRw7+BBSClVvJBvBI6qJXuh0D/Keh9N91z2B7nR4rrjgHJRzys0vW64BC+7N4UEugg+
ViugWJQ9tDYSHhmkek6uCR8Bz4TaxBmA2c4xwVw0BiTNpNnYJ5kddOa4bvrXuIaTgZHY7fpz1WlB
1/sZPUnfMaDpP50dZebZXa6QGzfDlvZK/yesFUbmiVjP8PRUKvI2LCK8TkVAVwA6CS2+EgIMulXl
hDZzyyzw3bcrU0M8sLA+40HITyCd6Su49U0k8ZPlxPRItS0EXyMdJo5dh7LLYxFFsS2b5mTxBZGC
Va1PTuEX1/wQZ8cJQFYB6UJhd4eUeYv/pI3D6tBKxrW7RmG1sOICWhWj+z/BQeMzceAWQ+XrvBqo
FmmaAxaH+T5aLJWDagOgbN4Co35rAeZpK6oHSiA2LLKqyhYM/Gg4Ljzfc3pvJfPdOOrrn6s/nqyf
9Bw/7bI3wH8FNslveTUGbMSM/66y/63Vuuxzpwv17FBY3TqnubN+wbJutTG7X8KvS+fq+7YXgbUO
NKMvM1ZNiM8yTv5jN7513uy5CPQmYHWWZiDsS0WS8gCP6dU+MbnojRJ0LtzaRQQ3GwEIRHveMx6p
7guZxhBASs85lE4tg3wiMeZFBSsmsXRGGJVVQdDfzSR8j24u9FyTBOZTW/SHLRzgUFuqxQhdgO/g
qkNZ6KTUzbTCCdeoVNjSYzG3HudKCWpHSE/yOWtmWvI8zgvLvE2qZnCD6y5gboQ8dFJwEg+TN69C
kHftE2MxolhiVamLnhi+GNJk44YehGj9OPdWDw1BW6udwXWl7Z3PMGnRNMpbJAeJTOOUFtygBPpq
iHbff5d8n4AaOHjmwFQ6Y56KdUlpeYWk8GXthrb/4r7CjmEzqJHPmrCmHIuwwivmVXK4z7YeUcpJ
7EyXCpbiQPvipnCjCIEJ39KBa4TfND4u+aDYZXoILj2PirrsuIkSwsdzzXazAM1ddTIbSiHrNM2M
VVPudU799v/5Wle4/oFjiuvGQygZqHYXGUVzA7wKoy3VYp/+o5Ie1ktK9zCltHzUumwNX+Yj0LQO
/T/mJBE7Ya2yphRpCUSqRfrVdRXNAKTb7m3Pe6/MlIQRbCBm33pwxFcMEHWmZnWJ1OHJ+fexgJdl
/vweXU/OdbXxfHrU4c1tgNTFnocJu79i5ErmVTxLi6nTkdvN6I8qbJME2GGWuQriPmx3X7xK8ylb
nem8U+Mq+C/o4WdMp3B0dfEkqDC66QIMjfuCHI1aAeJSIe1UmscM3HsIgBNBwDtJg9x2cxOJD/YW
6jGaxS7prD8eY75NbUaoWHLOjPP/Em0zVUBqzGNImACohrjR1Ca+QOqt/PlXsQ4/up/QRYD1nTBW
QOXyS12TbTTDWRaQDyF9nlXmZsxdMnEIS+aNoS6P6PYasWXoKW0vMo7Or0AptxLMnh60oCQwzu+x
j/M18sJaFSEWHeZPasU38rKs37DinTDX7DNqQlm+fHQGpxtMP0MUEwFPPMY2WwFBDfwcC+D+lSWt
eopz2KQWD5UPrMCYsypcNvLiFscvFGFiFljPMvWVVOFNqsXtZXq9/HZHl+LsaLodqjMHAHJd7wd4
rsz5QwM4wbGJozc4Y1zrPVzXk1O21kALIOgJ8JzEvhZLpQNxT19yZx4SRsvWn/YLuBmjaN/L9zjZ
ZK3ifNDCjf7MGT1kfIJ4rkP2k3tWSnhYlv6PXhMjlD8kkiL6TULYcU4sPNcT7sjW5gHgpE/6p/Xn
1x0y9kyk/6ySJe9bHKP6ZJkPqnkraHod5soKm0vSsAZeB7NaKR6mH/iAbxCidNjrZJYR5+3bn/GK
3KtT0++zaCmVmc8gVWWDb1cNMzlncTcwcB27dPRTsHvr9BVWFYrOE/+l7e/HWXco35ZzT5CzP8XN
4PkNmb8fBh7M4b0Z9XNpnKrFk2o2SyJhnmfHQ6qk9VFmALHlxxR34RLqQ1DU2QUAOPwZckiv7QrZ
4fOuZdtU0MHmcM+S02xRfAjiPrSF1QkQeKdUKd4Y1WoC9ub75Lb0wdaLIE8xl6HzKnvEGhVqRfPl
Vw4SDpzN7XbZfUf20yNcBE7wWNXHqc0TAKDJXAOj8gn17Ob5sm4Lj1Ez9ai20s7emDPtwYlb3nvw
xcCuMpXEnZaf8fGqTniMFbxEzzSEE54awkHyQpZyrevaWWV3nifvW952/e8+CxI48Z0r7bp7gnEp
cLtLmOW2Hi9VapzAkihhxggOaoEm8/yniPTM0EWhdKeA0JPgxC6TNWna7RC0j7EwBxYuEqWn+mqJ
JQfP0gzOW9cSlh6ijO1nnDtrROgzHouqBk4ZJSCm9vJZoJaPeIqcKYy2Z1kdoV6ChPx9OiGwRPb9
di0G6ZJ8pnu0y7H5Gjl9CSDV8JMcklb73z0UZiQlbchkxEuwSVU3ZplvU9vYp2wmVlKN9V//3qL6
w0go1zOWoVFscgIL04GnEnIZEqZxSjnYy5S/9GbbH+LXciV2qNpp6uFOeZDXbADv5wJSvmK4VZHJ
s1WJ0qPkUD7uazrh6z2xhOfhRi1Wims4NWjOBSGB0Pk/zARTP5iWCX//zI8MIYQAbqZazS+c3Cuh
mhSYZPZKENuSYJ6qUK8TRwYzx40kYk0XPDaWOo72cPFRjMFrd8PqkSPiJ1ncGIx+5TWoiZSOxAbM
bhm3mbQ+CA87XPVjkJ6q4dE4fIiKeYt0s9PWux48CAsZJwWG1TaxMHU3FXzbfNcYt3t9rS4yt6Xr
c9DgKb0TGDJx/39GhaYBrHDMOT2r9q7RKrmguDFgE4PoYFFwr61KIabumke0+OPTjsgqy8296q6m
ATdwyVdJ/3n4DFzNZtxeEe1oxlf2fCEiHl6QNokc9OGbgfE6J+eizHYqZpg7Hfi5nax0mPsH8rZp
/WhXjIpexsRgQ2di5Ew7yAyZuZrFyLi7cpSLyQ1Vk6u3k/oNKHYVQeNtd1jF1IGAgJNXJ98pTEp3
3mK164NGvVlrnDx1L1+qd01YwMsDgHyCQcIY8Qnt6zPXvCo4o4YjnOh6qLdj1ygyy527pK6t1Flx
uwiMFHfv74DEOneAqCgRDbtl39ax8SWb2gPbZ4WB2bynll5BU7gStCcrPpNtbjjrM/gFIooMyaVv
0pERZ/aY0U9MfoikOUu1MWH1zgYK/3fFcWoYpnVClhYjAxPiseQFuab5gVo8or+vzRZk1+JYTIRP
9KykaKSMwmuNs8gt+eKk72Pqmsmb3lRP1b98iaq4CdVssXnP0bBZyiZdr09mY1f+BpsXYd2osv2w
Gjp13GcnSHhvam+NTwjDGBP34gJBLLs1n95dHP8OG8arTy1nw+YfhkrliPrHJlYQ7vgdWD+2pmMv
dfo/u8wfwGX+yEtFKq5apzMxMBfu5Hh4aVxzRTqtYbZbd1RM0mpmRdCv1HdpLhpMzd2WDR0bZkQq
qEUsJPg0PAHM3X9iVPXufiKVdtFf6O+iMY+Zr2IW/P6bKQnNzcFXHuUNKpR0PXYXfEdZrZB8uU7/
kL80CTcxYQ1o4Iki9U2gs1hDTwHY3SGx4FhVp/YZIVGVPArtK24byZDMwfHlz9ZF1iaihdMU62h0
pbrvEVlEg7ah067o3rvkUe2SvJkzvvZ5NO59OXs43g0TZBcvuR/N9hGdoUch7nfPkbSethDvobhJ
qQrMfnNVJcfgo1D+F1z3PpjI/Y9mY+W9mo2MNfwR98on/8DBmnncii/or5gzeP9m0mt2RTbOafDe
5VmxizqIakY8W6JDsUUPWJUgWjGBJPZ9vFmzLsYyp7vtgyEnk2/uRXbrVqbC01AJGvLMz4aNusr6
AdEJAhAXODot2g41Ajvtgd3FEv6QokHul43Ore8WOY9p/qH/NFcqgVVdRV1v1lC6Z56lu/3xDOsk
8r5df6JqI8q/DkYoIES+bBWUABstZQWh5pRPeaOKZfN9Gq8ysnONQFdW2jaNkzZhztwd5MoN2j2j
F05EyR2sIcGmcsasqj2ZNbUtDOT/relDGnxbXMcO9tRayOu9sTHp5hbOpBFiVd1tCPw+7p3Cavy+
P7A+nJagOJPKjqDa/XiK1Vo+NyuXOIgY6J8CxKwbhsFLR6gaiPEBiJeXAf7VEupPFuybS0GSo2Rm
jk3bKojsFm3d2wexgAEXmyc1DhEI8B2zYkNH6LTLyJrFxtgquZQg48xuyq4BcCGAQACdeO3eKiLV
towFQDNS/ev6XqPgJUvSxdikNPcooEVdr9vq7tIagBoo0qiB0RWyoDrtWeTb/na0oL1EYOMKaViw
qyeY75N9JFPkEirz2n0yRHy6DIRHeHbTQ0JnFdXN8WnUoxoZpRJ+zG6+CcvVkYQWzlE0mxW86zv1
m9m4vDGZBgLT4sS125Y7eLzw3YU4HqEd4t8nNNeFwejWbbMY1JcKQBvVrWSoncZXIUYDGlaZSy61
Lo78BQJfTQyHtwtMLdDQ1jK20IcJ4cKwgvWwFKf5zzzWWIGmYJqWFWR+VldSepm2WImNXSOIJQum
s37ng6Dsld5W/8kKhY24isB1PALEVwQaCH0XRU90caUcbqhzqgAR7BzDuPkDfhVuvm+t2u8ENsyc
FdJ/OmL/UZ+V/ElweSRGGHapgUnlckiBT9/5FaeTzMy+6p3ZruSyIXjzCIICHDOBdpjBA4/kpH3o
ug7wFbPMnra5LtGVULFkd+JYUgvix+r3yvstSAl0zeQv3DERtpr10EtTR5NMTNydABWMBfPGm5Nd
Qs1MPEZrlVS6k99Hsn8ssYOZwKMg7Cpv1yYc50Auhqip8Ca7NVRrPFZKKMR2DG/59il1ww4tMlXk
DADg3+/6Y1AIL0EOGzbcFQR3MWb3K1sm0DUinG/62WB/Lhfz8Lzd73APldVGY52io1afzZVThW0x
Cm125x7tAv2BpjpYXxTFXvLXeTYLkoI5LOeXZo2V8espX4WiC+gEIDBUpRUQzyqVqhjOajtzXyvB
+LOyr9toJZlezdYBzxBWxTkysGU8xrcSphCtT4j0p4uh0wv65jsuNmPq833WS/2FJpyCYipNjHeN
1pFS3upwpc46G/Lu++0woRP7aX2y/q+ifOvLaL3tUzFWU86QjpbmKdtZI7VZUSfRf4yr+KkgtbsJ
uwf3TcbNRbhvq97W7UKibNFWG8o3rw3gvkV19amawZGIKZTlhhWkaJ0zWbe6Ny3O6MP8XDFLncHu
MFcwqhR2cMIzDmXOA/NuWFsrdSXbP2z4gSq+pLytL6POz7FLaFxAucCATy1GF7VPj8CPMhDrxmrw
Ag2MuUkkpEPq1yS85KnmoHtVKBjtB34A5j+/4PCqBC6xxGEltlcVGp/TCMLZuqBgOqI21+yzwyow
R7XmzOwgc0vJxHQSvz863sqz76SJJBZ0gzG+sVn5VgxAiIWVuP3aPLIznoatonj+tpGIjQE6Lspe
lXQsS+7zE6WH7S4oZ5u/tr4Yeg39mRzIoOTpBuQCQ/L+PB5X0pKhkcDpIlUzXazKKiqW26HJ6DNZ
t+YP48dQ51mUbqCkDm8ay0pauo1L7rQgVqKh8lSK4ZwUmh4JVlsQgpcOSoDwxNrwo/XwFsWBBROw
vNXZEZWCI3yholPOyntZN8677zkfRTS4+jrofJdobZk5Fsrei6GtwqfEdiWjdu0iWS/oCQOoPa+I
oYqKb1fuaDEIMAh0g4TJPzjoToLQGW+aM6YgEWwqvzNxY9t3AXGoucMVY+mB5G8Tze28YLaajLMI
A3qw3i2iUZxb8QZ049eAEQfJ3ci5wuzh9Qzk7HsoGKPjfIEFslb8ahrdFrNfoQg6UouXp2CEbZew
omlQhJyRkYfUidX+U8DzF/1L2pa7VQK9bNFSqeXguidC9S6M2dLJIeMKm4YtmbtDteuxhuLLLmRR
ar7DfxqRJ4kRGHOr25FGcWUVCwlQIdfdYcnMh2HUV5Nwl6L0Eta5MDn9E+lxW8SLaINJZGr+gYIN
CTRdPtEQo+x8wT+luOsmtkkgc2HiDYPoFORg5rpjvyinXg4Y2ieoUqhEOI5QwVI5m1M6+JkF5WxM
m8cUkmAH0+ZHqp5lytWl/a93nws83yneUzj2sC1nwMwdqIlvtB5gvURhWsV7Q6k15C8Tycm/fly2
Bu7IlJg3MiDPQKJB/vFB8b0Uj+mqUs0VputbS7jh/4ixnbjJnAhgxmtsfOnYnBD4u9zozqKcPE3a
CZyII7FFQTwQoFF9G3v/Y4MZJGuSB3cBNtVgVJ8Xn2GpK3a5gRJxFkEBPiexcRydX9Zib3odON3j
M901wqWkJHHlHjk9boFMOUYYoiiYrzMeYOIXm9DKW3IcY4DNhwt474QZN46ZpgfgD8atJ7er8x9O
gTf/vQhsUUMJVdovp0nX8e12TRcj5YvMrMEgun7hMWtZP1P+4aHLt6OOQSYwZu81sj/RdOpVUdKl
M2CKkWZCt22jsuQ5aLkQoF4LYBSCwrG6x0lZF+asTdRs9W+l6NiQhnRIAyT8bBu+cOqlHAhXe7xu
ikYj9RBvo0Ck2m1FJH7ERTBkeADVCudNVjofU5Jmkg5oMo+WC69dGVUXuhFXsjY6+NIng8cCMuQQ
oQGvGK80NeXRl+prPd03KgI5MG80RNf3CawqMJTyDDD8qQgB5pAEeT41UZnae3vn1ztgp5q9OBBn
aBgUxHvUn8Jhh2BpLk/FJHPkmaRTyQNBW3z+kMMhZma9dj0Zoddw0ywn6qzomcqznMwQCnIy9SZu
cY1n513fahw3TdYDb6vfYi+EP04Ukp6dGbbW+8INSw7LzcsvfWNnJqt0jTNNhAJgaH+YK2sypyzg
whXac9leLdDdLDv7AMG2SUEfo31Y/dOE/3OO5PkugKwkAyHQipnCwL2UE/sjNgbDI1iL10E0MkXR
IAeMTGxQSNH4W/U4tlXK2Ko05IKc6Yg8gHYd/Jjxjwx8B1tbC4A+HKSr4XUri+h9j9JWZGojjqPg
DaYlFck+X1t+vaqPcTcRUEI56FDOT8Pus8x7vUr0hIIZquELlZFyCUCKCrMPKP0RLT/tg4PU28Wp
D2IzghWWK2vbgpQTRiA2q8F8tQarnEjLzuKSY7L9pEjBXHds54FRY7AUPmvDcqNU7A35BsIzXS61
RCsrH59d1M/XPtZvtjHOhVckKBp4DJuI5hT1ooG504i7TgnGcp8AAXmxk6hXDcEJr3B1o31GUOjs
gFPrl4OMvp/Kh6qhKyJeNDXNsBiakLYpUpQQkdlEH/Q64Dk6rZljl96aYEJ311RXzLwhfrqbCzLk
O6MAEP+/vs35s8OWz8tTFAkDqn+7/4tVcTsyF8IX6KZMzH/R9xa5n2+b9PcMREw0SD14TfK+glXE
a4b8uDOgILGvBxRoa9SyToJRQC9WKDQs9WvNqrl7/CIBI66ZP3GLLwPIaoS0AGjmu0teOcYus66s
xQHal3M5Qly/2cOyf6nDjj+vN//qNv/Qv8qiWIahOo8bjBhurxxhHTW1DXUIh3R2EOJMbwWM5obd
zHOK1BHSjFzqipDKIliQ4RpyQ7/8D3LbyTr3f7hyMCftxmHp31eDX/Vc6ldJ18I0cFIR6Essgjrc
uvEbLVBgegWJH+SplrfrapIMLymDmFxZueqlNnn2Qn7Ty/IbqoRPUy9pyheIVfikYpNcNGmKzTW2
J5b/BilzvboqrY59qR+P2RFE/1UfjupsbzrZb07U3Pv5suDbs2BKBYRwf6LJKa84CcE9C+n8h1Pi
20uY2Y//LzlV/45D5rrp8WKP+/JHQ5vXa/YLSB47oXc18ylXEPzRyHwE8bjDjVmgecoa7h874rdS
dQHy3lwK5UZwHW5dPzpxe3HMK2qrGbIVgOhsHL9M++5c6gNzvGEddIxCkuvu/hQhOh4v1TGZzSRl
dtcrndWM0atpeBEkG87p3yLmE89X45anXe0dobUapGMTEBnF3IEFiYolqYoVYeA1qqbhse4HCwrQ
JtTsgpABZhMwYpjQH8myWQAAafysajQiFEdMfzlC3HYdSoZ01bhO8pwu3LgViU+LLYpXlJrEVc1o
hjPAPDZvZpJvOU+1wsybufK+od38kmImZSYzeoPlXKG3Es12vgURJLyLrWmulL/3vjtZ2ThMnMQ3
1HcTNRulq9OEyRvGG1KLi3lc3VV6SRE/KVXQhWKsCenZSyZP6gGhnv8wU5Fl5jMOBq8+OVsmGgTG
LCF20B+4arY3UbC9+pabYHWVLQ7B/oOebQmfEeyqoGqDRM+cwWlhRIMM42SGepIBwfd6NcxHXpPQ
4tYlN2jI1HkoMDkgvH87uG4McVCtIP3LOVLYUG68CM0ejM2KR/Cr+8kpAUA5lUkNk5nvsyCzv//y
kOdL2I6FGaAlu/Zn5Sh6xCo9s7d0iiylGzKjHKnXBS8tn/dXW513akgtVmzaLOy3GPb55GQVGt9x
q1dlQ1Ohoha/0ggjnzcxA5wn1of+58TR4tEEmcDnxHjEl3I74YupkGD52uqXRLGcIynmMb91qvrX
0FF/pxBVPlwEycaxUk8OabxXJOvG6UG1Ap3dHitqy4UGHtOZdkIzqGk5hwekMdmOOsjXakwguROa
cROPRHH4a0Yk03PaOjkFfemci5BoIMO5kKr2RthXXIgexU/b2nkdoOnz8RBMkjSMsqKXGLhkUMSe
SzZkgC6G74pKNd3p/szLmdM5FwdMM86eBLsAsERLhbbg/qTN8/rozTMk21uVU3AZg/FAfeMFKVw4
z75A93Yqbb4C56Sh07LvjQBj1eVcnIMmf30qaW89gvp6pflrTt0RjCkR1X+o//8cS5Zcj816Mx/5
YTwR2KWbXgWwJFwXxHIhxg8kn0bv0PNVWcNjIQ8ugO/2Gcel5DfWhOaQ0sSgopD1x16WMSjJEtib
LM1Stz1BAdZ6GoREEfFQ6qvnaQhJmvmE4oVjJK4A2xtfbKFZSaQmjoU2C+5yhfjt+rJ8HAjuJuvU
3LgTiKb2Q50CJo5fw3lXVxfX3pEaJmC71gj6zs0SJeunJWN9vYFN8Yi3moZsWFYedqogB/PcxE3w
X7TUpKpISj9wQD/furJUSi+rALCddUa6s5wwGuWRsneNxheK9p4QsPnHae8qArvcBHoBx8DOzGO/
4G1ujo22Z9AkOsS6r5loivSSu1psJrqIMrhZBOUhHDH1MKpoQsft0MqJyOkmybpMIVKk9XQeFfL0
4TDyqTQ2Yce8sIe8PT4mmVJPMTU7FDXWck06dtMvA9Sv+VonIl2qgiU8hAd4Yy9ZxgMYHIRRsobq
mbv0PCovQAcroL/voJVYPbsZdJfw5+v/49GyI467hMz3shwEoJ7utaoKEQDCoJULeiWAz4TYmQgc
eWwr9NtEXSz2cA48Z4vNr/IPMDsc3TyoIr5CNnIKKyQwGDx5Ump2eXjeR7HOhXRjSauB5VqBsNKK
N6op/eaGD1ijRUR0S6+4ZeZ1zoz7lwGPAXVyo3qtDF2ciQyLUv3teHy6Q1MAWNxrWIerpJ9agPLl
UE2RqYGMRBV9dcHz4ss+/e9x7csOEBUBmUIJ6Uf4G683jXjw7nH8pRI4dhCJtfPE3/SQykiOiS5R
jZmnoHhur54/Si74BevFdlav+peZumRfx/Q4vfhJeU/vOsBuyI2AI41U1qHokTsBdPxRC/i8z2q2
ICunvfVlzplFBS3wMhT7Qt7C1DehVGlPee+DGxy6S+ivDekjNuK6kEll5TQRhceBHbs2nUa0LZP4
ogdSrTcFV2QTzbOOimRDgMtlAupvQFKMHwi8Vq5UWgREJf4xedCA+F78tAKVKOJAfYoSKuJMiZ5c
1QMAgUz9mplj4jIWt/Y6bYaOhuesmLNEBQVFT83qdd4+ZXQVB40tVOP702CVMBuzGYC0zbgLJQAP
KzlWtpMlPKK2mjyA/FEx9tfXH23JFk/5Jhhq3N5ZPtsBwUAU8u8/AP23rJ7zK74N+QlIjm2EUabz
wRoWaYGzfWj3fhxgiMYpM1KZwAwh3jqQJt0wT3kXiz92sUzNkVl+aCc4kAWVM/7NSDI+fU8I1dfj
zNk2DQ/21aEQaQWIlOEEQJmz7Rs8PKjY69iuSTIluWMYHW/BRVnThJRSibdo1pE93picpuDO/jyh
G9FKpU1WtubEulVAq9g2zq2LYjbKt4/KGyssi9wKsh0txMAy4bb/StPtTIoUui5dsJWZ4CEbf7R5
ClFkBM5dpkIChKQL72EgBOUejy8qfpf7VdxNaQXQr5VBLIE7fCW73oqmCKRNJw3hve6B971Dbkq8
nf5FpvgPC7/b3KlMtgD6f+tU+wACTd95nz1GXwF+taR5dkDsR56+/6rkNbmswbp0ec8XAVOK2sHu
BfJX71r9gEKonwAayOcUf7OrM3zijegCqN3AQ2+8sDbpdIKFutlRM76eZqJ00gZmZ7n0yDC8N3k3
mVdJTcR1kgV8WaetesAfCveDbflKl7gyCNzitfKmBHzCTG+JRuvSobQXEuL3isKR+9qFs5o+MqIC
hBKZVCmxXoHZMyrjZh3L1nyEjgQdRuQhfM5LHZc0B2cG4Q2M24eXkvSo7T7D+kumJi2VD1XrCsGO
S2KkjM7/yL2mXqRgYUpAdupoT2zhQRUiUrb/g0+WWLM7Vn7PdvZi35nZf/LysfRIEq6yoFRde9eH
hRKNeVeKQ6G8qUT0bX49wYgwFD6s3WbJDyyLA5K6zvBIZ2WfVYvQhPrgxM5S75BUfqzVM9Hp0/qa
8m0j1QExO2TY8Khio1oar/zTJn7XB7HSPTIHluBtKC4YvsPAIzZC5X3LuW0gflt3D2pocAAiRjCA
39uuPtBm6d2OhRgc+5VVqCmHMvHoc+WamkICAmQxF2q7BHchyKMGgSnu7LShg1iygm5/QYKwnW6B
jxbP/0Fcl00YklQCHjffkRQleLqQLShhWqR/f6G3rqeFOCIvEAilOaafFqxs4dbxWPRBlDiMlCeW
9rj+6uy+Sp/4IBic/nG/jGo2lIbUKYmv/U5JrrddxBpWnsam59R2Qi9YTF18/fiViWJd7tu0mHYb
HP3g1XYCtLIDghurS2owTsQblDUzesiuOqzaCaRuOWdU8DRascOo2vvz7YcQny+tbxjw3wnCaCVn
u6whgeo4i0egxDH3YmD2Ksy6r2OgyE2wU0M5f66G5rZlHmHMZFe0lPI7T/P8i4MkQfsxojgqx/Tm
AXRrO6mbv2Po2gMmbAbq2IDjjd7PrH+cTaJoIJTQSx+isEgyUGo5cMCMMEq2/m486egWJqZrWJj0
i9W024tMzOFPaQE8c0uDHGcw5BAyb1QxaHmsHbTKebVHvNkQbt+mnLdbAVmjPuoAWUgtc/0J7h24
4neE9eMHO7s6xBfjHfxfyRCcMXtpwlN2xDVUgMp1IXFGsr8svxtPzFQ39g7vFJtiADeJRRW7gTci
3Uqau8AgXrT4z6Oo78fnxTUAcOLX6GzDCuhN4j6PGVBXBlrbJxxuvgUnU0HTmyOnB1mJ/B3S6p39
vwiMVPtO3sjSWWpnKlsRnDiQUsmMS6gD1f4+fx+P7A6QdwxMD9bVC4B65B/7U8dVjhFWsHaSGhdn
263Mj9b5JNQad1GonBvB8ad3Nwi6i+WGXE28asRkjFkYTzWRUJUjSwudV0I09MoT0Fx8POwDDv83
nPHDHPblhYxuui5h7XKOgG2v6yUlyG0p1YyY6LNKrGm60yFL3Jq6Ym5FmUtMdz2XZwDrF0YpB+tx
wBt58LzBmUl1l0TTn2n5wzhzIlJC/pSUXOvTViLRsK2P9bbqWrs2eP3r9gS5QdhQpiUzepe35Cal
6PXak8JSlXWkJj1DeksvmO8m2UvPgFM0YupbcDv1jO0uaQaAbEbBPr1ooX3vOqZhnklX4XxTl7Wq
H6O40Ksuwo1AZxqFDtjCtX0o6RlBO3D26PRLYZB3EuJwobh7qYeGrNQQNG+8UqqK9UnxCajJeeda
6JO9dLLqg2Ia6nPyVj0zTJxBdAXQc+/xz1NJaheaq9M2dYkyj0Gbdlog3nnlhLVQbOxMSjm3ysp8
GIdU6iOff++b+wc72qTojT5lakR+j42TAXXG96gtXH4TG4dqKlvsgBeX5aJXVK6dufEf8//UB3Er
WzmuuFhOG0zZVfDizVF3XTv/WMRCMfYls8kDsBo3Hp5saF7tzqRHMw1eLUlWaabqsniLfSiwKMqw
kMpqkzETGLCSHut+cr4zgvT/2cDPCv0JJgg/T1wd2K8EtKxOxzykuj81Xl89Id1fcbyWm0Jvb923
Mda7Zaed8KUy9GmpPShOW3S+M2dim+GdVcZmlw7M4N9V9mP5F/U+l0XCTW9hTnxHzfHw3cMdO4r6
iSfmYn0d15tQ+bIJ5uviebKRS4T44gJypM9QDD197iSsRc7Td/hZSf0moZmXocTojfwA0LRe//Ny
Z3mn9FggSmdSQOm6EDvcetc12sfnuib9+r3PJQxr/8hmNGrHOk8vilUvECzYg1tx2D4p6vnTS17Q
0HzxYy9wnZRBelP2/e/lWUpHHU3VHHLlZg9XWHetMMeX3PX8GNvgxo9qZYWkHRWaTBnjiVoNcqv2
GSFTxKjAzUrwrSRd8sImR/dk8dB0Otrh/Q3KlCu3iWK/w7YA+yUxVnrqy/ZRPx9412nEhpIaSswF
4ag8vWXGWnepbjb5iFWfQIy+g01EO+kLQwPYJdJTcs1yio3zNBoU0ZX2MbgBEbvQLH0qybO4/dRZ
EtkxxmtBgjeI2ayKmRQ3TiFFN+KuZ/omjYRE7c5F43WMf0b5VHZTR55VKQZluiaOEZrhC+uy8psr
BxdSU4Y6B6vGL2XiC5JMA7eAwdk3Dyuz83UOfXJPTh6Q0Re9qkolpp02T//VJ2b9YNOC8oztpc0V
1eLT9fB+JtwyLx7wJPKJ2qZZpzJOabynEMP3ks6by79OGjq7rICj1hcljoHnmpxzkQC7iILIYSEx
I9CzgMZ5mXWfJB9drVAxslBfQpWIJgShtPPwIpC702CNPHdGOXWrlhtXg6TWLFY9H1qDNZh2BvK5
FlwsnGjbhArNH/9Fmw+FpWN595HFXbc94s+re9nWWrmDroJLleuvdslUIyU7opUdDPfuHihWw3U1
UowH7rs1JCRJg9LnfLVM09WHwpr1gOFdpZqy+pkvCHII2hFPSp8Y9AsqchDJrvUSKOBOijX7cfWk
9vMj1gcDOj4UH55hsChPvG6BGK3L4Uljxu+y52+5ndeeEVeqsepS+mfnyv1zpEHoaCvsFxf7LQgO
xYv1VsTbdJgQW9gPb0nHkRSneP6tN2zWSgRHrMrl/kxM8VoOrCQqG2ia9oxGXGaRfr4/QDu33LU1
wMa+wz7rWiS74Jya6J0QdHb+ifMgLuy2/JVzkrz2pQpl9O9PhuROTEtWzBaazqsooUUtB1z1tmyA
u1p9lr/ur8We/AEvSEjN2y3EWndkLJ27zM8o2anDSBWOrlQm2G/C7fPSQ9TTD1MEAfuejt8HC6lw
Gc6UoAwHDTa95IGV+0jGkOUR6B9DWU2dP66/FdwK7SKv68GC2DdS6hfPw3/OjFnO4v+EsBa0Yheg
68FTSOUtz1oexzLRBC6i9gmADRBY9vz/rNQ6C39WDJNOxB5T786oVNTwsbVEFDsvdgQ6ZQMbBNkf
ct6E0vUSOBfjg2EjrwGhzT4EizyPTdMsTOvCL/k6ftNur2MzzNIW1qPj8JGskElzmmWCfhc8fMPg
quq62B1d+wehR8WMNCSoXIZj7ryzdUXOm5mLzZt8GGLBNxG7YscWCJ8LkuwIsLnq472s1jbd69xJ
390Idr9AXdqwcU6mCgq7+8bGPBCmaqi/yRaiUe7jCA+dAu/PQhbziW1l2gCg9JGSsa1QCsSUfk/w
cH0n69fQuaE8GGSfKTkXLNsAlvmaJ0Eo4yJTSQHkBZaJ6Uwj3DY0MtTArCm7rdc5mW6qMVdEAh1B
IzUruzVA4jpa6p5TNWYwVp04h4oj8JnzyklKgRamUhL2FFa1oGVc00929X58mMinpCTV3Yba+qVZ
XslquLM+M6dus+frSMY8pHX4OxDNdqgD+VEnyf9cAlmtXpKvIWojAtQpLF+P/kEkq7rF4YP7WHwr
xtWaAkNjDlxeh7TGUCz5x/pLQ8WipDSD6afO0Qfw2O2wnMv5WcWlvZKie4fko1NiraRLQ0H8sII9
BYShJ9QavCHSYmxHDxqiDqa6c4AWgYCMdF27lrvHQq8A870dQxN3RPP0L+ue3SE60EWKu0p8VNfB
KXOR7bOft/fdTYdd9EttxRrm/WMd7lhcCDoLexLZ0V4rvWLpyQkQdVXxrYmB1dDH2clg/JAVLbyK
OlOWHu7PVgB4pzk5a87PA4Dmf+AA9UmQJ0GYmzvBBp68at3YDBTj/aQfVf6KMyCw8ZrIHQ/Ai5XQ
vHKvUHPzEfj7TMkETpKrjf5y7YeJt3RhvA6WxYuUkN7bi5BWoGOxgZZDF8PHs7FlydRiOYuP/GyP
bmoq1ySt8jd1OqXjAvNDPAwpZorQvqSbqhlGLlu1vi4kPEL8rY302qeMKPw68rgLf12LJ1Ae6B/O
jCOcO9pYP/o2Cf4U8N4g/vkhvvBOkehhSI+6wMpgnPvsz28/AqukZ0+EfgEaku8p2pp9UYUcjWw0
cazX3alm5GXi2+bpQN3GtGphdHDCtv9XIpHfQfTZm7J+DJ7KsU9HXt/lFrDRvjthDyhiuh/0wrN5
RPJ1+uKuz0pMiuElKh7snS+pZX4yFLRlKSbGHDtDSGi4QxYI8hU4RkJD3fN1mwrnrLY2staaAYmo
rjHcUnlW/wT3Srv4U8ZjhhDY9kNIwOnFkbk/JotkFNAgfV5c/bNJfFH61fzrDrm+g9E6AohE/H91
ZuvqziSC3Et2q2tcYgFFp7yPPGBRy9WL8QwtY6oMOso1/LFWV2AAeqqrE35+QXws1Ws8EEHAPNgr
n5rkqGXXVIuJTn1wDT7GqUy+UKPURFGkhYCM+6CTPKXM++0GpHQT8WG50L24h+S9bcXNEm0vUiq1
mB9D66ShYpECwubaa5XFrRF+VZPLCksG4CGcDuCMjrAoEq/t5G1oXitnZsSSqtwyf5hb0P7ZkUfY
clQ29E4TxDYLJvZOcKbJ0YqeZsarEwW3zplfYMp0L6pDZ46dxKDt5N1/Zm/zCpECx71fkfQAYDJ5
7wnJzSUQ+lzSWEPLqkoNmbXDgF5ZmnIsL7mr+RbzyzCFfa98UTyLjR20M66zZUVRxBiJbdj0ZB+f
Vvlb5Ty9A3UFUFYvrRTIIfiUXgDbJ3utFYXou4QW4gVyXXiO4CE/Ydx3NLvRI8YJBaMcx/hIWbAS
jpQp0hRn71zqYD+7HrymvYF9+kVmRO25c+lk+tfrTUWtptyWWkP9jlaJ7Da98ENSYK16g0pYsfI8
uDjcNKoYgHG+GpOe0ao285RwRD7xyTPLpIGZ2ycqG3qtyZLdcjaSSzcSPhgddpDE0OYzzNaIUmg9
sED/1y4Dbeo8jTrQmLJ7pUsnB36WsJ9gdiuZaArR/rup6ZRxKqwKlBYoAHoMw4sdsiOHE4Z8Ba8s
QiQCv/dFrqC6VqEymFQifcAXW7lh22syR7AnFzH3r/EB1XUcYxVvcrYZsbP/BrQiWdbzTL9WMEhv
iIXTfNUkGt28ZEXAazZrEphGDr9QpvuX+9KKvkKgYV6ckZ1vehMUobQX4ki7VNqYE5lki+l6YZBw
Qzn6WrXMu/1y4MhGqBKqRf6IkseJWEMTXsazZ6pueUSAOaD1U57iTzHAv30LAf65kx/CjAJhcdPS
j+8U/4acDapAxUZdpp2XNpof7Wjrng1GoofE8BcwQcZOmU3fEJ5rGea41sj6IBEFPeAmCGW48GhB
jjgqQzeUylNqkt2XX0D+aZQPWCtdX3S8b+/Bn56o0YQK0VfUIVrEDvOAawnOHO+xEnMdgwe4a+Kt
KWKgx2ELOusX1ERPngIgE9TnRmw2JHpMWBM1xaW9l2LAVr7j+X1gRlzuI0xOqVOLUciF6Ss7psnu
9C3iMFO/28pn6tkhYpYpwWptM+Hxv6F5i9Aj36nMLOsE2joOfI9L5fnYKJT4vN1PJcKezWPFuoNV
xaRJMGhi1pbut2wP+Npc0gmMNatVVoWwT5anJTaft/Olhc4HK24WuttAt/zvgzmQQclszOk3/NFi
y475cL58Um+0Sx/fan8oKfDHf0FderqwrNjLE6cguWv42sdpGxnYVLrbMWyGxoj/bm1J+3cNOeK0
abc3/mPwXJ3IVoPSQow25YE7X7Ho2hmD6hlH1qAxkG1nF2LUuAewMSY0Zrm6xQtO0h0hcPJcnhkM
qg81vlb/KktLHRHi0k09+FfNEX/q/VMKAoHrn0Ag795JrTAPwiiJHIV8TuBiFZqEFHDEkOWYfXUs
C0DVKXqFSH3rC9tRAzqJfFymsx5RDcfn5TjNI+1bGoRE9/JKnAI6TogKePjK7FjmZUDOsplBZRv9
Qu7QnHLpmFLja4P1wpUmcdG0p6LPKukKUA3w1ogz8y2qQ1tbzMYrEj3BN3Wj733VMHPpf4JuBNZ6
+KwqFn8l8HNrJ1uUo8P/1rsn0Q4Zf/QXgiUl4hUm8Hd4565/tTjdqk4rgxEIsLnK5J50nc/kf1Zd
pm6SBMdTD22BRANmqqiSnLdlhDj/r2P0ozkVy2ntXmrdgu6XzhjIXaFfwzjlesYjCk3eYZwGWEkt
4fdTXr0Se0CBWieEvrDZAFVch6xqU++vFQxePLok5K6TroH+qRnBkzAwvB53ONdImep3Nm8FGS0e
mWVmGuiFnnsfH3le4v1/LGYTWHij2Wdy3n/RJCG6oI6beFEvNNPARQ9dqQfNQn0mvNU7Qox52Tvx
iJHEJtaOUGXtybYndaBRkyPyteq9ACAf+joghTqh5Kcsa01qchiDCY+QxTJ85G/1w7tULuf59DPD
f6EXPQ12Q9TJXPl6c66dH93bad3bBHGXzxvLQKQ37SxxZUeM2NLjkcS/piu7oK6HDygzNxsKADAv
HSgZCM3MN85Avtpj3WgjBbD0d5ddFwXlC69iXbL5ZYnidwK2QXMtbmaIMmAQsIDCQgj4Wkms9Ldr
KL8Z4UhdrIfhltg+fDB8Ce2rIMwFFuo7wVgOMYIH/XHLnML6MB767JWuCz2Qf2mFD1JgY9TTUPLy
qOXH7Ttalg3Jl0Ziw/zCw921NpzrDEwa3hlSqP7evXWVdAt2sCt4lb30guPRSzhNqke80M+cFziX
d3sxI3guIlJ7PNU8evCCf7vdnuO5SBrG18HGHXCKPkao7ZJB5ThXFHWPggo0s2kRc/iqwNS79ybC
nyUD2gVmVNvQNI/U3EnMXPIYz2FdBSKvPbDetJ6VJX68RRyptdO65myFU4Fo/+JbvohagHeB7Li9
AmWnfn1F2IBGQXKYO7hDtr78s5Xf8LzDIw+GsNbd+r3BlZl2IjdxVaXfJ6m5RUNGd+m9xknGD7qx
bu2hTkVWaWhXbKB5TisKdrVTlp7qArua3DAyR28v8Mbqk2VdHFAM+V2mzCZLXpPQDSeSA4mqJzB5
6xAdcX/FWJc36O2VoZWPRMAFerrxzP1gC64sN7W8OkQxENO9upgz1nFuvSI/sXOiS1VmqlOWhLhQ
fuBP7UxX/bhcrn5DsJh8iTCpHkA8sm+s2fjhOtjk5QRBc6dFHQHX4//uP5NthXk6EOgiuWv66G0s
f2KtyVl2qO74jhcItQWcnkLFZvz6SssRrWvXKP/z3L34hgg4hQcPDGXQowhCuT46kt8H09z73Msn
riXXnDdH19TfqZ0cs7PEQV65aCFJ88llEfpfx7V3At8gAz0PpZjuzBLybmit26UE9nTZjbcT7Kly
nOqCsOytHM8TKXd0XFPn7rmI4mBOX1GCN+Ch2l8VvuqQQIXA2u5ATavb5GeAVX0SanXnjZL2ibaz
vB6BT/tFCkE785X7AE/GA5RvFhIT+ASNUVaJfPHVNU5efAnGIAIVz2kvhqsViMjCtpNfwrYycpPB
4P364KrIXOm/XcChEHBfzejTcWFnqKLsfR2ipkIms7E83QvNl6Mp45hnIW1/jiDRj0OoLw/svZym
zRS8SOs0vm9olJ2K0I/Mdh2as/fWYepvcCdWBqw7+V/aZVS3+5+syOoG9Wm0vXJR3KF4ecKuYivE
cSjpmgBHGh3ye3HTzFKErJDf2oqy8+6U1X/rOQUvKfzSLZo7Zn0O8upXbzSRi3dpsf9k/wQxfBkF
a3k+SjAroX742LozPS1smv/OmIcoALPFjjqKAfJ1cZtHuRChxnRZcQLwSBI0Ge0AHz4LK0iKj/6w
vdNR/GAXn9EafD4KTI3L9ASiNHAJPFYP1/RN6MIH3Bx81o/vFlQYSs+WjUS/2icgJkXMgIWXtOeH
/Ju2cSu8m3PT7Vk5H/OM0iSkMboy4MOv67YcwwOnQs6e8KyVZVUHuYHZvcNMIltjVAiqfIaZXRvx
C8s+4CiKNfrt9qo1FvurfYYLv0edFmM6HBtGCbbVfD5aJVVRKbuWBlWniI6zWNVljKr/5AHiA8//
UKZKPFlFx6jixAFG/7Xtq/s79dDgxtZc5Fie8EkZHgZJeBpJMqfFaqxjP6H0jQSvTlMBPH5tN6yy
DHLZLUgIK/MicBsaOTGK60fPiH6A0739BIwPmlt19luXciaqalaGCqnh2rhWDA1fgghXjxOwqWy3
lZXTOFmUn+xZdBOqGi4qin5RRj9WBbr7cpMVDeVvG27XeGwQXDa+4ADpggA3chc4oJpsqhuNOAPs
UnfB7onvVCD6OLEwQd6qkI/GcLXZ+JAFEF2WVWJ+ju20oXhrrCKChQQernm4wFrDZ7VRKwzhiJky
ZSZk6+ebeRP+ssuXezXi9Op1W9iFcecZr4wwXUqVDkqFak1D+dDSIerjepjdPUjxrXU08c4vcL9t
w/R51+w6vBjzp56g1+Zw58crZfBsYt/bAWOwFYfIOSCIxmHuHv2/D/geIYKUm/D26r1P4u2EkgyP
PGeT8WGRaJw/5nVqBPdsXJ/nzuoeM2ShXQVccpIyA0yCOcW7AnTIiDEh51R8dRFUREtQc7Yp8dB+
HMVbpx32eyYctvCiXgM8Ckexxkk96UG8YKKhCntYY6FYePjGJRcjlZxSsvFp9v3hmDRBCi1Ru3Q8
RhVmIFz3dNOsTwVkqXpEyfOOn5BvQlHkQxiphpnzfYujZdbLtF3xbz2fHQm72BDkt8ZdvctxI+yR
kUUCnA2OJjnZC3QuavjkHxcay5vCqijBNam92bWplxALug6p0tPMNjPuoh4yFJok4ZuPal4V49Lg
KxPKMz5NdbXNLBn2CA8zKoxZTnOWxs9pmW56CEtdI6zOBIjVv5Xv6C6/ZLKEJ5ZpvAVF9mPcEiT+
dbN9pVdzjaTURtVzTYtxzJXEhYXNloZkbQpM+58Os9UrTzwi40z3wXAs21FQOIrdDGvbXNtQTJox
BnE/o6glmI5w6qKsS1pmBrrNC4PekJT/JTFufMKW50nUmU1l+pWM+WjwVTppE3DkYl1y2U/QxMv4
ikGQRZ3ligrrceiKIQUezImzV0D+ffDFLMuBCU3aPgOKf6dDsKjSBYUqyvj8527a/8/epsmR5pOB
m/BdjK/uoBzORh36hNTtWbHosgCi0yVVSKf2oqjsidDTSuiSK14nb0UZrx9A6bhsJnxIcCvf4rt6
HdYCp3y/J4/ApozYJswo4WNqE/ujSMKV4ptbrXguOV0XM9/WqMH+R4UYhVnu6yyzEOj8bCtl4cE/
8xzB58ChqSz9DIO9HTuILZ4k/O5s7WGWAlYPpNHD+madpy5UfxEcz5ZilL3kaAy0zymRgGnKUpon
JXsmHcURD9owiut1AS4UpkT+aD+oqHe3JuZe7m69PDOiUo+9Ldq5PVGIxGVKGlEJdNUrrD4hkfOg
ZgpLkKFGHAhxsfJk4S9Lp3ldZYeRTBjQwY+mv7dzEiiYwZCpynywRAJdwhOZ7byNAnztZyWZNwCe
BYow4ZMaJW6lvBzfqsOr+yJ5qEDjx7nb1PE1VxMCUIfbJLdaNUx6E1W74QXBxHWd5WDLJKN5DCoB
GLb8XbqzFdbJv9TbjZnW+k6+QnUYn/rhUyQs6nZ70iYS4l6Ey8LWTsQhGpMdjh14Z9yixxpmPq5u
Fy+y6NsWgjK/0Wx7J5aKSZlwisTum7xOm74nLn946nuBBl68q/FiXLdZUL4E+sTx1QNRJX9N7beB
qMdSnC5ZQi/h61g/Fsc9roCqhBsAevnFYdutdnr4DbN8rtkMn9nDwZR0+SQkfugBgs+c0cmdClXK
BmjqFxCcxTzbEUomtK+/0JvSV7pQAStBjOu7uVP2/MXiTeyE7duxZpBZaD/nSXl0cNdZ+VcHRlq7
9Q6mL+uhUNHwYTAHPLt4duRIqLWhQu1td7NjtNeC9ztqfKkC9u+GjHvYpug+zs1EygMFC05BSchi
g9iMIlx7msxzyaXzDmXk7867zpism5fpxyhN8DWph9K4lQbUijpLYfwMBwqmUyzSFnYKmqhwidTy
C+JZ9eXbpEZfKL3lC3UUVxkNKtXc5A+lV3NqnsUGMADb+JYMhm2FRt0AQVaF7behlhu5xKVpWxdI
PUxSNo5EyYIkyUOsUeSV/fA7JdDQeWilRs6xovG3uHelvrcYwwWclczUL1LBNLrgN96QA0Rbvywj
q/RV5Oo58JWUO/lAtbzHxcuJ3Gnw1YFxCvZvvDhyOIKhylkjoNWu6iNcw2+Pvq3/7DziEWl0EdvV
SPOcJ9fMwTWrnTWhYOloOyXppcse6vFj/3yOe+o+HemNStYknHk7okC7cmPZVjVEo6hP0P6bn9a8
QPFcxpK3elVAQQuArYH9za3HSYurpzXLOpD/hczzUxfaDsZ2uFzW8lbXFKjkpfU1CcJbjtiJ6/Rw
mREgitWyNdaRW1f2dG94KqlImfynQ2sczyu7CMwSN15CzyUtv6MGAHQlF2/UwewO0JhZYfR/zMZH
FXkTW1uxgPqolPf57DfUq9RB5Z5Bmd2MeeuJDU+Q9iP49epY6wwQ+IyqjgLbx7i1GtK+t/XfYNsp
EfMw5zSpFAgE00/iT5pX6XUpz2XRWBS3lGXx2kthMhKNY+hpdY3YXsVT/hU475/ALSSqc62ZOdIq
0YZx104U8sL2DxX3OmtyDFOTbXkw8mwr1g4RSqpXzGInPsPcaCUCg0Svk9JmTmslZWiy9g6kl4hQ
uL+Rj6riV02pGwnOvflBCV65d5cbfRn45C8YhJMStE+6xfINgnECJdOSNCNEDw+ceAOcygSfHqlk
hUeiNycBsVIe0mwBrJH6LGFgjHptkprafgdOJErahS1A3NyObRgM7+kh4xjToN2nCWAPQyFCStcM
l6EN7Chvlh9+i+Hzm3Vd/E3pGiPsKMo9e0vxY9d6ccuAflBy06WUUxLa/Xa8fzwFVdESVNfV7nDe
3tIPKkk1s7XpyETzFFknOljxX5wZj8sVbGN2sE+J3k01gvjSQqm8M3onF9bzTUxC6qShW89VEPgq
DTN3k8CnOC4qweAZH2aRrviQwKy/pcF10xQ/UHU8H5EYJeGpY2tmfbiOvzyRtE1b2fwadjMqC59f
wN7eRsCvcVmaPr4k9/RXtuAD1TsqEEJxjNEuFTff+l1VjeOThGyt6uSEBmggvP5Sl12jVn/dCGBz
dT5V2rgbdVuc0cUtW2kmEVnliHAIAlwvfBurpk0opJtJYKj4Njm27Bg8hLEgFwcU45WdqxGjpOYD
gM7EdcWurXlMVjwTRQw7eG/2bVoH2Sc8f32rWFae6lOetYCZUPQY/q+LvMamx7PstV7sr0nnly8f
vLakxxBa3ZiQAuLO+rxbqbRnNDtFBORGopzkvUOJtNj23Yn2ukZn2TMFWOGNGWmAU8YXKAwnUrpT
ygVeXHlPMX/XgChSYy8kSkNSnuri3Vy8Q6hhyjsntvwlaLRgQxLun9iU++70smfN5NqB55j97++8
0O1G4dX4kpe2vC1OBrNMaKo1zqdU710qKzTvy4kq4KMS4MewrXxP89Ul8oWpRExSZD3NU5eTz2ct
UieiMl86KTd9oJTnbNYjedZXt1d2d7Ky23v6rpjdoja1mfUi3XjU+WnjawA6O6lwGSiMTE/wyyrb
sP0LQfzw0Qs/lu8IJzpraVy1UcU38rvG0O94pd3uHnyjeUi3YY5WrCjADgD/owOSFw+1GjdChHB8
ZYS1WPHWCf4cHDNT80LfzVgbQdut5oUyvXCauhVWBzoka+jPSQ4/ZhZiVozqPuiaAD+AjzBtwg8o
X7tirO1VpiFTdCUrdjsCNR0yW6acnoRlGl1/UDJkCXLt4l8fGFkz/9rBkx99lGERNenVqtMfnzmV
NNI79b5dhqew7UWFbr78nHtk64kWXSW0r14JeGslM9ZFOtbIq+wpgCziFswqnI8exRvdhaDaR6p2
ogTXwJwAMZcH7JiwfMM8DN4vTeH55YJjEcxkeIQ9GjQcxq9bMHkPIZd5fEVEZkwl9LwB//oyvIFo
6AYY/2EJ5NGCHrXv9wFeY+aP6Tord9WlxgnCq7PcSKZ7tFPbQmM9wlaU0v+Z0HBs+iP48Oz261nc
+Nwf/iPri9CIUmwFAprlLlcAUM4Oi4peNrSt6AJgrefqyOwmst1LW2Ua5xcjDMtPmNIIvd3yEp50
kYFedt5p0Io8R2Odv2FwYRrETO6hvQlIT6bBXLCGxL0Xwx56GQ0EBflM2OHOp2GIuX3bXErRcW0b
gBv4hskhnZGtoW3VtcE3Ons6lUvLVo8zaIxauey7bm04phOB61tw9hEuLuDIlNY8msWZP3medtZe
V9RjSItkF/3Utnhe9ud5ka5X7jethxvDP35cOIHHbpkjhClZ+w+L5j7op3mMZRqQ2DByoH8QQgV2
+5LRigf/rExsOGBu5NZAZaC2DLW9InxI4LtPgTWGWB5nAwlSxg5kqvfAh/gCGzoBejLBTIOT0czO
iGXmRlSeftbJHfujOFJ2n+lNuqCwWFd97YrQNZaHemm3r2ixZDyj1JaSZy7Jgh40rrZ/lmEGtEey
JzA94M5eYdUI9kxZt2VFtFBHGY5Tu5H5kdT0Ym4LzBs7WOjvbxY8AjtfNEMi0YoIyUYIWICWfAXc
aaw+zzwttYu3N5oulJaSHbqnZjgTw/apXEDReOJdrF4av87g6QUMDMaHeBA0V7jNp0l31mhD4PyQ
/qcJ90Y1VtLLCxR3h1RyPsHOjYeBwcpwshiNpaMJSwOM7P+jcXfniX3fSsRAdCs/zhKXqoT8/Jyv
ZxsiwzYq5w1HkUcfWxySlvS39i8Vr0ZR6JJ4wwSjV/L5egfy8lo+XPvyabYlIX1otNc0q4UofmTG
m+Ir6NiqRlz2MN1wpcNnuj+jdt3fBGDenLxIYkFGP4gk94schG0pVU2hZqlPM4lZfkhgP1AqV/fc
N/VUW52zHBSak4nSBciyeLAuWBVH+eEPUcHRNjo7E4iGHlaK1RVQCvd3K/9jWdUreZdqxNjEBG71
/cQZq0L1RBNBn+HrL/sFaRk+/tE9hsH/y5KwdCvVlwg+euLiagDXpkLwt+JGvJg0Jq5kNXsvmkOZ
7me7IEDCN/6DH/fV2egGmwH5IHYFGzUY0qmFIDqoHlsg9SaT1oEUddUUH//Ps/B1+uWNAFUTGzyu
IYTu+E03KRIkamaamw82+7PZ03Lr1eFg5Mh7EkqP5gi0sbu0eAXBSflpZLfU1WhXkoTj6dqlL8S0
axkzcBb0ZnKF/TsD3P69ePeCERDhe22Pbgu9Lb4gQ0tD7KxXBddppsXga5+FbIiDP+V5baHTyx16
LS/eAQZXyG6rjNQDHXUKt31Dczs5H/udLdDYibSn94fYh8rkLim49vOiImn7b48+tv6h27bUbnxk
IOJDiM+gjWzfrSDiOaVjU7r7l/diGQ9nIa7NIZeU1AlmtcORXmfVRsfFgPY6OGKiSX4mo+c+R6ZA
j1jpVc8e91XuJWTCFtZCvzbqgfLiwMImGuVCjeAZIf0gjK0fOThP+0N5bMFUXvN36rqWPQpPddeV
u9bkJNCuqFKtVJVWtVAt6aaivgZscsNmUEBv7F4B4RXNErV1laEIa4fG6Wz1mO+bN9KPdUiNp1Wp
lmWO8zMxhLizWx9GWn/mVrRpx1/okXMbQ+mjOpQCeOyjTMY3hyhX5Uc1yqHZWZ+Kbem9zWjXL313
BPWtKxKDDoi9HWGQWZHKRDRdPKb1QlxImwFXk217r2V0WJ++yfAPHWP7iI+Xn10MABBU0rUUlSaM
jHfsAsDR3Fn2HVPuqoetqaVumYykX78AoE3Bl6vFQQ+BWR8NpVot1tAhZQxqrvBm6FFuexu3CYal
5yqmCyw0Fa8hv8BwE3oS5OsiAqc2mi9puaPs4YGgIJvzFXIkqDY9fh3gdWqyXm5I0X5g55s2/gF6
lE0yzlU5TIdByLNJipcOG9s9Gsbula3VDokV0hvDtyYCTQRF6mhuTeIi/BU7qrf2NgNDi4SaztNp
X4jcLGFGBzuKgaIFfRY36F1bbh5tKjzLFetgCQvioQQrr6r0UPnSQe4bcwuPTzGVySrAkosTyK1J
uw2LVc/9jLPpTqKbqzh2////smLLaSaXHhjnMev333MrDW9rBBG/pMsGsA9YyqcNsKNqR2kuHI8j
WUNmTytIs4vdPiI4T0aR0BnEWwaKnpeJBGHR4jIP9OjIFHEkdY4ta7bZYXkutOPXLORey08bwMhj
VE96qBg8kA5pOoI0mxtMnDA9tf3/Ia0v/ibE14H8Q3lMv6lG3/0FnykHFFqZSBo+3r1Ut/NGE2DO
BHsZvbrpvCP+ewIqWx7S0cXMDgaCNIrSV2pscCM5DVLXWi7j0UnzPjV+gfys2q+YMRuW+7RnT+hJ
D5xfaqRG+bHkG+hs4icYT6QkVW8/2njpxz1Qi0LRaCAr4zrf+P8U6tkjuJrm/W9DsjVzYtZK3Cq3
MowlGfwQZjK5Fk2qY7v8gxgQLIB5VeEftwPawScdPJYDqL8BUzsjXoTCLOPdLkdjYQe3wau3ja/I
vlEZetT6wwGU4U8ShFYd9LhVn3dvnvJipVj7SCBrjcAkHmdd2hAuB0okJ6KPh2QJ/3UEdxGqNHxv
GesBtrST6vI3dSb4S/lwAyfc/KiXoRzTqWH5kKlNdweEUXZmnifyCWBhRQVYtVYllBOKutzC480u
MOVKEBZ87l0hvfQCZdTpt3LjdlprF0QzFZKvS3upGGveSLe3OZuhJEGGadviFzp7bvR1nZGhOMij
EVZiRbA8G4oqinDClbyjuStbwsaBuXSthqiUWTF/8I4tWycvGG1Xp3bWTAHzyXvtNFyaesj6Svkl
9IyNnQMFMBY0trgkZlUNt+F+Fg25m1jDXU755yY4cw698JRI/J2gHBkG5YrYjoReLVEOsO+jvv1R
cO/tE9VdodlZq5FVxfI5ITf4xVYw4QXq1lqOkA3wrVtoBUic/gm40jglJPCGgwYUYV1kRNH5Sohu
S1wwD9Wop3by+MwVBl3M96YK2unkyUfGA8LGAwPe6CJzdRJnDtRU9iy7oMSHCBxUHKzpAht4V9H2
eRdj6vePqzSpRfP9x8hcQ6XUxGA6sUwiioI4t6a1N5k911oCMS3MAWSdFgwAkP3VAyMP0q+wX4iL
ohUPFMik79pb2p2hRynbrwSRnEFJkguWQTJ2y+/1JN3xbK+NkUP83+375mfLhoRB6zvlT3be3NwN
EXbhVJXX0qBH54ARgbPQKLeYIgzpqlhimu4KC+8B4uxIxOPnKoaGsJ1ByOkvdoCDeQm8yLEKFy3o
YnIALvwa/e+GZNNqaSUduE03UD1jce9HdQSg5U+AFWC+Y41CVzjO9CotBJLqVoLSRtxeKV7nOeE5
gsVKhM8Tq/COp1VACFi1ttmkXZqGjjbKqvHpDHJI5NJTXxzpAl4v1hOKA2kSNTrDfHSY8zdY5v1s
pwu7YdA+sjmSUEAOkMEJXt1XO2iLaMypRTedbcwwiWkU+zC0cgNvnjjLdyYznmsFsNowc2RSGgaL
CvYQUIks8e3cnE0dSsA2jdmpMRxGHBWZJN+j6goc+t/EASLhta3A26vkIXdg9RtY5BSJJ4+pgfGq
37MnOr7ZcQck+Ds7xgVexc2YK2UBctJaHkEj0oAV4Lx8hQ17L4+vAQef4kqTph+GSf89FjQ4biD5
7PLbsP2TirLuHbxjRx9rS3I8WIpyoiWOC9z4eCG/0JmNwEV1D/cASEAueSzeR5irh8Ps+xoxJacs
KLPrcSp2wHu22hVFtA4LzRvOYZmf/LahlJwjyJeQsTjBgyceN771Hh52kDrPgXGoeGKCvSPxuhl3
RolEPN0Xn6kv5A5GeJszRKlltaBkPM96iz4Udohu0CB+DKBzKsUAx+2B8Qx7MBDAzGZyKvsONNSL
TZaCYkAWS3FsNl9So13XCQmftBhDdtDCShgmvRqfbthZivaTdUTA/oy+1rLbYY2degkceWJ6D1s7
Mj13KlEu6GvFgIFp156qdJ+cg/H4y+YfAsvPQ/rA6RCM+MMtuTD10bY5tXvyr5GHMfOcjfkK8GmL
TrvL0kIIrQasypcz5B7pylEeHvqCxVRIw8+gqpRiJQjqPZnSMWwCb3CZZh7jtP7C8UVcbJoRoFFR
JSJpZMA7GkULF5FDQ8GjDm8y3EyOFqX+6N5qN6UdnC1mMYG1hL7m12b+ZBFInw7fgSwJiKWubDU1
0RE0Nhgn1gUdZa00RSIuC4hXYlJnVfIpMlHbv8WmfUD4LyqhvIuZjTCCXeK6wLSAB/hJu5ivSkbA
E8ndczfGSXpJvT6VXifHv5Q+PH7oauvKWWr6s0w0yzj62xQVLYDyBuA54RuoY2VP1vFyvs4Ry0Il
kQJIi8eZCNHqgIbSIT75QS+cFc2jTKS+TzOg99IHLjvkz6mLMReRmZVhwOZebcNeFMnqkiFQu1XD
YbetYX8WXHU1gXyJ9vhcXfCz8apdHdaTYjCbwcx8tBhxT2knseW8vBdjObe9DSluR73wzzZPEgfM
DmS3Rmj6JacaNSPKKVvAhb8N/aysiOfgvH8wdzP8Gg2CniC4nMtrIFhqGljCok/KJU0Jyiq2exXU
NIxzYpUdrrjt8E/dQgycC+f7V1Pv/YE0O3N0IMiu7nhznv1Akp3bAxd92GuvGpjSKDQrcug0nM7J
qGJYVshx3QGAleZBTq9nGC30e0UUJ58QRMyltHTa8E9r3fMdRSXd0r/yhrbD8eQJsexukP8uGuKV
RR8rt8OCFQxv86Vyxd861Hb+HA3mbbVHPW6coV18VR2vQg8DIMLVvPZpsWNqPyTAGMtgbmQW5sqg
orazDZZLGtUDsdFtrz52Ds6OHCjCpWeXFcruZfmdbXtkW0bNdmI+UCJmwE/39oYAc87a4DUvz6cE
7jB+B0S02mPdDO9K66Gqlhq4l0WrJPIevvtXLKQWKPQ/tBSe03+2dtYZg7nR37xcZqAiQuaYlvzB
56WkAodQwbETbwKl/bthajmYQ4MBlgPsbTF9vreGMbEppo3+mjeoFGJqsfJNl2XbP+2HJGOc+CMy
+0XjoZfR9tmO4hHoyJjhiKQK30J/6kmjV3fpvctgkyCjL5ArhJQTCSO0Ic6NyzvQTPk8kE1E9WA8
36R+Z3Z1Ono/kl3NSBstgqAD80fNE0bX5PFc+zY2XzfuJFiQewHHZfY+Apj6b9qeLCcYWqbh8XmB
tjjMbkpaG4OS8caYe1D7eYUxVB5si848lwIdlPla0cEGB75MeEVhrJegW8vhUO6mK6H/LgQvVOIa
j/tYx9d4S53P3grmHI+cLLuMC3dwZmgekt/uLasNsQNDfrChdRrD47EUgbLOiAMagnX35Oh3/71T
1k6wxNnHeVzLkNId3Q9bU6aNsmHJpPTOr+B9gecvCjH6ROwkkOfX8ddf1ovxj0ZozwYS6Q1bq7hu
5c/zZD2ept1nEu0hakni4iUzEHuheQinQW7geGVAJAfijVerlTlspUz7rH7e6/wd4OydKKvcGcv3
IB1lfjC3rMWSNjupnw9L0nZSrxYa6hS2iUH950Q9eaHVJNItk1qPzlu38KZQuPpMT2U0KCNSPKKH
PC4JLjdU1c2MUWS3HsH7cJ65PLxr7U8cJaoQkW7faFH69LkqXomOF7EG4txleOgK3o7NZn8bfZkC
BNpZd5dLRK4f80sOb1QTFRjaO3ucGGy1Xuy+27d8eSwBzgtlqby01MBjG0/Zx11rzpCs3IFsxXyz
r1L7LukCn1k2ciHe/vgWd8WumYs1veFoc6GpYhbzAV3bTCM41eKTjXGlFk0/Hgyn0o0wI3UDLBZV
bjW+xYGXnJsLjYnW8Df6H3gmqbEMC98iO8lis4UBJRsdDN+Pv8bDXpFR+JpJMRR3kqo+0PJpGX7y
ZXUle/ceW6S0pZ9h1JW8RyPDPJ91At6m7KbfHv2DfkjbNQntqhdpHRFUe1BYuBuKubTOBz34E51p
cJK5UikxOBGKcBgedVN/pJuLOrmtGleuwKT92z82Otk9Vvu1H/MsDpkD7e+5S1o6XXR+dMf6VruY
O1caJREyMY4LTkUYx7muNf+4g0xZgz5iWuI4mVi/0LTKBi4SR2bnpDnuLXeq0cOgnu6R8Nh3jloK
v+3IXivi4x9Mge96BsrIQ7bTgJ3tnji9VefwsZW/+etEX7jj1ESdPmElfXzThOhKrISw1cYlrBwT
k6Ch2tNqB4QZvqgR2RzaP5XGV60kXeLyydEyT4pEec1ErIAVQum9mti/XmTrlSpPMw6vBptFWEFs
7PubOBZFBRzYDwPdHnKC6dCrYPHDjYVhTT2HyevNqCnn81NO1QbL/AjkLIVnxRUTlKzEasD7hm70
HUApD+vEl3v2TtJYpb/IVgfjrgHWh6Pbf37KKSqR0UrlU76Q92yz7mR8nAnTF+Jjvg4beHCDCmGD
yklSAmHA45HlA20iKEFLRNil7AUZ0LNbBvPN54d1zXsUFO0GChF0JWlVZwa9MjFIia6OuVnCyn23
+HmlRr8jaSBtcHJMCvaKxjgm0gUIwDrd4qbC+NninIRVUPolnWiabK1zGwSSZlWwIAY51JeyXf9r
RY7Nc2WV5BRgwWLR1lSPNUxe+F97uNlVIBgDLdh7YN6a3N50jmZn/Fa69nWgLMWX7cokQXy/RFKD
z4DxSYDH93Hb82Y4xny8Q+UtQJ5PT7qZ5ulF3LzY6LsOjCLVrUWDdQ5FjAVlAa6I37wt+UZqqXg4
AjgSafWfcrAct8loXfOfkNtlcYB3UUZJEk66UlBqX+OpVa1BG+kI/7FzafyX0iFs0l4tk5vhvV79
s48cQ9XxLF1C9s4qc4xjZvl/G552bA9806q1eHzshUwoHMiquJyRFmdqVwtxackyJYNcnJRtOSBS
vpGNEUmi0kIGwFxagzZJdrCOUJa6lyXtXHhng7+IFGRpZ8kl8PIYSBlJ9758jGBiOc5ScG5hR7dF
2ZsVQQ2u2KqpwE86A3hdPDcIbhBZpgPos6clju84vYimXzPh+/D0dn+eqrgQVWo6mwwGges8i505
FN1YzgrMyu/RLti1whsLiQf8jKLmDoim+qwnkWTGXdhxhsIulEwINbjHo3OtfNHHC+whHrpROXwS
vJPSUBWv4GPEPHnBZSfIB75xe8BpDm71PYWxXBRj1Uc7KS1TwQ+7CkGSemQ9RMjtEQCu5UpQHWLQ
cdcVNUZLJlrvDG91WXAOzxkWZFpdypCDs+6lEVzhwKhhEPhkwP4WhDSSmmy7WZmfqlBxw8/iwAL+
7F1iaBpCaabHygdX+dEsAID0P75gqCP/1cGySYv5HmUyY+ysR0T8la734/HQPePHlTOVSnpgHWvM
RA9FNjEosXYbdDaY/S3/5ab7knw15a5XSIWZu69zo8oVkDZNFiWyWlUwibLcWk1GEPz6hJRysCvh
465PR4fsigJxYDnKaEiVs2xGmYakB7pk7eobLQ5zx/oQRnzdFRfhBujgTUUrNUtMB3ddQoeOjnYN
JzCdrSJt5UuOzRJfqaMXVs2Gl5vfOIdYB5jr3GvtjGQUo1BjskBQnVFjOKNDz5EMFzVhx/BSEa19
n0VMN41k2ZfHNzBSTcU7Thh9DkDV1g4n3Q/qBsYhuY7jr2cXwfslFW4iJRVgtQCj0kGxx57DHJLa
//SZ8PGUv3U7m55y9ez9Jj1PyQOSWgbEtvNYYkqfaBjDo4ectB8DWX8bgYWV51ppo9d2d9Ah8P2M
GuOe7aWgY0laMb9lNuKMMQ5CUVegf/Gz4SsBjhLmNLopeA1JB5wHJp9+b8dHYTBRRFXVjz9G9IMi
fIZUhHjBWQBqkDS/O0sSWn3UD+DoLE8Ae3QV5/MFTym14gdVwqibTQ4oHQ3erX3Hlo0m8J8myRFR
s75WnDVDYyAr2Tsx3OUzh3+TyXLglRA1pBhedKZLGy8NobVLsMwHg9OcFejvLYhibPHJvmiv3fwM
wSmq+IQdO9JuHvD+FezjYbRFShSkIgoPrZ1wWoE4iSnPdOXxhZdBtjyQUYs0JBjIX/eclN2Ue56V
WxINKBGBY39Avb6SADf637Kiywxuuxp0VGusFUJWRsyOduwocrc1LPfz4/0o6lAQmZZBz87ww59I
YbDnDBAJZgXohz1CElNWJwLmSXc4sfnqUFZVfu7TaNyaMZuBsnAI6R3V3FCHNSVdWpQDwpSAE9Ue
dAxxOXhZxrpCdqjY/jQfbbMTHaYQ8moggHasdjLXrQJyMjAQmpnDrHZjYD5t//Lk048BkdsgxOEq
0+Lq/aQ+75PmKLAUlA7xWpl9nGiWPPbyRRvo7NpLIy/M5vQ+vb8zFACJoBZnQhV9tWgzoJsF9oYv
GObCuffEJaWsiI4Aht++mKDsefXzRMFjKgKYRlQsJ/ayiY9yIbCUxcZspmX4kr84xoJQ0q7K7YaU
Gy4IdH2RHcmebcxFkOvYDQCbU1qe08N3V4muaM12kBz9ZX85wOdIq3fbd/o5/U4XlMwnryfNurRg
b/xBMpko7J3EK33xrcTJXyPRmZv7OplKe02lBX9OISngCLYMXelX8xLzKCE131RaMHd7BGo/ST42
6HVXk+/DqYZJKc2Iu2YqL+gdHIoNO2/H8Gq5oMn7RcJtxGjjGYgigtL+S313kCvQih7bpUjcPuIs
OGAYsLhGwdMQKhTHgJRVFhQqpP8K1rgzr121kc99ZRm0oWuectSVRQnOW3+02sPtODf+TavpZ3D+
EJTWN4PHRHv+8DvQCTflqABTRas6YlmFW+LESlWAt3hmZxrT1xhpMO8N8bkHKuy3nzji9ktmsTjK
DDC/jM2Tyn8TIF6grJhatvUgeK02DxASaJf/3SIJKbKEuhM0e9WxaYfX/Udak0zCatsofKpovxgG
tWkUXU/PUDYiDDtjVI3rKkzhejDCIqBLBBG6bubs65DVEazRRcfGtrB+m+OTyMfGk90uuumwyLO/
yMqc/jk4WhE2faU551lxfhV22PtONfIq8EZyT75L2x4okHy/oMIgkcS01G05Xzwg6Aaxb+F1Px7I
3ovrda8HjocwbdZtqPK/APBwchJvZt2hWOXycPoft56EOHrwhY1c9iCAE4Kp1otD5z/+tgWlaGt7
JvkvRVucxbUGtwliiX7PK8/ScRxN7bHFPXv1BxoNEVIE7dpc/SLy5pWqi6gIlm8tn2AC+o1qMRAs
Nt7H8OfoqJJXpIfPwq5KvN/Hy1t9XBR7YS1DOzLrthwJk1/B69o0Qu6rMFKaItt6ueLNlVXZZL41
pnzzYN0vJR01/D15C5dFgJ1fSqjoRiENIAwRSQ9YEX7zKS14d0YS1pUE5dq2qsi6fz19HlXr3bPi
2tuwKkSENJEdqFGN19P4dvacc6k396CsSIXwg+HSF5OssemC7R1kgdiyfMcaf8EwlISdc1E9WCci
3XP1GOAJPjc93ClqonzeBZscCtIHjWz1H+0S9Ow6jNoVV5dMN6YP+m3OW7uTZythK973OnnD45EF
p6qwECJUAmgAfXgFlHBoKoAl2+UYWLFoZGQeZGQxMmDcu5Erb1vLRQWY9lKTp91jT77QSCLfk3bu
J1QErp7huYQzAix1M3yQFH6eVJP5lxGoR2J7ihulAl419OWdlXTyTYARGnwhZvyh9dF5MjuTBCw/
7OePh1W7zLf0JHX2SdctSTRybr9rCr/SA4CsdAYiGBjcQr9JVdQdpVgNyhZUyV0ehvNxEpLolz0t
vP9qkKbB34NJvQiAuHC3JgOzOkdKjC9KkLX1YEUn46SSBARP5BXkZS1gqZrl/Dj22qmLOCIRp/O/
GMKEtLUPOM9yLgF66bV2Hi0dU4nZvFMw/Rgp2ckea7mwBVjd7RTnmfj+G+HCJkrt658t29Zxnqi/
KHPu/JLBd8+IVDXaXjR0IzVXJbX5LsVlUMtcX2KeGhREUSlMHhvGaU9YHpXky7NfwafI42x4yDWs
rZxLDfBKFOcpLtQZTPaAJ8I37IydcOP80sTd6L2rbOkvos1U+0oKFn5Ce+RJUnRpf2kXhHd6KWM8
nsH4xekkv1laVXWllo3qSSEvOHqDLCVp+sBAp/yK2gIsNXviWMYjaNkaEdA0ijLxjk1/TgCziwrQ
tb9ILUzEXPw3ou0Xw/mmJu/D8BWQ1tka4zV9blmt2/O+6Og+et1FYE9rSyiC1dtsRrXzZ2qsPBDX
kmK6A5YIMBI0fQviQ5xicSmONVeRoQ0r0TiNwlM7j8qJKtfOYVnQ6RrIdrKoKQqM7czLLY4azETE
WYq1sQFfeMOY3yZwNKv45ycyIOyntT6m74s7L/lvrN5ONxsnt/JLZ+3BBsxGtEWyVpW0ZXAJnvti
bIMcdhiVAlRrTqcWG/4Voea3DJqWRkclkcBrNaYuG50phxYH/CTu5Dr5Mj8KA6oXWW62m5rtrXVH
RIW6XdQbyz9u4swd/pWzsHrsme560EuiMyUf6nZ6tZq3WuLYDPgdX0Lum/ooDjTkdE0nZWA9rKJv
qtNTzzKeL0SYK7V9agoJIaNYP57atiuEZwnKKm5/4F4zAiMttptClMmlrwaFNhCGOXqz8T3QXbIk
DUnfZuX8S/YxJr5fXsWAulRrxKrI7GLv+o1K13BOrHIpWT4j1W5ivH3L8OrpSXl+oiS3EORlyG+s
3R4lKdz71UQ/Lxq88VT1xjAcLQEziPcPV6w132+koWS9zhs8fTCGuUQx2+ZS0ZnaxY9hQ2ueRpjm
aQbpDr1WylbWlzeidnUg8+XLv14AhYvBVlHwZKis6heYplRaHqRN+5xXehPd/VvmcYZF4iHKK7Nb
SuGDiorcceITEu110zEDm2cIyNgf45HkxizYLp06VGn//2sTTNleELvZ+dWWzUZxUtHF5msVrMGq
sjCAv7eEznJ1yXCk0ZakGQy9zc9czvvgFCx3RRkSQf25sT8EeNzqZoxyWMl/pWpW3YfXlU5h/3gE
hZZrjgHDAQHDqP651GXBp2zJymOUExN7D9KnapftY1j6yBXR9ftWq8/Ve/ms/3a+0y1up7pSusU3
ALFhqd0K+z5DjiTTJ7HTIUqygl26zpG4974R7dOufpJrfUWk3BU/RyDTcYvU6qCjJ5RjIlBAl0Kp
Nz7Ak3x1pguHXdGGr6VN/O/Nx294SyappJxjrm+yRT95SUWEoRuno4n6TX+QsF8AgISQ4A139lCp
5OFW3aW06BuUZbNtD4PuSivVhu2tLiSmNHA9c5EaI7hIS/blOGB+cBGHaKYuTu1QKce9Pwz4+hon
eqFjeM9aJ4ypCanOWhPKjZwNCYUiNo7pHEWFqhufFyY5D29v9i7z5VILCv6kSZ/np4GkxjnEIVMA
pdB7dqqxi4Ge2m7JpZqohCWULeNJAvX+UwEktKCUfuLs36chzDTVZNMP32tFEu/5NfgOW6XPJ6yR
AV1DIWSAF3bHppgbAflnoHzqjbIA3csWKOMBIXXSoXKar3F1PQVP2/3hGbi5DGZk9l9Dh16wnGHs
ID7qcg+OFpbybcmq7puDZQq0jzQ9wWFN6ukyO2WInfUnPvoouGwAsevAMOwS+oO11N4sv1M2SLf3
w4QPvtZ1dAQtmaqBS2ngitRqWyhpM5cMEHBySdriDICxBG81r8DbXi7LPuIZoJb4+CNl/wU5Iw8v
1sAiurV+rbjBUz3nSqcCXpEUTudHn6HU35h8cjUR5q4YptsB73TPECZWQ0umfs9RzAXALyE5k1Ov
td72LajG6hMZj/QejH45v5zZOVgYawhdN3oOzrHEY2QKauTYlESernq1eyFfKrT/IVVncf9c7IeZ
Awms3IhYnpFd7zPL5gRgCrV+sFGiOQUrz7mdCJ/TLjlvfRGeGeCXE4H2IwJBbkgevuRgA2Tmyd+A
zkbPXWook01g6wfDO6Fp5QS1PuYJr2xGRsWK8E9KsTkGBEJ/R2aGx7aL7KFRxtki3wLIdoGOZW7R
seIvz/FF/0m4Rcnmcz1bWnjztJeIzK1xYK4YVZNRz6BFEckgHkdu3OoKlhwN0xLdUyWLolcgsOKr
OWybLsECGdaA1wpsFwOjLQMSQxFF5tc2f2Y2U/NwvzS6Rbjvf2m+zCboQwj3J+hDiL8txKL49kYH
YqZKJyw4l3IZvGEPjWWPMfKTtOLhbB6PkCSogq9+K9L7fl5aDhy1Wcx2qNpDDEjFQD4AYim08Uuy
eE8Ym29w4UjG7EwZbr2Az4n6hhbyxwK6eUc9jBrPqjKc+IqgMHjyGAS8V5bSWKlVx6IixnHK/xve
32esHJ6hKcSvLrnS9h3ZJtYnEKCRyRtBmFxgMDqZqlUxoePLN0R19kq3WrJBXMO0CgggK7W3/WTW
e31kwl48tjEwxLIlX+qxsjLwgmkOEADsMUbQvJ/0IfwOtEtB5f0eBWVT+dhp5uz2Yb/gPObAP0EO
TDX5rv/YXhBwKnUrM3lzw9sjGmHEE933acCn6urCOJOVRMObnhlbGxpMCJFpl+k365SVZiKK6Grq
lNm5UBRUXe4igc3hpUu2yJKtFqdoZaNXWBNAHTO/ulBUcEhxyFm5pZqDxqt9Gl7Jw4BSvpaLloTr
yedT8IuXgY9lwsXeWGkVkF0+ZBlNeFKQ+si6TN7H9K+Ti0EG6j+EG+egJEa5nTasTWs63oqS3tcK
yJuiNu0msHk4c0VDTI//BKeASoDyETmoEOCkxpI/vHik9tTj/QK7DqnnkDLzX8XHPe1e6Q2gOuIi
4arfRFecstqtmpYdScWpM4Jf9KVq/y84Xk8kWGIH8qEwTwQhXwjyCD29FgvHYuB1Tk7przUFE8Ax
1t7pKPtM7MfvhIsckMu1AjOaXfPr4zAT4ZF032XMjPNGdNBmCkA3KQQw20ESkgavAOgDI2wg1tsq
FFRt4S2teCY0I42y0L3caeifePQi6Vu/rj3VjxBeZ/l9QZkTCtwR/flEqifNp8DrfZh7gZMXa3ig
sEISoY3I+EgogS5Ds7PBMH5AtgDEIAqhC1bahtbSc2bTlJKc6a1qduOKubhFp4t+40dWzgEuQRFP
sGBpJwjH1H/dEg7SwImC24hIYBN+XE0YELabWqRyFbKFgIrCstCK8PxOT1p6A9EfLsfIQ1m6Lw2f
WkP+3K3e2kLpZRDYGOZf4onenPwuetlt89iXk3i5A4s6qv5oT0qyJv+Y55Ng2TLjvFweUX3uqvwi
2T4P3QPqMPznxiKxZqedOO46OgWV7t6LHoXB8ecPnqlJmXl77yiHWTa4iTI28xaOTv3RPnsTRKz8
pvbW8FIHUiZ5rtNm3HZVazmvQeqdZ6R9YnBO5fI=
`protect end_protected

