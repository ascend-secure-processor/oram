	parameter		NumValidBlock = 	1 << ORAML,
					Recursion = 		3;
	parameter		EnablePLB = 		1,
					PLBCapacity = 		1024;     // in bits
	parameter		PRFPosMap = 		0;
