

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Fs4xUNl4QGZ9/2RobM8vxTll5QHDd4qxr+8ow/53LgEfIeV5QsDleD+KQi2q/62p7J7eL2uJNefv
dOD7ngB+fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SZwKjWKyFswYO5fKG/x1o2qvmidu4iy8aPAJyBthZaWSvmPfeWLxnCjQUgycb74tc3rj5pxrkhII
S4UWVzvhAXCSwhYMKoaPmivnit8pTDFdRAf/kL17qSHRIM2B4rX+VdpfuuoOMTcGTt76ATGlNmYB
uBS+iEKt65dD2WdPoMw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rMdNON4xV4Ckw2bgGE2G/px0hqcMCLofeHarfz9xCdmHAQeiPFfC2RtPDB/Lsuefota0h7fibQ3r
ZJhuzws5jH3a2/k4BqZveDDMpPkjaMRcp2FgwF0EbLvfaLz/IMSSWcOzkZXNKtA6riF0w4saVT+Y
q8UTRkTYS3GnWIMh3g6gKDpG9jPBy+cvIZ1bFNHmPaDnE3vH0hkqmmd201q39ZOGWyb6JwrkHf6x
NW47NlVQEk1zy/46nBRFHuML6gmYOZjBpBsmyZgvDhsVZCB8P544qN5UySmf2vhC+Lq1226E6DLu
wct2X+qNckI74M/WZdW2bf+tx3ftiW7MtOORUw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fD6sx01U0ZLTwXq3gkdf2CXEwMGDnWrjcYTgPBd6ssVDotZ/2YMqTP0/AvuYbG+bEy0bk8I3Dp06
exmrg25nyh+k6eU77L/jaCVnNqhtxfOVf03MDfx1pIR6d+/Jkv0OXYOmka5MOXIyBAnGoiFcLHG8
qvJO/0bMeY0TGbHn924=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pqBVb1i2Ddny5KrWb+4O7laTu6ajYyHQNuBtEyj1HLcXLzsukFOpd8kj7kODzgxwQOOwsyJKVzTm
uadSD00Op/d2S9zYpOiXrPljl5lqOb/DkFfMWeL2ysi+L0e0lme94hJ2Cdk9sXYiWnvOCPi8oIHp
t25OcXfm19dCFYEaYUdH23S8tcXZ9RC2zxcLGKCxnn9wEp1DUJfAMZ3wxgfrbY2JAgzHcNg5Qxsb
qnQVGmRnCsbgU0edfwWC54Q+/1wnlqOf4N/x9NiGAt/7RJ3Yp6X66vB0btoKM8jVB+/TyQbp3g9v
X/gtmzeuRjO8bue9Eudatq+jYPQGDfFp0CVFsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5680)
`protect data_block
/YODsBmETxjYyuQSWvoHMKVjFy4Ec+PWIMh6gHaVGh3Ay07FTDQssbtJ9vFrrCWtrUCCsnDPmf2J
a/EhlS7ncz95nLt9CXqe8AOYpSa+WoEHVMdP7bJztTi64QTlkMJxvgnzMAQjPnvD32q9bvgFkCJr
AFI2VxFCYO8Mw7aUoPWtsdl+/CsXu1JwNOvv6UMo99H0ehQdbeeOy49FKcDyZ4O5WrySrqLP1gf+
sOyRF+GJQNuiCzJ8N5fitgIhX/nT/YqrOhptKtE8nKH7n9+J97NJPidsFEG7/2Q+2Uhq8JYoP8W3
akB0yUyw9NC9KV4RYbmq8NPW4/BxYJxhyNU5SmTB/w1Xs90+PKL9uP5IZtuSwAC2tlNn/c7jkiSZ
h/wID9J50K35PGAh1s0Os+lvo9U0OceDgjcDlZGtLq0pJoWhskKoCK2Q179QE6gPt63u0YfM2fqS
RPGIL0z9Nug103MgGjPERQOiro9PbsF93A2yNxLo7RfC0FdZFS0+IWeT2nQEw90hdRcFaBKvScIb
G2cHlpwHLOoVRNymfPag4XyjRbFIqGu1X+16T76gzURRHKAtxWY1dvm3mKIz46O/lGMJNe3LO2HD
Bp7xLQ+otpG5K6Vzq4IhmHIyHdMHYjJJ3Pkl0QXvSN+mZLBiPqeHcMosI9Rw3obA1lgCJGGUsUMe
MKN6q3JefG5FRGmSPeeadYdLyRGx2W1VE9Guh+cz/14TacdoLaeM27rirjbXOD8cVumYEPAyCMcE
+N1GkieGZzE5Q6/OjZ+EGggmlC8Ea25ghJCrI6OCdZUSnBhJ5wL6nuzmHccY0U5/PCiTASbW05nU
1gc3PiNG/drHFfZSQXK2zK4NUMpSCp082vdvtK5dicFFbbuO0qnONW8hpioryH73VzUUG8iIAWG8
/Q3ivDDLS5YH6vrxRESC7fZRXzuzifgkcZbLv0jZ8L9UsEecc9IU4S/bmkxb4j1l85H5tlhvZE1V
8ZtihRxINWaxTmnZyT+/tK4g/34L3mur8JGEz/5R/GCDc29w4NxnWbBtHUEXumvZeW3uZGY91isc
Tzyz6C81QZGG43DFtVn/nCRwIL3+Fa5OuQhovOyrDlW75y/nE0N2Wy5RkLYJdH7x4KJqEECfI5LT
LObMUsIG0CyREZOkQkeoZbOO5XgfwapHFe0XQQFAyC+1rBn9tq6KVSf7GwGkQP3c6WVAhSLsP0y5
e/Il8k2lLeJTcFRqMgAka8yyegb2QJlCrq9flj4G+HPa3NjqUvy+OTp4S4GsoiICv5HckxSEgN2j
8LJQKJaYg6+Nwt2OsVvXijsppT4ya6cSMxOWGcrfJhVCk49rr3nKDApAc/pjqvbNx95SNexcZSz3
0PqZurbuhbe9BNqUHBny4KLhIO/lNiNAhuI1FZuBh5uyrmg2HM4YlN5yX7Eg/sGR7RxJWCbADV6g
ERRb/8Cmy3Cg0nkdiYr2+hgbBTXEAXMrBfoFyaMvHGVrQylwimd1EwZGjeUTqilhfLVRwgCuRXHa
byZboHs0QlA4PFYRTmfotcCb7bxd+m2Tz8Hx8tn3d75ePW9emclYkS4YlYEQIaXQR6ooyhzzbJ2l
TMrAdaC1aCrEvyUEjNZ7vR80hYM7zfXwAbq5CTvo6xJIKaKq8qG7V1Oh5LiqOGxENyWDS9kS/JG6
Pqw8RfkpBz+q98FbYiNeIS2JAhxvTdW+HSPLBGI3pGEIUTvC95xN3uvqtCjFDrfLSotoBq1ZJo3u
jlJrvaV4x/Fnqrqp7MVh3Wk51je3w1sVj58pp+XRy8f/FGC3KWT1KKjB9wckBNj6LSgzmtIjY7hG
FZkqGbJtqsYbalIOskEGGAC/DLW/b+pm7pxjtTISQosrRlECZISlzMOrYfTX9sNzO4YBuFyvgaNN
QWFxwA91KWd5vYWLvcpF/q3LF13A5Qi3wqP2nKJAhgdZBKaJWQ/vN+wuZfORiOIyexAdtSH8bEu/
jjlGnAkLohX6GEI00rHp3cFFjMqwDPyoCFEXR9beBx1woQbpHjJlCd+op/v/G4c+Pi8HuwP/fom/
QbCjwoMYsrFKvnVHalV9wXWIMHc1ayRY8gOo7bsunPHzQnfp5tFBvqUoS9RAeLphR/imnR95BIr0
fcd2mGBxr+kxVU9mHDgl392fUxjkIhL/AxVmbFx66hUx8UyfpPyN8pa1OSbtuOMzQBmgxbkHAoDw
5mVy1SutjjrcvLbzPYJOY0MPWBSDUPWj2WI+nk11JrVe1dyjVPqE5oWcXfb+H8Aa5y5mwyPMrfLd
D/LmdO6Yad35Gf+4ycl8ahmCzSQsD67UkjZ8Wb3QYk8j6SAmCcgY6jve9CkQimfwHas1AGmawrPw
cNZMLXAKoxZlvMlWRzfzEikiIZORmG6LKaySw5mlC1VQNq9CzKXE1nk4pqZ4ragtRsiXWSR6ZDwC
U+QumYSbKwj4ePF2gYZCHd4Ywyn/eg9jHoU9m+w39zq65hcNFr7cV3yPEjlP6k0r87p7vvDjq1Ay
TDnVNUIFHYHTmmon46Nys2UbooaGR3Xoug7sihIoA4igwuDBMLi1dzPZsj8Xx5a1Ma3NCZ68ZYuf
14MC3QNu6GGQ47heFs1jZnYKwqOP7w/wauzsXBqjOuJ3oXyetoMKZfoQjga/r1m5RG2V7seoCYB3
D8qiP2P6W5EjTfsUbdBz7O5uaiOZEO4C88udarT/D4Hz3nJrkSpxtAxu2XdrRrS8xeBSDoCuaTCa
w0y4STDbEqgsRtfpEQgfK3VWUa7RlrC2SymUn29uOgZ0Tl8nCZj/lRF+j+BlWs9rSMSiEYC2M/nG
8gWQ5YVhoep8zrRywD0I6PUrG3LiztAYZjQoniw/fOB+LPSD2ryVhyhkH1/mpYThgtwA5wapPZGx
WKOz9DHvfZP0GJaAHMcV5eHCNNWqwHMbQnkMERJg10zTHRK1zyM529ZJYW5IVYBgJERlUE25aC/J
dZKyo0nRwc2aZBJjAm2+RQ0wqLq/4qoYR34Hd6y9lAcAz4H2vy5fwE42ep9e1budP140h/Ehtt5V
1z1YyNTBr/d6MWPtuS/IUQmGU7HFACWI6tkNi41VIT1w6+3jHhZRQZbzun6Dg9Oof4BFQo8N/+Y7
Ja7G8xP0b2PT7Y5xoGl0Di+0WDc9plW7+m62ZSEQ/qgfN1DzqfQKzZxaCzI79KlLNyDFZINA8l/6
o5s6Brq+iVIGfcfV7rkIQ53jPYFV8siAz7PPN9Tg4Mhqr5SyOIb9MooYqnWSHcPCw3usEGWGBXn4
3O8HDe9610aImvleT3kc2lRAnvDEZ133MH9cB5ITFTeFpn090DhCrZX9b5cVix7eABXAHrbArHMC
wHi2bwR+6S0GjgmJA6DZNkVtLcgbbZa0twqSaeru9wKysl4r+7J2oZbHgV66AdMV9w9s8XBt/8OK
wTZMDqI8IwljqB6f3uVVeMKU1j+m/YYmXLt05vYBopkbjGXgiIidgUAe5ZX3ZsORyZ3JDTKP39tu
GpJ2eoJ+jt/HGZa4Yiu3RxYuX3foDbGQaJJiIQM5utg3Ti1XmhKVHkX+MoUfXwchCxMUIDwp7ISY
lRiXpjINusTmDQj4g1hO3SasTKRthjKH2XEjuhkRmf98EPeg9LoK/9X5pMRZ1yIFD7dYzdlUWRIn
uwXdoKh95h95m2T5VY1H7zOMwne5plDwbVRcCsWeu6hXvVu+sQsBk2v5GrzDKz6AHYXpKI8RJAM3
faegKKqcxUoFQJrIk1pYwR+awqLfIBYtuQhGFMkWpBI0Q4tKgKSDQQpH+sqDX6SESuR5M7lZ34hH
iMddt2tyImAYTmm4Q7gEwEwp1iOeE7I5ImQTECl4bXSHyqj95ofRdI9rnWpUHBjEvtMVefIcL3jd
7UCU7kLJkK01Q5EbUWGTHEYKvDmlUgUAmAP+i1bDMUCFlSTIwtrT+TyShrOkyFycLEFeAwMfGhby
vFX1930UwNACGgGc0ZqTtBziHj6toBaf9FuvmGoh4EAkEB9LdewGAF9wEz30CjESIzSjp+MKy6eC
JSIXMMBwfPRox04V3xJneZfRRuqjc1WNPZ1GgDuv9cQoIuWR4UBFh9xJJR2EF35DmJY3rejImkm7
BolTEdxBmdiBQ0vxNZfS5VPwUt7jSRtX/+S2EXbiPgdcsHS4ylJGYbKZQdi26ISQ4WoFdFRCSvRE
A2N6vfpqdDTzx8gZJkjvy4CiJHOfcqsrC/08D1i4Udl++CIsCScXbNcg3AKE9c/8PKqCL7Gq2cSd
D1uUQdJb0ye6XxTwxicmKk1RlEeNTW+8BZ43TCu1bySUf6W1sVsW0pi4s2N+r8NB4/Le4WqhJGJZ
tlOWnS8ctMP+43JPWpKnlY9FGJ78QuuJUB1RJSbk/VgK9jhPQZi7HYHfD6HogA9OgsEmrA/FHlDk
fGfRoe6a0x9fOffEA7hShKUZu7Ao5r5ltAfkNpk90tYhN2HsJT/hWK8HUmOkqHvMrvust7St75bl
atTHFs9gfHLSxE201TtXmbKyyS4vBru+GGw3ZfxD1qfj+xjVl8MI+2nVUyD+gLbGltHZHrxeM9Bt
pSwhOb6m3dsvg51LKXmt6akS77V710XW1TEuExbtth2i2sMRxnIi5pPCoa6VMRc7Jem5+Jm2ZL/q
bu+ViI/oOJY6R9jomxRzp8ZJWAr6VNYiE2QiSES5CH8IXADrtafX+T8rQfgCYt1LB5rywguAlqsD
pX38Pj/CkPEEKHcvMROsvMLf2Ea5fAQDThz4+UYTZwH+YmSV8ZYeXmvAKWLJrqAdJ+KT/wdKFHf5
PdCrEJv4YEvw9GhA9bJZ7TxO7bs/4c+q+DttU+FFqYJ9uIJqQ8uUttHCe68oYU2IoD00KcH/AGN5
/JjLd/HAw4E47TFzUrEXBftQS79+beWH+wogL231DGnGU+CPTbDx/Yj3xOPoiiT3Ie5FCVyLB/eC
WWukuXyfHfz55VU+GBecUnVQvupBiXhcc2L4/KR4q0X9orU4ChCV879NbY2geBiZCTMoYzGKxVZn
dKfnLN05zqgZlsWowTFOl4q8734oZin0k+aeLrJFe4ubVPsHmECiQbbqw1ERWAFvjpdLGA3ibjcS
xFDbRPb8AxynmfggfQHJIOoImUgJt8q6yWn7a71Q7biGPq1uc6D0RnjghhX+teziOYFnlQMIa+JP
wXWKKEv6HsZUt/WTpLZEa5o1bL0YnARd1nJhYInITsrtyu+rGm59R2h5M8VA9IFmxz6BrFGOkNsr
4nXE9YXUKf0qB712wsBZpMttnsd0lXvMoPl2AndPbsxUlcfLaOGzBUsl8qVWt7yzp6JJesXJ9Ccl
bH6Msrf7Yy4aYinPKy40MP2cmp5moRBefu29W0f0N4XusiJbdbeChwsjaHrmc9pKAxjuWun+mjTk
E3SZSlJYphUC/rlIWUCqW3za4E9CPo8+JmVDfURvrTs71Kzy/17QIer2jK5BVXPWTqnd5TlZbe2V
JtZeqMZPNwVDh9DuTUqnfyYb6EpwHdjCOBniLj8IFS/pWdLx+b2nvet3xtXqqw334q2zsDK5Op0H
TfCRLY5jNbZTi7ZCHiqH4sQMtLJIdjYpH8AVfBSwgr63cKT7AXOxRJ4oWzFgGZaI1dSdsjHFfqpw
JMF30LkBZHqzpz37796b1KiTybIdFaU27jcI18N/Us7HHOyvxvtZTtkJ9QuauS/523cUMMj5etkD
tJNNNuyVIfLLPvSuesG2uuIUukTztUKov8wnXVmoLm4/C9B2G4hG49iPiiRAQxz6sEfUTdL3Jj9R
+i9eMbyRmWgZdGwE+a0QiEpjWnixEerDB4ESBmsA6bzt2DS6E6hazknxMJWAEWHJc8lMeBwNzCkY
On2XriJ5sGATMVjXdPj/fMLK2m/uYtoN3R6j14YuaVqYbNVrxXXFYWcHkzJ88gdSYyWY1zaZ4cH4
FmM21ZKbDiwNLOJRsGeCNKkg1BwII21I5DT4wroqJKEoj5Yg3XEUrpsuHH5oO/Tg3pIShIRrRu5/
RKr2I+vHUpk0MUwFoNJr7XgT0z2pBlIugYMpWxJyq6nydFHvR1bfXZDE9gBbhQjNvTyScyFZ6w8I
9RVpNPRbB8POq2BzLkhA4w8xY8q5cI44zhFu3ZDxVnYjCn2BMe9gsxUsMFf0bENFjDP8GQl4iRKB
ck+OZsOVQb84TNJym/eQE8gbrk42lXTcRYmgS3lnMd9WdNJP1RBZZ3I5svIOV/fuz9QnWjQvVXj5
Dnp/RlXEv4JnD9lx4WzwBKQ1QHYfO9uISCc/rUHXUvkQRNoro/y/7ofQAEunhDjuPYBsyt/77XDo
Cu5c3JUKdwRO1EblnIkskWDQdMJ9rUp++8ngyy+f/FBZtW9GODeFae0WzdZpgikG8oBpGLbQyhw9
oZxYbUk6vKijorp9Fs1iVDLXq6zqxxMIjMrzANkKFdPN0XDDv5/3HuNEeHVjyXiT/KWMs40pnUUD
F17QwWqdcYF7zvIIyl10bTHaJHUwhUTSdDmaBBdZOmMgyDLbrI/Km+lQl5c3/eK1MowP+eqW08SC
DczhycFivAlgkOCoin1mNuYLpAPmuaB3/DVYLPIXx9upFzzIh3ybfdt9MB5pKmEKI1q19cZ3QBev
u2not+whWgm6QzYV6QuXXDBs5k1Oa1A44A8o0voN+f6dLvbCM1WWAko7ABeqGJ4LF8VOPdQKDZ11
Rnd7jMMknuzNu/36Y8hIUX0P5+zsr1uXO2ihPjE09RiUEhSo3m/CW+ZLW4ir8CQFqYwELTHCzA1Q
VZ/AGWBQ03c5Z7U7iycTAP9hrI2FsIY/eBf9CNZbELE+PY9minodKPyBRYTqI0NvhjWelqVI3Zj9
r6soy46ut+LyfJjH9LRykviFdClWXWGEtSAK4xIiy8labv0osJiWMhhs3mXWU8+/9XSnYBVfiEkK
cemJFKQRQlHyM9rJXJFWTYPA1V8ZLe096tiXkRMNHv6bVp1T2WABWyQ5ANsm22FRCQURHHOeqNSK
0LCjookbxPjBAZUZqzX+eqQ+iWYgtffVzHcHROfSyNHHoRhBArYmvlr1uHRkEfaLCn96Iu33QA+1
ZDXjXG6Z+Q5+w/nLwDE5LoxIbjxviWpba1kpqfbT2yi6cY95e+JGniNMwnxh7OCF6ScJfQTGoi1j
DJZG0OKnsCUHO9gInTCwE3SJPRGiG40xWIXvX4llp/7IxufKI0+R8EH1SiIzOyPDMMEszBeIjWwG
PquLCEUI90GhIui8Jfsdgqm8vN75qcgg5b37/d8Bd7/usMIQw2fv3kkRhUMhF4+Xv/277oOnVz7S
xjKeSNd5+4Bqw+xjkabkZWgDtULz4+KmcCz9yfIeDs9hZTDPIgdaW16UJ8SQH+Aam3YVSLaaUb6D
0hdH6XQcM/Q77HsEM7sW37jsII0lWTvkAQ44YMXDSCCK9t8QkTME1YHVXgKpqHDQelQQAOMI/UZz
gsf0fctEX/tCJ0KyAHrb4xF1RLhbWnTw9Bz1McM7oryBeiwRh9PG73iP/WcMmbz6Gas/OHQVk1r+
sEDYtHsmXMD0VaDmScsP8afYtpfKuD+trKFeHMTTplTgDFlJ9g==
`protect end_protected

