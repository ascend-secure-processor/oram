

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mt1j6kuu3+cb1K2ZJB398+FLDRNfQGSIdQjXp7qmVQmOQHPx+/rlWaa1dxNuR7NekpTe+npQXqFf
SXZR41Vk5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GzMy3XYHpujLbH1VRMwcnskKBc/VqM4rKnS6c0cP4yPuUMIsIaAk84+K18/IiLBq4VJntGzVpTrK
nNPZphAJn4V01s5T4oFw/WmMDaIuyrNZ460qU6SNP5sJXuq3EhbY4B4GR+o0Hvcuc8QMo5QBzZDa
k5HDyO1dRtAjgPYgYtg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AJGiGYE9s/Mdc+oo1Ze58OfO5hGRr1kGvaGRV7aUokiK6HDR9rWX09vVk3hohi0zaihQ8YHHiE1J
cY4XbMg8CM4Wfx+OiYzs34NMMZIFCIKpUfXISjObTIn6h1DDj8hFqmTWmiyEQKqqbjglZEE8D4DW
hegUO4UFSKebZI+ZPGcxR0SSRD8ZqmJZMekxNW7SEr6wcoys5Q6AfOapNGWCmMR5vmGTJiAj9gtf
Fn/Kl5f/qnZmk7CzgrCaHyfJUP8dLNRR4skdnbLnJzy9gBFm9DDm+PyvyujH/QAANF69u2sms3dY
3e2Jnqg8hjV77dbxF4tUhVpRVKMMlSBoAxEEew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nVR7EPGvZP9aSMp1TeQGqwX2IVO58loMmrCMMVAhTm+zov2RVpPn3PUQ+P4NJLddCCxS4PYmRSAA
a4qY/1LBxLfCShfwz+Ry5uLC09qFfQJ/9TCtlAxC+0xnma3yZtiqpKsYjnNz+APEV2SKZsN8T/lc
QVi94H+Teiux9vcF8h8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gLA5GVUJ8mNsZtD9Vye1GMuPTQRcmBgyzSuTdfHAcVLzMuc9lA9OMZub4mklVtN8nuKI34+By7UO
63jO8lXVUDTrf86yc/uAZZGp2C+XR5TQ9zjsdUOzGdzOcfamMfLKG/JBFZRIFdvnPwCp06hlSPGv
S5p/9LKev4ie7V37qCXLeNZ4PP7BVM2jGTUqkZJMGRMVL0GO4Jg4fh40u5OGonvv9CqHTjqp1ONO
q9rkMDGQJ3Cm8TCYgZDnjhuladgRFeg3HtihzT4qJlpwyFJgt/ywu/FS1FYOsYp8HEsrl+j4gNcr
y+Jo00Ir4CxGea0b1CdeQzk6RR2zoqbAxDwoEw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43328)
`protect data_block
/340aLidm6JxqvohAejKTT9uMz2bAuuhCqdx34Aa1nK4aEnUnIkgbPmVfZt3R8nUCAIcDCFEoyLm
w+kfL+ACFvlv/UETote3xRyMOYBPEqPGpr6lpCWoo8ZZzQ+8jnrJpXwXbuIWEYxo9h1bPLaKFG6/
VCw+UlMf/e9+bSsc3C/TP/Dy92h4LTnEkZ5Nm79f4GfjMr4Jej1BK4EJomJ+EQ+WZqo+PXg4A5bc
iNf1n6eaJkAacWY34Z1btzLOdhOLS9KsHAFFPBbFBneQ6x4nTC6rAT/U0KayxmqALYF2gfaaTR0R
5YmNZBScb8ylONWkNH5NXrHdEpcx2RtYBXJzfKVxHMsPMEaSZePv0daj/g5Tnhm+9SA4WM6NbZCY
DQbPx3MkGnxxo7Gs1AZ8NUj+da7tZQdi/2WX4tEeUak9+4ZErojVe9SLL7DZLqyn/OcovGTXWmsW
Fu5jOmvVWSPshmdyi7byPcikBU+ikBx/CtY2bShNeen5qfgu/xbM6P1KcG+1Er92LqpN4HW3t89F
MHb4R1sOEUfSpktEoh/RL6Bxk+5U32I1aMpRlOcEKvrcfnN6wOAIy2ffWLl70L1ebYilJC90WDgS
6cYfnldaCcSY1CMDQUxc41U4AsvMVFqJE05iBpajXIsdANsbDWrX8hr+s49pPZwkXxWDrSi7P5qb
TPccXb2rKV4h70XWIjeah4YmLIt0eOni+0SE75/Fa9JsudkoSVjPpyJNDH8sIkb+I8rk53fxtr2v
D8XkjQGbXfJ7NgkvXfm3w0Fp12MCTVkltGb+ErTgFtAQt4lDruQzWEPMA5TNI67S/GzL+EqUjR+b
m5HAgzuuGPW3pd9040jvg+1AFrvR7vt1nNRRVL4hOn9ThycVNGRhcQIOChUNzoCwdEyCNhOS4kcO
5ch6gj1zLANLhZvVB3WUNS4g4Oj0F8Mks41u7Fe1Uoz88pTXfBNo5YENalL1GHGQbsUX3/L2PlRn
kCofefn5GWq/t/DXXiquUjQOFM4uL78wl9aOKCdIN/+p3dHzFHXJkjGWPVgH+Bu6vVl7QkG3b3o5
RfA23PfPx0ktiVshrBfXdgSHsyRi3pGNTPU6ZTkhMYQY2ptJwWEBscHOSenLl1R3qEl8NLvFVfIt
nX/NtX3jCI/vMlRZ5V7anZUqAaHhMrkTlS83PuEIiFF/8/fxljBTWLG0+2AL2k91NtmiHSMn2DCZ
sthPEZmCtfIcJaJMcYcBMvSL/wM8UJl4JQlfAkoR/G37qZ05Fu61/9IQFsHtYSXfC89m134XewqF
d2ISFYOMW8Blng+qBagfF3zLduSkeD4OblbH8MLPhhJ/nqpWRfsKo3GiYjHfkH9rlju2IHfyCp03
EtuATX2tZszMa2zezniGw+SkVxzEi32YIOg+pfGI1XEKteOlGLaCBeHJLz1wvXWX4c4Vt16RwnII
gaFfF4IB0GHxH4sDz7L1SFztgovFtwWXYj979YiYo7FW2Gbn2H8SR//U54qwH9SC9ulxRcHlhyMr
QEDwLQ5uRp2EzORU3EJl2pWJDo5+dinwUrls73JZXVtaUUl2bvnhHgAVYlyYeE4VEyhqUr4u5X8x
zK850Eq+kC2a4w3W+uMinUP23LHhxF6TrAKH+hvgraSaYtb/Yv1hsQbjouWOBTtDaPzhSCOHLzTX
601VulMPzUEXZPO+HoflF3rnQ5yEPYtLHvpe6QxCIa0bQ94Jd3KSg1J/XJC3NCelTO9nXWz4NJUj
Uod0Ye50fTF9BFIcStRYnXoAk5yQK/GV6/77zCJ+m2FBCpPdwwRZ4polE1DDOWH86GHmZeSvtGry
Btl+7yXa0delvm0Xu3dBHhz+6zL8Yx/aezfTOgHp+yxMyJGaRVM4bWc6YbcmkkAdZAVTM3r+HR3i
D3kC4F49mTuUzgrlVIXFZ6+p3UucteWXabop7oa4LDkuE8R0W5eV2VEATwugPxeKt4uXkqEIyild
D/n4ZIlac3MD9EMAerqihz1JCP3CkgkZRB2dzCMvwk8P/8wbXUzVhNK8b9Z6qo9w+SK3m+wcB98/
I/q4IXtq1FIHNZjeNFdhzJDMzAYM6eK5a33AO4uXC24O/9pQBgOPeMV7/VYxukriAJ0xPYCMBxcf
bdoltMcOxJ+K5c4XRxnQSHwXIgbTOiAd0TFSiAQgp8uJuxmdYSrZz1Zbw67tZSUu0vs4xrXz6Bbl
vZqETsxfufEN0l3oTQkCngzhF9ZsWLqHfoZikFp7jdVcdN4MMOytGoVt81Pgiy07NvjIFrywm3Ho
udFiIOBvLgEWA5xIqHwbUXi4jLACOZ1Az+TQAZNKV5JMwgIM/eS4AXge2F3WYLwWdxe0f5u8Iw2h
/mgM1o2SbTYXK42x9wWi0iaIjA5Y88sVpjY1yvTp29V0+db6pWm/EnfjovdGJZEE0V6Z0UGDCEih
QHHynZAV3gLpUCjtbN7oK7K+Qo8d5oY/Z+x+fswIfNo4ynSZkk2J7TH23ZkT0ZTf4WDgIaGIGvbA
OhkiQF6VYiBVgPsFTcScoYMtjaVBDRd7ohx0K0ZUq0yeioYXcmztUHoQ2xDWFtxcZbEv8hI2PFnv
R0eTjYbzy7NR13K6DpJQ3mN7QmU6fE01YNLFUdMCz5aNps8/n9a9uaCO8gB7D+dyOGKmLkLLNuZE
iZgl/14n/EHM6bGr8C1tlpb2ft+Efw3aRxyVBZRMF0E7LxX6sIqN/KKSprCplRWvct/y5DkV+4a4
IHOQht+7zjXUFJCkdjXVf243qprxeN0tF5J8X8wYSBq4+UJGUAU+ol0SOKTYujKhBtbRatxHYjZi
tSxKetMNxyfxuMQbILF8xRyWpf3lYwdMtKNMvPhafW2Xamj5CBC+4lenOK3fhuAX+yutDEhRlkq5
7c6FablgtDAKh9qe+vbR3irDOxb4ZoQ9pYw0nej6LewpG3nlqftpdy+zj73hakeDOadK8nHYmx6x
+YkVCztk0lpFox0xHePe5DlfVJNGGapQxkfEyWvR/k3epg10d2gNExMvc8PRYkM8t90toKv7sMsn
zrOn/LSgPkfn+UtIlmAH8a11pKwWMCaxUTor2ejWUFuoDxoTmIw5wXUN9jhjRxZQDBqc6HprU9nn
DKBcsRTfv4PMY9JG8Yq0cHpB33LyoAqnfzlUoYhbtnKoNKaYi+VUHnwez4fSvvGSh434GqvSZZsO
MppeqgLdeYXJfV5U5KAFf5sNXQSc85FnmYTXfbmdW2F6PzPjjH9o9VlAHOozR7Ml5Hnj6LgQ2kjP
8hopk5TYiqakWWpIcNmHt0QYJe8bEKUSY3Orn16FBMoqeQNz62g4a6J9rbhv3EdcTAqd0GOmNKmQ
UybRqMBZ91bYRgktY6ImOA3sNFrHw/JqLhHHulEXWherOj1EVRzs+8I2Uh/nGRW7/OagnbV/wVr6
03fb9LIE1v7ndoEP0KmycCfh5V3QyTiDP/jWYqXCFgSlzlgs7gbkE30NvNVigrzwuakmR/UB0KnE
Zev5TCTeZeSNCmu1BOgsNiKqt0j1mMS68ny1lry6Xl/97Hu2Gjcx8LEuuhSiikW9dWwlZPn6v0IB
KP1K8u0OQQY57sgWd45V+e2UFYPrR9MZ+HqhXRyfKXSwvlR/qK8GlpYI3N8oLDlqpTu0LMGSPsLx
IxiEG6qwQL6+dpmIUzialg9DrXPotL6RVSgI4bUgPGGc2y8J1pojaZnaegeSKMhWMBsUghYK5QYY
4CTsYSfNrSuoTjoE/AlQD5ZdUXCbdWizs18e0sTwYQsEOlhQfbbumFJX8a6VnVXpWwaNXvAWdPVq
spV9fR6NuzYzSrVMduHVHVmmWGH5iX1mm5bHUc1yf/mZPu0fw2YXTWWlqS5B/JrecXPivtEdyAbj
AVBEHGcgLaL+UFq1O6yFiYBtxpfjTaRgyvltSdlFdshO+bcnLhANLsDKoN5Bg9S31YtJ1X3lvoZT
9ZVIMkZBNo4xXGkA1YCuqfaPLGLZ0GHFvR4rmCDbO0a0ocZGcRWcyY0FPUQtPvVihYLS9SJKqSba
t5bkI2Nkh/NryL05Fnn6se6xj1FHQOUmmrg9/aUW9X9/KzJH0DBZHfFYsJBi5UbCHZ/Zb/6SaaPh
PchL2fHg5VgQyAjHpofUkWjhGNqcxgXq+UTv1W6vbm1UMxduOfRbaRNdjbhioJIZBMVJMzJcjozC
Ue/yY6sJAJmaSFonbRNUFQFYHHA/VHVdyH/iFgXhKr+uWPmCHA3Qi0hX4Z9Esu1XF38BkzjJMWCk
h/OElQi1sayBWj3UfmhQ0pg6TVKpIcU9XsbZIxnxLG7ldl0UlfgsraT7HUVsyLVzKcIv5YGzaHH0
nh9DovE/mZ9XritBgTKb/VdyrJDPfDF8xg7kdvJ88fW8MBteGIC4RQgL6cEVnGuTifA2MA+wjj5N
3VrA8HSG98fBmEqeVKR/0mFjx0s0o3iGao7higV4vTrlojB8+vNmYg2YK5vcXzpjQJRXT8CR+S87
WdXjpvrRjMULF4ACyCcrYLckmXvHO7PUrmM6OAosZcPwZRzGKa2NE1dbi6Pyc1wUFSJJzW5jvcsy
sVff4/n29UNMUwUtxmkIsNaNZC2ag9t00x4R+ZecJVvQIw0PHufh4w2NZPS74edRF/i1os/CVrTs
oJKmRzZddND1Bz4uYCgRmhxfqpRU8BL34MoMdgsc58HJoJ1EFxYx0BqN8/efXrPL0jRzAxesKPKq
0IwY3i+e+0Uk6dhIWNE2l2JOQRNpuB5ew5jW00TR6LTyd3yRGYLmwxQI+61UiaBDHjhnR12OyXZr
Y9BCFk7vvqsCgjlBH8ce8y4t/JxqMyjkMGkRzoc+mxOiBXjAs8GkJW0q2VPn1fcVdhM7nvGbA+vz
wQmCXZQsoN6xqwKFdwVw9vLzuUiW3ky4WOhUtguLrG7WDAwTzzx6fgm1K2HLivY2Ogc6fLpu0v6s
APcxpKiefFWTfEKeX3/T8wP6yOjmpaMM8edeJq8TjkBI9dBcBK8ns+84/vUj+oJbdR0QW77ir9wo
XFXP2Vf5H4KX6x6l6nws8TWhE7Fq8K+PZtqUAJh7/l5N5hWQrgnVu4/alZasu02lZS5Ws88Qg6wI
pfrFYb6J26YVG+SrErqswefOdFw5SGvwjJihJZ/mLUMN9bjI8ayAzuJyo3tVkm4FvJLKZSxZ2j7f
3nLcuS9NlZ7xF7niEgssY4f199U6bOOATwPO7k7XlourWW5zvINixFr2fWQMMLKJjH1rVNwLVR+j
wT5IN3gJDeZUhvbs4+0Kg/t70UEjEBQEvW3OG8bzMh3HxXig3AULL9QwdOJeuCP4jepniYpvv20u
z/Ev+G22p3l8HX7Ou4Oh9DXt/t7p7EmIM1P+i1qzs5wuhnN31+wKLoLwhvM3FRmgPBXmh/UtXjEL
+pkq4hBZZkpqFrSA7n8fU4IQ72/mRj2ibPdxjwwEYC7d6D5LuRk56zBb7iyqfdBY8ipwyUCCrmhn
6LdzwwiNH+7dTok7tlTOpmKdR1AyVIFWJxl7v8hwPwnuokeniZQNXR9j7kOEOqEZoqVyZA9mGq98
RwBaIUIgXxJcw0uZU5DoFA6lyD+Bvy7Sua9RhHXx3F47xUiUEXmIB8oW/VkYF+OnodqoPe2ev1KU
+S/n+i4Vohz1DJNgaYWO9kybDxJGyAogn5xeIYjfdCW7PGQv0IHOaf9GoR7OL5JBdGbA7qUK2+xU
/b7bok33JUjznmJGXHZGDKMmG/Suusd9xFzh3d/77jPWlhRa7lhoTrrpJZaCGfyTuEkRL3LzNNzp
mpsUuPv+bX0+nYMpINpznXYs79f0aNAKSbCJa+7aionH7WtoyywnYTkZladUcnnycqYv9LuMftFL
p6pxibi+Sp/9MG2HZdZpwuybWnUwuY9A9ECmN2vHVE7+CJI/OCfbE7YdL/bIPOnZ+tqRblZgxDJe
wqFLx0rVY0pCTuKPLQ+lnrzYX+t6DATTlMBoOzkQSiFWTyAqX4Ymmt9xmQW6Xh0rkVD0u4s1v7KO
jhRbvfyRZqtzz8iHtJibSYYU7Ftfl+nf62WR+WhJnU6rxAdVTQBScN1nCLNYzrMpPPkWIXAP4K4l
JuxKF0H5MelnS5wPoMM9dLl3GqiVXDLg/rigIDsV/OeZpRQU0Zbe4AWLByYWbn8ztqdUQzv5SD2o
xrpbTGFQydRnsuXGQB5KExrLn6H5IYobzmbgeOE5aXUNtwETHZhg48ipwZKKiVpEkb5/REANRi6Y
dXsgDyH6BGEbqDIBK67sr3Nh0Gu2+RDTpa+LKQH2Xs2ZKOeMgYex+NieH3aJErNJvvkKgncy7vLG
STMq6QzoHrvArG3umPkTv2ImwR6V0IWVCICsjJeHUbObeiFE9xqyXdt++JDi1wlm88JoZ2vB1ork
KcWB76b7x5AjDCAR4Bepo9xwBTtyQ+50jfVTKg/38yu0MOof8Dr9EBeJ1Mzz5rFdnoxq23avP2WR
mO14YitnDbiUd9kCeIl2SsAWVP7haU5PS9jWvEiKqg0BLe2L7e1oD8GcUM9w3voK++2cO5WWPAuS
9asuH5FKr9aSQhpWcBUjlfoeyjG/IqmoSfnnD7wO6DJjUTlURTn4Z8fUw0d8uU+5YtKORXIOXhan
e4yV7VDPn+GxyxNpyLEI07uaOXvbmWT8lDb24lFSxsTnI/9t8PzmtksmLxSLdKv1uXyf6HzKVaI+
cJ8WIvYqvUavbjSJeY3nmIuBLiwxoskowjmr1FuGXW53B/okvXOa8bKeH5i+GcNjmM6QQrmxghGI
tT7vYwDWAYDXDqZNu4PfcYp0tLRFWMFsJg1tIYmHTupWO9PgjP9XXxQX99F1TrBlLMS70zmEFhwS
c8aCZPfPquvjQdjvF83oV+BVmh4hf/ZmwAjmxWt/ScRb7DqaE7/MgZGnGnUnoGu/ycLRWVk5Qxva
uKDwUvAVheJZHpUJYguHs/mS1Tyh/E3eRK7QLCJ2Psi6KnoYVm3nSoJ+aG74zfIppA3qiu/YWhI5
nEe2xt3VdBRfzX4+7g7uenf1pj93PFUnxh5DKjr3Qikaq6X/O2o4oe7BB6v9dWY1d1YLpRxDwK3/
D9WtoMOm76FwRbmwyZfDT91o00silttvsDnm619alMHsYyD1JS20EVvqITFwS96Oed0uJQwJayhf
4AeN57LxaenL03xaO+JAxekqTMTpZTVV7IZwjbSKSkYDsz8FSRAJ93+kwQULORZVWuqlISeYgZtK
DsYesUNTpdqbXSYaVFHH9eHPTLTCtNL0XPrmfO42Ys94SdX7V3gkisHksXR7T/+Z/JLDSmRm2n+h
u5rSUOPg51ZDZ8oE/KyCjAm5ypKPn9P4no7ldn0te6pvq4fFwkAwqUOmNbxBsznF3C72sxSv4/CI
S1Q+bQU5sS5N2UU/wSiN4xpo0prI1g3lFgqjnhA5hGFHotq6kYoYwKsF+QS1Qvj2ED0T9pfgmpcR
dIELTD9W503zWLTelU6tyP9LNE5ovMGLF9V8JLJT9kkd6YsNwgnoA78sY7PJLE3QFrXKexJBepYL
KmuO3gObEBWDAjL3jVGXIP9uqAwyX4M3RG3cWNKCK+1HXnOWkptbZFuTIjKGRr6wxrAJ7QfvPWbP
BRqUZirqfTkBtubC6ZWzv+NeHHtvHAf/61j0cYNxoCmbK++VNCKEnPKx/J2UWGUqqlFlC2BxG1aZ
md/QeemLYtLMa7VXWTw/ma+fBoTvDm405YGhzMxGPlJTbBJXsXJECwk336lUS4WvPDid7fpkQv/T
d6REuC8AVh3NRpDKIpSlteW6lAtq1qgZtrYLumJX51iMco2KY3LtD/reft21v7GYPm/boLAvlJVD
F6qgYXDyClPuCre7fv9dtKj4xdV21ZEw8gZ61s+RF48mhPflZnhZwpRwRJR8e95O8tzp9lf8Hulg
eOvEUUoBnVvw3pA7w0M2BoxY+v3nXQ6PPny2LuQ6kOH9/glOMZR3H2UlupgJFT25EX26vzsXokwa
6CAJf/agLb8kjjNCpdOEi9IW5a9gOquGOty7ldRSty889e3LyZAQKcCWP2DzW117x9jUAk4cJSOH
Qh7ze3mCnrjV0c73ptxIMTHUTncwDB0LzdvH7a3HQFIaQaPQlcOJUYg2Y6MjZVMJiEcsgWauci4k
nEp+OI72pyOPMRbJq4tstnBYkiJbHAZO16KmKaVb0xhgXTnAyeZGrA/OW2LoJEXMwFd6Spj0kxh/
WJ3Q+gxu4gFdULK4d5gG6gRoYE5zQKlGaidhOfXTccXtpOBrdESOQ8i2YTm4fXbdC//SeA/UnN7e
JyvBWk3r41HGzUFBDNvTSi3tdSZq9k/6xtSIVs+ncwIWcEY+slCP8YNOGcptvsF1JEgGnFq6CkRA
kw6nzj+0qcvCFVUHWIyjHUaIgTsprUNcM1Ic5NncY6oi2Fy0sbk36iPT2Y18pM4uDV4SY4yjmN0h
ARlWHynFUiXjuKm4sk9whBXBg9O3lH+eJq07K/ao9h2KpPYWjM30YZf8Ls0XDduYuurbNmuhq9Uo
bBLSm9+8tTCVXsKtPyFWZOfEqMIILVIfDmoVB+j4ksobVJ1cU9obcOwaeEBXPTB3UOJDM842NZ6u
YT/ElaZPsTaeZCB7IHvnqDQTHl2wdgwvq8FtAdSG3rpaeiHzfKTLjS41Cn61BnMAEJaQWj5dtNde
2Gvr5kD1cvc9fMjyjSriZ0DYA/Zlix/LpnKhdVomIFBExjeWNJCbPb7z7ui7TKNsGTFoWNLJ9GoH
I7tnINlnS+ZA6SXirATN9W51kHKd7yOuAPX+9e6PNDqDY/IsQGexCy4uPBxcGQUDatxlvrT942s7
1pk+opYfN2YisCzKXa60RB0x76YoC23aRelw+DdDz6Fqpzjgti4HJokUaQmH7+nEMhR1OOHMnpom
I2U0yfjJ+/GOupM9bkVhBo6m/BStrVlytKq//9t+1UOiILYkm7qCA4Fk87B+fg5ruEwkzkIPUvuj
QnVFHEL5RcT+Di4N4bU5Z/KTBKYlgzflsRnNYoR3EpBkNg4wEt7R5jXL4XJWdEhkSmhz4xLKPiMi
JDC78MUgWWc06RQTVrCn2IieQiNC9bzkLXnYqb7VkyOJCM9tLGS3vMNZdaMQ2hAk+a1BSbywLh2m
2dFoP+D/hYr9iL8dJJ+2gIcgp07iW0Hd/9XqAE5vsJx8Ve6u9rFwcDOpvZpHYwJ2iULIVuVFtkhM
zdEkU0B2XkE6FprEgNpBOOO+o7f2FPjxSieosFjPqwXH5BMSdEtYwWFF3l1ekD8fj4tjUR03Z1pE
ODDFy5MOTEQHWVoIwiC1oaYkh27Aeum7a5t4R0BF2H5zC16pxRlOuer9clTAoBHYExsSkyOR0TB7
C2yaEA+RQKzJKLu+W5yg8zAowWM1SYX8SX9foZM4Ot7V/txi6Hs15EUxFjLxPl0z4ZLr4nUGkv4G
3tnMzCxx3RHtH4BlhgW7FFP93X/MehdFg6pUlvfMXaU/R9jXN2rbmYqYTNudwXzX0eoa9ifpCX/q
BQ7/SzhpdriVIDukj7a4KzJeRfjJ1rMxHQkjhv5JU4J1Gy7MHWZEs9exSJSF78xjd02ESBaJjCzY
x8hynFUTlRLPg6wTmci3ekkHYv9YJxpgtjAIjB2RkTcwkabBQcx1gaz+BQxGzFrrOs4OAt9KK6kZ
3IrorgrmWQH0xoTHdoyCvqb5Ag12v4sesq2UQJmOM7EnSHdJdjvIxgu/9jqc2QSnemG2rFWTVjbz
7KkFNTiJJgrPqCQMRZX/hgnATixksj84QOpMALXtpque5Fnulhf2iC78xMiAV5Iw/AqdvQ13IG5e
UITuTr9W26SsEV+McXDZvs3ZSmOFVGV3KE6iwtvyeWwrqAUDvltMoh/CmyXrvND/ZbslqzhF6m79
Y9OXmPxsuYHpvqeeSZhZTSp6hNoxSB8g3vtciM22rKB6y7LP/SLlx7hYRuuO43cMbIQqGfAYdsAG
/9xJ6XhDlCTwLkSGnIR3i69C/0mAsGJQn1twGHo/hxmYs00YlgW0KNwRZyFiY8LqYOYwYYk8D/dp
flYGfOGSPmuOpt3H9EjfNCkHX9f4pnxd8t5KoS581d6gwdcsDft4ji4Wo1h3SlY8mMUg1fnElNuj
vRW4UmuP7Ene3ebMUU5N1gZdM80+/0S5gNxEfI1VjjMoei8pmLqJMRo7aAIjvhFgkoBKN/X9RF6t
LdZJETzWA7bTLE3bLpn2pOYRqq4gwT4SSjibrZYD/8AcTFbfQy29Ufq5ZXsccIUNkfTv27Q8nvYi
VWZ0u/5XX7xptRaRKRemQMo9tRm6nJ1yocXSZVWbYSgBqlgz7zJ1Y/zvlWR+orcl2R2VzXHIeltX
bFON4k7T/vaQy+s9TDugS5Z+jNd72lE5EnazAN9cauLew1NGONVqmaBmg9hYDnjZeSbQ3f0Xcls+
zGbbRvji8ct2jW/Luqek26ljt99l89iNQxiVDexNX5D456CKEsCQu1t5bEhEH2ePLVQI5JxwKNLh
oiDMgaB5pw7UVxLoRD0i84iiKDKTxLwxP+6Qomr0cV02dwzE7YVnXoqfBgeuKv5eCiyS4piOdL8Q
dD+dDu1KVLT1BhGDLqzJIIpvjC3NjtyU3rOYXLJx/Ok9/dBU75n5oN9EGhKOlsAhfVpFf1XUvkHJ
iJ/1NijltSnMN/WAY0Y5qOqexURIhT2qamN8E6a5DWZ7CoKN7923l6StFKUAOZQ1uW2CJIpZEV5H
6Dydr5/UOAFR2qpLldoeZNyogfgt3/KrxO1WPMwWUFN3+NPhetsjql6ebBOXS2sDR2cXAhVYwQUR
jKWqUiFP0XlaDCfdS6y6GvDxxq76iyAJ3njBtJ2FDyWaDbUSEpr0oKScLg5k33vv34s0Eibz9ysU
NOuesYDYP44cK1gQdsBoN5KgJRuNj+hyIZgl2zxf5XtLKdnbDS9Mps0XJnfklOmFFd9YqvTNwUFO
ajsrEx+JPcKYmJ/5Jw1cd08+pnskYlCkvqY1jtqvKxFqYkea5PhebyHl21G/3yYRA589laGfS5Qu
fxGGdT4l1QvE+/28osoKBjs+ukOFmJckTewAXXsyjJVQ60iphq58Saa3f68pCd7FWWJ/A+nFDwUL
5NQb0wXMvJKIbPJGHqKxc0CN2c/01lflLa2VyQwTw/MFopAj/g8lNq3zgmkeXmU9Oou/KK7rQXEM
aXrGHy6uUDOukXymrodmz/gWoly72IWmMNj7/F4+MLPZYxpd6xBAfg6Y+jU8da9p+T8R1oD21hCC
WIjMRQYRmWtfNeMhEqeMMb2bcPeyHjHnJvnUZxOt/Y9zTSdiUlhm5jNf9CZLqZ0y/8OHIebxPGJS
sXKyhWFlxx8eXmU5b9cFcz8elfwoeO9viVZg+6SaH5JoVYMMhaq51xuwVJCNtAseqUMG1H+w7/gs
xKyd/QngB7tWqpRFWKrWvYsxP0MJ44l8CfQHYMMk7OECQNWgUPifCJJDvkhZyEusz6NY4Q0Vj90u
q/tSQbPTq5izIqRFCap/slSA8eYR1bgZquaxPr/q8L56xxVuJEcT86OWQPUsSN8bxr4PxbLa15E7
rgs/TGEc9aGsyYsX1LeY7//Ycytoinewbi/7nKOVLjZgiQnosXFgxSdxTTHaM2C8ICnUwibCkjjT
Jga1Ybi+/2eceYFay0KNX3IoKu+m9ayvbGhWRRcT6OgIjIOYY6gGCDG4Ob2AXrRa7x7uQJgkl9Kw
hcQu94PQMp4pIVxtJSDYF1yYkLLNEELb/axNt4jxR0UZSkebw/LGfbW/msdh1ktPUIYryNHZq/7L
dHrTcr7kzUia/KtldrIfCaM6Ve4JfIaXdnbaxIsYZY8NvrW9gOWiGg9jZjRX4ib/+/RjZh3mo3nr
Gy1tcq6PsJqCtpicFXMZ10PxM+4uV+LE+ZaJeOBJ8YagQayYNY6sXgu2uD92Cy7pAhs44oAXKdGf
EaABRP2mhVsC4f/xhgUQMLn2QgpERea2Dg1lP0Pgjj9cXMlZoeSpEuFe0ft+PshKGBEn+qpDNiqx
6gwuOC3wwxSTjceC9Rea9mA9UUDA5L0OQtMG6CcMcSaWaRpeeHHVns5b20vzLMEVDqHTDYJ1deAG
sK3Bn1dNLAbPt0yLR+2CTGi7cZG5XwL2Cngpquc0Ra8wh2j5S/66o4Yv/mDIKyVO+rtr5qgQOcl9
8gspabWoyxkLrgUPxy+D5o9C8sBJPBCLYiT9x0WsWjcxiiA1ZSmJC3iR5wvcSwLIHLVdl8qiwz7O
V7vVuunKKhFtEDlQHUbNma8OG9pnX6urJNFf92SgJUX3ZYxM991MXi3TfM4H4vqdp3buHQbHjISH
j+nQc/44Z4KJJyme7OzboFz958e63Tu6Y63M8RXHtHda/SAEEbKjYVcDA8BHwtKjsAMAMuVntCD7
LGyzs42mkXUGNAXwKJqOKXMT9I2caNOb/MPKiTAWEIe1Bf81164Vd7rEtGzX+7gYCfF63XMQpJLj
JdonGiaxyvRcdF4Sx3yvGXxTqJUgMSMQHnhgLAEoyW4b+hc6jxas/zc74GVXnAEWHHFzo6jIzW/U
B590+YLEEDnPNeqFeAcDxVD2UHtgRKSBrooGHYIn15+3x0CRBssXvN9ZRNj+KrFtkisHEDkhw6qi
5PZiBSpc4BpRh5XVa+0bkjuN3BVZR0O+MMgjEW/OXLBqtXEqBfSi9nmWNhgWZ9eJ3k45QHHdCpZP
bbggdJ0VXd7iK15vVXn1wloShPwtNfJnVckCk20MNXor+lD4lBft5ujAYWswb1OLkJNrQ/SziaI8
Su6f82PscoKNOly4DNGXGEPCSOTqZT5/bgqCtY5cDgIPQuPTxFnLk4mUXjZLJemFlumGoBSXc7RD
E7UtOz01FwqDcPqwAO/WOneTiJ1XBg39kAdqImLBjrajtVhYHsixLe8s0A4FQLZb08Y1mNHEGNbB
5IwiIhpC5/Na3saHJSGGdNXa5AHKyJ8rEac+hsUDi+gjN3WVc7qgIPnXRs2lGIjpRY3AtGuU1B1N
pzZkkfFASbAWe+iWffA3iwOG4ZgXQ1v6uSlhdEsYl5ZHxiaI+8JIWo4CZhLnOoLrJLiRY6mN75NL
/6erQfGfz++qDlCeGeVJFAYxcNkmmxzFjwADsfJ2Ys7L1bTnTcWbgq4i/25TukSpET0OuHesT/9R
YywT4P2VPiGnejjY3AUFNIHQ7cfrMQ4LE18UvPNqRF9zfT1NwxriuixzF11BOX9Asq3G489F/eZm
rWtMudDqOQnsA89He8VIOGL4cZ0kAgroCGi3DUU9lOEGpfAbtCdAFcF5VMWeDgYrEeRkFKdSZ/Rc
+zcdwHV7GJvGqUiw/1pcK5tBk0yRqOSd+JHSYIH4FKcGisnTEDBvLoSLBd+x0c9ddhrzhEQg9ZEa
dHkOvbwLoONlVY0xByR+/OQsREEAbx0EL0z8fLOUO1uvMhF2tVmQK7zwaR3/BK88od+hBoRkwFCw
sli+vEx83WhVqfsY6HH0qHiATBsbiD6kfs/jfxRRlSVRGCdGncVO6kicv5bB/tErUElnPwoYQZvr
RC2WE2kjHv9Ps7NT7AQPEtBISDfFIS3FUvEYXE5036VjU86UNpYZ4HyCgMUSZ4JCehhtxxLL84fW
fmi0P/wEMl46OYAlP3EyMQMQ6awqfGcZClGptAxS1YILdmDcmUI7aYbinkklleWngmENRWajA0Ov
LFaJkMDlEdDbi6Wu2S8hYCDT887CSfrM4MxDU7T7EMHapY81rewpozwafdVGBiaCm7KLDuU0xRlu
7vufsL4QScJc37bkx8yGKQt0l8B+GX1TMDfaCbsH43g027it6OcPpGi7JDkspqyYQqBeaYBn2jlt
elZtHMhfE5vRak24CyVTn093zv+vhCkpr3BlTRlZM4caC8p/Eu1FcXMAw8nJ+/MXxt4aHHBY3Lhh
/wEyvmY4fFXzuOaqmrzWJj9bkFca25y6NNgFDk2F9hYx1O7XDznaNhtFBbzZg+znZ0uPcEX8LlAR
oJ5a9dKuziGZJY4YQvEBBmOFFgiMb+sOFbiQo+ItMlRUb37C4Kbxp23fCgUYujx+Jtq1N3Mxm93G
VqJ7eZ9oIa1vp9LzV+6QYoefoAi8xgoWZ+a/cD3QJ6+Ki4tNibnizZrmxydvpKxULJ41+QZKODRW
G1P0hxk7MWDFeXS9Y3T3JBLfvDcUpe6QbVhrCv3bE9jNF4ICTCboaHao00OennWoUTN+ZxbqH0oQ
YDYw8yu+z5CigMT8fo2NANmOm49GrJdQyJIUD6MGouJrbpqP5RXmDeWjlnfrl31ZMqpEXBT7cTme
2xdQJ8M2Q/aiCjg+i3o2dJD2eD9HUeaRFPlu/HXNf4YiJb5MvvNQjkmHxhErmzQK0t7gu5tu7mPg
kOoR1ZPrl+JOsjKRrHnIJYwytwaeuoC+P3//skgp3+w5nlpLBxeYhETiRAnzMIXyFsYiRJFZVEGQ
a0uqLnjGF2RJNOf9aFhi6rr0xr1tWLo7vPatK38vZ5YZmNMYRsv8LANDDb1qzJc3PzACQr+FKk3k
2iFmfaNBFeFKAtCJyhX01SULVWyA8smECqxpALvWrjWMi4QKMc+Nag6C6qnUOkXKUAhfxkU84xYB
ee/RvufdchgcPV+QywlIozbdvZPUgAYwFRTx2O566CezD87tD8+wYReBcOyJgoFYQ9aBDxZHixyF
O933w6grKvAAPITa8Jg8NUwG/96sZvOmW13TO0W5j4lhhrYU8nM0QdBM76FkJJe4Jn5R8uNHlYiZ
aflsbqb5eXWqA0jQD1do5bVOPFTN6ypecs2o4zfU34iNnsaXfssvTl8Lu7q4D8nu130nq5XyVOJW
leGbeirpxpC2xPj+qLdrxrW0vtUMRjxo92+Iumw+3uywcpJ/fwHF2CWJKK5D36pBZFHX8Tis9SSu
Y8d7BNtsZASXoteE732oBfPySzE1Tbu7jAa4LoinO9j6JojhxYWpG/KRjLYfqzCxvvDPuZHrjweH
dc7Pjzqm77MFHIKG1lhEEa9yAfS5A7JBjHSe4kB3HBTy80H36Lf7WL8qVcrC3VJS4L/BkUo46Y65
3ag0ZF5vw17Rgosy92NO8kVAIGBLzrRqnFHu44YcWWQ5f4LXasNeI5Ym9qoMg/16Sqm+dYWcxC5V
q15bZVRFIrtvs2IQDZxuOKjBKOmkOp0Q03b8gPRWsam8KOd5fuUI/D0yZARwKRePR+B4s5ktWac4
dEvOSrYaCh62GVjWvC8od7cWjZCM4eW9vmsyNpm6MHwujhep0EN/30zzzxOF0BaF8Adc0xaiDPyy
j8FJZWkAtShGP4TVVxMpbqRBtRdVSsb56+egWC2EdB+xAaI2xryt720iX6ZGWq5asdndKp5OwuQf
7O4ZuFCFUtvfgmmzoJinDtNGDzvbgxw1nMvp73oUHpzYMkNU+VZKAZGEV+HDRj5S4pGTiAf9olom
1K4K5HTc7pcQOawrT7LJFeg+PuQ0m7XIFo+rGK1qAVf8atwfbhwgGHnSQNrth/zKStfVM7v9Lmlb
pbrFjBCGcmOc5K+H5BIs60Ov5WcPZEbo0I2l4khZ8St6Cnucp795fMj3WX08b9iInjLFrEIOM+pR
hm0EzKXIUMECUw17oYRP+LDJ69E9dhtvO3Wf1JNR0YfzFe1E/Qf5JMvqXOt1YGpPUnQfP8lCMUhM
suK+sB4MjZJcF3oYvUDr9jbNUBzcGl1CUdI5Kzrxn3o8y4OjlacN6deldn/uU9RhzM61lt+NhcQM
DYw5+IFk1QaFcVipo+8usYBWFK0quZKUlvz97Vfo+qjMAxKwLBA74VpO+bjoIIzsZk+M3NT1wm1g
pLafpJ3RJV0lKcfSuoJsKHqhwP/6aV4uvwTHAuHsEhCO1S6BgoWveekd8XMowZuzOUQWayG8GTMN
M5MrgKrC+0nG+FWOLNhwIE+Va1wqqrl+FupIPmFEEwzWetDuK1mf27PknGnm6/KmTSRz/YCBe9di
FmrFNwrRkjutD341FXymXxnK+1kMiiCMVoayx6zspkaJ17Tdki8R9iASbHMK1Cwr0T6Z2ejQDivM
mDeydT2OqsD5KYiEp84P2FV/z3dO+6+dckYPWYRo/saGfmgRSZ3Gdr3sYEA01oklLSz28dMw8J4G
omKWkA8hdX6sU6CyShq1F9JMHmm7gQod6Qjhv7UX4Ap7JwP0c0vyYuLZA2Bh9niSqgqMlmkNdhNm
t8cONCfs5bLb0c/vOG+6j/PzyR8B8BoYoVwKzR50qtRCjMl0vt0nZoc0DyD61mRvziU5IJITJL5a
VzQMCeJGrB0v7T5Fy0NK0z4lLDvkucHSGGH6q8QQY0U+oZM3lQrHS+pmfd5fX1Zh+Zr7Ppoa3iGM
La9pt7mn1dbf++gQyDtXwqyQgumTQTKzH6WQtBr0/mn/Fufmf4+wZ1MOhZ/49gNPHPvxpIbBAwtj
ZyKm520E3zE0P6une6P/PxtwJD20uJEWt8Ar8NdF1jAkDs79Fd2O6FiDHSnNpZuUyocBeZGRos9C
34UGkkeRJJJRn+bXi37gNhLD9TTbH2NsKIDfDsTBSJ9S+96IK/PewlzesCT0bBtKCilubTdKbMNi
yUaK7BjU8pVy6NC8qf254cGOWlc5R+TSGciwWbgvkwQoc74JTYmWO/2gKabxZh+OBI2pJoGkV2m8
LdCiqwcM+uIB2vXfKdsldNaULf9KIW1LE0gtnKcpCpyZWHvFhi9OUxS8l9fW8tG07RW7cUIt7/nC
bNOfEvWkMvE3ooXk865xQPU7kl1bMrt18wDJqhSm3MzBX2vJhuHN0oKwwuauL+CeVRp3BiAJMTWP
wIx53j/l0diODIqBSOlzi2X3Onjyb/7Uvwcw133lMj7fBPyweE8Lvxm/uviUeWxeMzxFoGM5GiZd
Uv7iZC4CQW+2bLDIOFwSd7NRKVSXbyGjYxeO0nHQ0tyCZPYAiTrG4b/2cW3v2FVgYJtZfem+qQ5s
HbN3ILQRAwLFWiOAo54aNEGcwbjgHcSf1LyJbKqXMzgexB/tI0QY6YELj/ah/FW3dhNQ7CZ+eD94
TJHWqXus6wyhWvxKGb6kca2/XuHiyu82GHpcbE19ajhykk4CvpOnruHVDiYqYs56Qbu+gnc4vL8H
PrngvjmhDOGAPy3499vKhziM29m2RlwsOub4I8E+jLiLUMa8B7u56gqKNDcYa+cjD9sOpuVIku2K
hXnkFvrOXS32Ca+9vkiDG5vP2tkQKSXxoCgTT91ZJTSwLZ2Hdg2xExgUbe6BJMotCkknwmNOty2u
76pGdofBgJq2xWvY/QRQtdoBfxDJo1JlYohyZIn2o4GNl3t+3BEFrbLHHDbPwuuWNOmi+vNLAfBm
OpDueDjs9hq7EgNxaCU0ztN1S9hIuqLnTm4TvW7fPsdVQXW8cPBRXCIpSflEWfU7DEyymh2c7Uz7
um18REn0hG0E4dRPz6t7SMNMO1FmUb3Vdo9ultCd+FZUkl7CeH2/8Ji3/Y/QKj10lD9pK2+NN1gR
1PJBvi5RWL2Gjq1R2QsOn8B8assH3KqWVHRSAS+fyOOWA8wDD7gFAowTYNPKBJKu0ee44v288zgy
vfd525rX7beWpxeZZ6Hdo+WSxDgAidsAfGOcASj0uaA56aK+wLMSAM2SWBjuhyl/KRNLMY+VZA3A
fxDN+4xLWSDUidWTD1B2n+m0hdYESEH7DE826lJG/lw+bIVK/mY9wgzQY/1k/UBURLCnKG6utGKq
PsOo8prVRBo1/Wsu+rAEErrFFikwyS2O0FCCWrL8U+BP46eLl9YX6Ag7r6kkeF8XsDOyeRA/e5EF
twx8ALvp8xselqIyAzjLLuK4dw8wPj9gZPlVD++a5C4atiwDFCRwELHm2RNrdxVKaLz+LLxjhd4K
c7QvPm9beJ7a8r8qh4Dc+d8wk4d32bh6Aqye4ajuEbV/NYHoVNYb1l/UrUiSvS+14ex0FWxAuRLJ
X9VzLNJdNY+em6zZ/qbhWCdvjo3fzV4Ki91EV5jTiEm2Wey0sz/Y66MbDe0UQ/+LAghe4ORk73gL
QcJAWeTxdq4LaHDCVM9lPelWp0mBcJb56fdegs+9IEXZY0RbxKzsXq3x6SWm+iX5xF4Exu6oQNT9
YiLXWFp23UUqHSsu7A4q+YN9bIfrI+Wv6ijHonYSfPK0dYw8Rf+CSTGDIFtoOvepbpGJP7ZCQnsP
HevgILGSqttBW10+t7rP2BtdTpuA7CIVleQXR5ePcz2swjcvgaEXxvgSFx50hLYGXiRO8t7FseLF
20dIJRjVIPfocdlWFmPylJOgNsBtXjX5Ozazl7xr6VKcrfWnzOpRl0lj/lToq4+4Q1u/RcM+PfoC
E3OI6QfaGcmHd/BN3Kiep5a9+S5r6wO9VGFqHJOA8yRVLBwlg0sJbUDh/lSUixpW8fS344a9u5PT
LrA5ADy2YuGcZjX6qX2dMFrY0GTkDhs6RM13xi6D4PVAZZRCfPiEoxu7NVyqY9vVCSG0Iqc76lcG
TCzZDSAvjwvRgMK1vpypf3qQQTUTruqvT86MoKyKaRsTPxYGzE1uJ2q5QZ2f3UCaNqLVpPWJGPfo
yXo7l88TxsuaHruAyvdgHQMvCt0kJM1fJVjBRH0aKgsTCu38rosUNyz40nEXkEeGfmzuvMAsl0FB
EsNwl4vdSbBRhnlkRj/gd1iZYqM0K7ul5i9gG9UdQqEVieOsFJ+0PmgUzHVh8JUN4S/N746dCbr/
Qom25jYYNkf5PyWgx2eaz0lBdyo8rd8gBPk1WRGbMGfb3pLWcQFr6hHdKRbwYZn8uc8H5Z92j5Uq
3wkW0VOhQ6Oynv4lbvJUXazKrndbDTHHEj/e4VYLZydFq/jFK6tbQDmhUE/+fIZnbVWMrmJQ8TNY
/SVzruwGB02YGstN9VlkpY3FvUEMmPS8/ZVMbF0+FGBpc96IMB3EsFR6ulRusttRuO3Y/Gs3JAsE
6cNqU3Cc95K7O5TCnsreU0/aYC5yI8bIJAb8oijDUF8KAqxUvmep6O/qGzL4JhmFf4AmovlN2JjK
utp6lAZTAZAL1SyJAwcgatbNQCLVYSdTPRmGLqTql+XqCpVQj8dkVWtXyDKJakGx32Ilohi67wP3
IdbToQgvr6ct+Lirhw/F5Fv2l7oUlk4sT6Z4gMcaABY989nBOI/GZZPIXNtLA06kPl4WA9wNHWHu
bxrcz3kFjTwoqAzXyvsnoctLDNFOzm5uURrweMSomFqj3PZkUvmxGEGgaDd2nXYn8csfleQugA1U
TtRcSiGpQ4m2QGlDMpJbnP2VKPF0kk3YNDSujv/bNP+thG03KELZI1v3ebjskZEbjY4yLG64OMK9
ynIrPMtKU2pAwbJ9xVQSQ231KBMQ3rBfToSVDyr5etySbNtEchA/lThPotwNmY9qE43ALT2y4PRo
DFZSokImJe+wNtzqjoGVBX9Qg/7aXkBUIIRBIksUZ+8jVkgqAOwutnDxWrRPxjh6Dinv/PdT2rC4
Edw/7IQA6c17mJDz4G1UFXki2Ul4Le75jZU9yBDc/DexD/cYM9o5uS0skilRcmb1+o0UxoB4h8gi
3CyL4eV8js6Oy+vxcbhGBDigiHcdxbK5Vg/dzpSlBv8ToKnMRmYpX3q9QoJXTpRBIt1Vrp2odHYn
Cdn44NaR6vpyoOMfTxygfn2h5hYKu/eH6P1OgMZUrxMR47naUnkYGhoomKgEFW8D835GbT5De5QM
Yc2WyDOXLPaiZMOQeWpvQ1VUyFrRdZjfR3wW/lihrKd65rBNz8kmZPbRUVtEzKz6+jH7EzF3U/4l
HFAY/TuI98qlGW9P/2pQ+UBdu//t23teXPeruPfdQPYa/JEeye+iuQgLLFLj8Pa9lw/4nm2gMnba
iHjGM0NZjV0igdyeR0ZGh+MCP/cw4KOJxD517GsjBOI3O9QMNMAPybpg0pJadsRHo1w//e0wJDLl
4sZd0xE83n3qTc785SbjLM4DBYQ+C3uDZb80+oFxBB4D53gQSpSFSsc/HUmWUoKPFwskpmoV+SKH
3YdBkJH58I/cP02xOgNi625ASo5EbBRzaUf9rCm5fgtaRslIDEwbbl3nYfPFcjdQyzzT0Nz/+PYl
jCtFdWk0MgmdvLQ/JwrwyBGIOKxPqrFzhyL65GASkFxRwK+ohIHeIHHxNTAC5s07Hbicy5lHco7V
mbihMNHf10iKUbAz29+GNn40H2PsUd3Ounuzh6mIz3XriEgE+3bR+T62RqVIKYG4fxY3DGeGcADN
t3HYH2FHocBKz+1Uq564SU8gm/BpuScUqGNxZGvatIWAqmyucIc5lEY5mKIHXT/iz2325uIvbHzF
9eDWdnJQu7/0lcraP8zemk+Iu59oyJcHg3rGc7KN+o9ceRYijt2IZWXjTS85RT7VUCn3HwWdp6WP
3Lk3mPLdTVvVF75i0u/ghx14qxmtj2rVtz30yapZdAy7nmVs09EOoS11OqdSa0VQxZ+gFW0SFz9/
vyKZzNItHkyBf4tNEPZv0wQI+FPC7OSFuBElQ8oTbuKwqenMEpAXjBlarMRTrMOOuBeirxJ1vN5t
2hug4ZCl5IoMvSEPQqgm5uOg0o89Pxs2dZ9jMAZ5aPo3o9MUMuK3SG4sdhu8A9svpDim0w12D9TH
YfxznIA4XDwvkZb84t2Z6ioyKIMLkur4OsjvmY1b40SAXloOIAgHtDorAZu/VfEY9t6STyC7F7f4
/UhZSxDJnUWOR4u9getY5sP7xw93ODDPWqEhL7UTOtI+e6e1dDNz4PAmi+Ti1zmKXiRw3E3KKojd
1yCHBG6ik/NoUg/+H+JndVXp3C1NvDYHvVRVCNzolsgRmmeft6Hzf9ASsF4hu+iGBsjdeekSBWHi
SuciRHpqLeGE5QAsG2Q5qypS/mTNgKIGDVrVZQXol7aoqA0TXHOJ6xXwuI1PNhvfE2hWjQZG9S1F
FeDdahPXYX+evZOG8cGy/C5OsnC+CbhH12NpWEaPZ+ES8Z+EJnmzDhJi6BS62pSg0jKi8hsnI4Wa
gU+5giFtq0x9OjNbxHzgo/AAur6LWpjHicw+GR4QC+qsFqsGwbO65PavNQnJZUZn1zs8rQCS0ffa
+nvwmSiqUpGxO1PcyqGsnJbIhToLQ5PBev1yeYN33d5aMgKSX8IBdQjvT1NLh3YBiYTEpV+61rwu
f79i6VnPE2xpK5k5phVNBoxaBRuuFbwYbfn+2U1jgSmWY/qkCe7g+FbJDyTh9t8raC1yhuZdmlct
j6LufXU2IrStDyszx0Smm7JQlPx/rgc77uOb30GAm2OhYvSPP8aFmM6psBRtdiN0Yh0be3uR3IBf
owdRolp8MFEM6xUpsOgg5GefxZoQdJ3Pj6Rjhi1KPJpJfgEqjAGxEDQn3WbulkUh/CP+8/qnr+hP
lnFhB5pHegupuywen28eThlU26M/9J4yHP4520hbPPSfT1F1TgtAVreJjC05/OTzUJewvnQgxfIl
E0IduqJw6cnMFmX2nCLVmTrp9MjaaVGVlm8dODi08LU+eH/eogWmL2rjV2f+CL57GhssS8n6SJf4
+dGKzWwdKjcrdh+r8lH9K3L2buvfdAqtzYP/8kM2ZJyrbr5aLjRygvWqB09oIlAWK79+Da8bx26y
0+fyqe8b2OHAWwAu0c0gckuELuBkBZqHz87YCx7M/s/sOxqH0NlJ/efoAKtBaX67pLrRVhdZHbDt
fGcKHqAy1CSCcg+Gc77AX4jRaijCvXYK1u4trX9DHs7anXh5gQcN6T8uuZIbqaFJSAy0HgiaLGRv
JbKLJuhMRubSWLtAthu2k45xLMxgBuVkcvyljjlOrNKLKMN3a1HJVJptxfwAoaMSm80kMTHRhc+M
Cpt0grgUfQEupbJweMVcYbgztJvqP+dqT49X6sWW4CeSWIH321bbbMXkw1RoN7MdPrluxNcY4wrd
+762wTvNrSD1EusDD+QRU+C5SQDl1N7WB1sInTDcMJ1+l8dsDC3J6C7JnX4yFayE8LLM30syOB+o
0dj5xT8FfUFKe/BWnNUkrm3YVTbND0uyA2Apn4cM/sIj+eY3TlNb2NKKN/xvcW8eF2UyZF9+6CJ+
1QFF1ZSrIcSCil6jBGx3mkNQXX/dJ1r1qaB7/W7UkmEMBIEqooaTkZ9xHBxBFYv2+GLPEPkvlVqK
mgH+XsIHGnBYPJNusyGsS4RK66DlXDV8dD+xqBQf8tscPBpWfW/bKL5CZd20Usfw4KOZ9A/uDs6Y
RgMQf/tKODgHHzncp4PTsIo4Ktsxw51oAzJ/cGIBYXfG66WoowjUIm/0+P3NlT7IGYwmVx/9CNa8
UDMyvc96JTk9cVcEKiKN//s+MJ7kd4Oe4gQi6s6jDw1GoJKfQIHbibq2X6QKeU878MF/zDK17DMd
C9nK+iigt5aYltzci5lA9XIMJ0S8SzyjT6FN0z7hLQVePeP5yS9VwepCpB0wd1v/alGuaWSyPDiQ
mbNg0wCLARm6xgPulPwn1cYUS9ZV5J3r72/8gba6deOMzpzyWHg+h+myB48mnjIfTf8CKd+KDle/
+5xNC4r5T/nyaCigDB6B92T98KhRk9Vy852BGwlocohy9QAfK/D2aNp8ehYikDzIpGA6uJKD79fq
c631oRwiEc2cqt8B81nKJNWW+Lk4pGFQc9qgXVQ32nKswDZcWbbvMFUQUapDQ/4YqGDL6B9Afaqk
yJkVpOgVaiTxyPzHdNzJZzLd9xDbMhu6AOh6g585uGTVs2zInzA6GkDFz6ik35Oo1AJ8rICQUQVl
PJSddXxPakuWBmyZ5b7Rb9qZW1NhGfHkZWD4sfb/8wsrVFaz6SmXiWzWt+ZN78i/PIoJ8mXMmxsn
h87s+W1IuSB+wRcudhfNmdAVHlTKHkOsvEJExk5OZ8DtGiyRdcoqcO4g305lM76de/vO6VbXQqNZ
Tlr9cYtrUE0snTDqS21CId3rJp/dqTJhkumaPtZjQgmfVj0QdFGvhp4hI+0ijFxmPFZHa/ZAoAu+
TK/Yw4Qx6cJBUV+sN/2wXQ96AG9BoOpEuy18BBz3Qla6t0qwRu/qBcbIzBk53LlBYkdfKMhfB/Hy
R27UPOS1lMML6LNr6lC9OMqvF/w23m5weuqu/r/GfsdKoonFXFawEKaqGKexnaN+aIHfdB5k5c+y
psfrC4TM/Thv4XBq20q/CxUjilF0k427UVMtf75Eu4q+rjDix3bZcL6R2/3QZ6ok1OTcKH31fhxE
y7e0opU0ocThdx+gHSsg4/yRKMhd/YVr89rq2YKR04wp8FZx94JnVY9BUqj9XLniaMJvJpAtSIT/
7BrjBe680XqNGdYmvldxOW5VAS8mVERw3grVn77K8Ath2nNl9gpHDudj/RMt+6kIPsznwSK3JIO2
tRRYEa8mwRdk7zh9CmhBsv66Q43KMZeCB5ole8qDrSwZaSFc/kc7lfhjVQ+VRNvwAifWY56DS5nm
bR8aoOgp31gPGXv18JObSb2xb2ObiBsRZArqfp7aDtKgCX4Ue+jWxfsn/kIdop9S/5NpPq3Lx3wQ
yPhrG4YExr+VLCca2PsmN/2y6mRBc+LcO5ZzQAXNOI8DJRjkTpkYqSlfxV9uoC37f02vIeqaJAKy
OnVrPk5z/VPIrdm38RZFNKmrbRVhJTvLUz5E54CI49rM5z0R7HPQBQXu/9UVxWJnxniLLR9ZsO39
xwPuM6nPgXnLuJkn/FAb3Eod87ulIsmnOExw1LCF3R2uW9TrNltbpF9HZfw1JEIj/mIovajVHgyB
F9iu0n35H4xjiBmIuCQWmRZ85D5C/luMfr37sZmIqs+Cafq8lP3iW5iMCH1O1ZpWWcodDxCnhYGJ
guuwc8xm0E1N9hB21vF5Ad7zpA75FSkGt1Ms4kk0mt5dv7Y0rT4iFpOHZuXncaUWTM2lyfJzsuAN
kKyYHXUf4dazdE5qnpnrX6Rxbi7jgr2jy8i/27NmEsWWiTAYowZ5kiCwi8RvNPP6rpnHgAHr6RG9
r6jWcv83Gyl6rCXbpOYzEiua2kWeEOyGXiGJLAaSZvnHJKk8h/RWin0pLj4ZUqQc521UhtWRQJM7
ug5o+/wPOMi4PQOWF9aI1kukLSR/Tk8iAs//xJbsHj9XW3IPPOVtJ6OopxTR+Gc0DNZ8e+RUSEXQ
aPmEcXHXtviOABxXBD89o6pkOM/BFgfq3DUYxXryvfesnwdAtgpaxwGRbcu3zYtC0hK0LoMrVrFN
OVyKO5VItplLtbZexmn+3Lkda4POQgDaeRFKOBQqvD+kzD/OqRu27f0yb32YySXmgfEmrtrYQ1Ul
Zkj14nfrwm2pFJQc9scH41vFvQ6LXrzz39+VbotxGTeG/gPJKImvRaSwOUQ19lrXLtbEyi3xO/KW
q0k2+8hjoxwCrgdtAWRSL2CU8nQEqmq6jsHbyFsZxRp13sntVmIwktNHCtAJqRUPrSaQglBDF2fi
Ux906pB3kdiBbEwL0KM5Vwg6nbL+guiCAyXPUzOmZHKgHP65xmDeI6AUtxLRNeAu68LIBAeryPVU
2kqHmvs6tS46zan9F/Vjh1L9JK2ecSP/fw05F5LO22JtVlw+gIMiVQPKLLhJyaK/FA4RbUD5udHL
V5mkwqjM111+Cr4KqKSgIprvhg2OXD4iDxQqa13IsyrpraGlKz8yripGhCzNI+/0NKLPaVjzYTxb
h6Zopa8TXRRaYS93lza0s6IlIt1tISAGQb/SeX0569kNNzwibVnPT3WBkb0bSYQ10bCEVtryDa7U
gmDiDc2ikMxiJXtLcnMm7LAt5kNvjiMpFZPAkLf89cziQKVmHUh+2LOo5q+TL9FLQ73Fs0ArT2cH
bploQHpSSqtDCAW65wkUsAkzWCYgbu90vD/IT+Nde+xXXnPpgvjGkAO5IpGpGVyTGQceoYvnQuhD
7Y1q6skbWez3e4UOMqi+5uvXA41dGuecPpnv3QlgVD4qgl87/T4LcTTGrZqFj/9kEtSraMqAJtsr
2SOUW6PoaoHkuPTxGJefUeuqlhGO6WGrgoHFh7kQmF5NecUCaeIGi4s2seY9b88xm2HR5lMXFFwS
31lLMPhI3CKkCpjhUMnwitOE03/srEQSAGX5kGFb32lJ1NKjdiZLAgg79XUY59+AtCYrsAonYS7M
5BKQpnJuzJFeGNBT+rhOKZy7TiMPYRWlT8Eu70Ksc/0qjN6Pn4ER1gRUL2Ni1TlUsaAthLqKfuVR
X3e2zFtqPEfKoa+KnRuIbdAemlKXLMgjdHzUsBMcPg+o2ModfLpvVYbONMSOo0BELG5qt6pb9fRk
NUQVWZLLk2uJQ61Utb3ko6UgxQMDihpevr6xo7BhbGtWyqThw6rbiVLYhFugwxYvGFD5W9dGBQgH
eKe47QBJwvFHLJEXh3mK1VFiknUqo6Cxwmi4g2/q8VZtOIfO4YuL8A/arngZxE76LBJUwAm2OvYN
1HvaYjO+HAFP5U07TseQIQfre4qp9kEcjx0W2zECm+Dk8HJXVr3vHvwnNtTouGgI1cJXx5lV0Nom
fpC1Xvl0RjlubJxFUbA7tMBjqUNVctYScj0fKm+f6rBtrfi8cBF4dGTgqeOrSRtYtuM+Sk3H4XfY
hZqZTPhQ2OIMJEMDo4bQm6MRTc8ay5x610zjx02TpFFVPBmkRy4Y8UBDQf2tEeRu4y8KHYNN9PNw
hAEFUFK0g5MgpEr94NU+Yet5qk6hsqalk3eMO9EVmYm5h5FaG86CFrRnLew8OOBDoQvQ0tgkgI81
ydyhKJawigvkwlCJZKKFsAjym/6lYhcHYSZvqT5jwdkdhcMyCG2vmtuUR/OSeJPQYbagVG9zB8po
b2jcpPO1kQRFe1u5C0jEOLzOW7EDOKHydAZD79Tubs0nVBDB+N5Jz5GqHpiHdaOxCjvkmR2nq/eN
8RRm/BHsiTYqtesjvW95KbNJcanWM0anAeI1SEUTWOXVDUnj9Mz+Gf+C6DiHBxr8qM1GFMNvFmZv
I8SbCXkrKp7dgabNbSktE1GhjSrMB6SaeCHtlyMfAc+Ja+WMMLVrEFGmWfsZ9MK99aNavaU1qVQY
GSO3h643r7m5eHstJbRfQesYUEOWEcMmapKvKhYfNZMXiiyhxzLPNWX50xkogeTac33lPhaTq/nw
Bf5KLba7jayzLO5yqnqeTVPx4inHELLrDEopn5kCiPOLYpWQJRvcAJ4oZeqh8TuUvM+WysZX/gMq
YmT184uQL8ys53MpLBgizeKObS/zNsqHK7wEtzjpggvacWcpR1W9pNhNGO6ooFtL37+MMFu+bwGm
IsxiPU7CUqHa15Rl+/rwPOVeReuEWSXwXI2DJWxLqP3nHHYMDdv/0jbDqq+pzdLHGDKIFSRJ/Xet
x4aHJJU5cDJlTkReNAijUaPM9Fp9lf1QdfhLrpTzSgvQhyjBBGWWSDM592UcRvFn0ujc3qXZgxsd
EHECBmYrcWDbwStgYpk0n7io5nSQ+VSeClk063MMRD9p5X/v8NrWINtDJkBd1BoBynpHNc0LjGLz
VDiIW8t1hR2AC/t+Ya0QwiN8DziHODFcJaPZWZc0Z8KP/q9S86iD9H3Jg6dZlVGc0J4GsSNif7y1
mkaQh7DIxBWpcMmH6ilhAsAO9qiu9ymI1NOUN0IpAFF3V5QA83c0xasYbf8qOCr+EU2OHUBTbaL3
YtSSYZuPNPYgXG972Zrzfi9iZ7II5VjLaVEGtceJvLGBCMQ2sBSikRAX8YKtiL5EEZLpfPX/q9kx
Zg3LxaCzx7jp3+mYvLdVIp7r8WZkSmpEdHuGBxwuh1TIr+jPAW0PhUlB2QghzguKl91rJchxmYOM
BOh+/3N/Mk+xjj12SQ5Nm8plyyA47TjNbOVlsr7os91Gr8KaLApAr0KX0FbZwKLZ90C8kdCV5l3s
UHvFUU4jwC9riNEo2lfoXaMtYj+8I9YhS4pwjP35InsvqSZPMK/PdDs02I8xW1/+v56/jb/6lDe3
CBk1rUeffhh284hrtlRHZHNbYaFWPq62Yub1la6t04CDVhjK3Js1eeQ+MomEElbLFN5rEZyJX0Rl
jTNK7/vWxwpcr3kUA7riDOl8AN0SpNPSet57URGt2z4QN7XKDx7oT9LAdijZRMZg6rQXL0pq1Co8
lEs6Gl9SdvZpRKxr+0ChiIR7YUMAWPOJBTGcc7fvFoWRT00M/XWQ+rEJjgtYkp81DOmv2i06y7zf
ogfHAHwqEy0FRUh/cWdFG9ucORIr8RUWVdvNlHAh8exGRvXJ5m6E0sh+BrvEq3okfdZwkxY/jTEg
Z+LztkLcx8Mm63+uRR6rmaumy0SiU0/H//Gq2W8Lglvg/z3VLzniUQVjvhpJ+7SB2XWCPf1YfriF
+45Idp+0l03+2PDq92SHG7XMLDeEB5COxbEq+sQJNAJaWAznbZO3P2V1tMWjUM/rrJ8GgbbBFcHZ
qSSeKR7lMzs5+DM4ni/RAE6tNv0XmBh4oPmUAtCDlmXYfyQ9/aN+j/KqPYt7dCVKLxW7Lc+EXItY
g5zCgrU8Wzctmj3P/tMHFz2yYGsVN0KUqv902kKxk79vUE2sPBkOL/MQq3WzGKyZgnJisJWuWAcl
xx2KPoAdCOEVPb8RQisLASsl04ypu66yyypuxrSvlEKOB+W6/NxcoyQQdvBgQ1/qkxeRFYCnjCMi
LRiM/WAoY6rFNC36ELLehvZAyGxDlHmUIZMonf0tb2ifisAUTSacdvJfOHgVYDeY4fu4x+WECC/Q
z7TC4VaEDbHz5CvvqRL/b3k5TYWTa/NiSkxPV7OjDjVI6IXA16mwmbXMwERQFvn86Seq/68qd+pY
5+dtimOSb+MI3jKv1MM5aaK1rH5/SlcMuFRxY4LoY0OqlxFVcpYxC19vmUgRmONUOoB6wrPnyjaF
FgAZncRhyiM22E0ZxdIB7lAuUS9XjEEFpjpog9mSmNxw2R2Tk28yoquO+Tk1gMwQNU6KQ7tDrzxh
+aeNR9ERHxcetDkgWplpg2u+ImzHczEK0qV5PmimmeMv9euhndTBs8dYCKL7huo93jWdVltGR+iS
4dESNrJ46Aw+eZjP+gIw9Fx48XBMF8s/g48x2LoUasnjExTwS/m8hFeUnG69asRuO1i5gHNzxSUj
hY3zBqAbIg622BQ35mPtYpj/u0oAhJsb3lttZ9Mb8unLfIu6nUlaKHrnuqf9bow2WyvMO+kyhVR6
RpJoGBJ31twFLaxaT1CfvXIJzoPZtBHhI3V7HKXu+oIXaI/sGPGCPmDWyaPKAn3yJcr7K9tsegCQ
bCamlapgCxVaPpLVbnOZP8fCOPgi/SqnbmMHB8ufistQuMZk13dPx+I/qvVKjd7Vaj4DlBNCTmk6
8t+nsFxStSg8j4ZciPPF92DNYefJ1NUkWgZMlJFFBunE930jOPc5e9d+ZZbzdtRByrlrrzzMprUX
FackGx0iPYcAmr3zoxyKPEkYqxAMCPQXc9HYfMRAprPwX1zhAH3J7Elrd/Kpddp1Y7DQFWwi0gwa
u+1ufKdLhOOyuxfMgxH4y9s43lFqa+bt30gshBTvBj57Y7T3tJJhjYhd28NFIfB9WvAWPHT35Qtx
g3sLmVhLgETlZ5BzXCMffsK35CoPj1cz8F0CTgejFUQfIILXvfwnQ03k7Xux2SlGJuAvj6r+Sngo
Kv8tWh3XmNulu5oFU5By62fTRzeaeHuUVSGsspk2/Io3VroakG+ZOJjkvZoN0HMICSXw9jrDOTco
4tLZfnBG2/6IpkKys6iJxOLMB34jcGWyB5q6ZwEHoZLVIpo0tgWzaTXlLITxdv/iLrzUCKMoIhBK
OpgEKdb9xYVVM/FUX4KAG/xvo/PxGVeu2Y3Ejxrh3Dz40nXv+96tZpz9KjgEBS5qvYoOn228AV/t
DicaZM5v5W3dypXPYGH0zVvCqe7a0tUBMrVnf7cXgkr5dHcGToGL5Od62hIRRZBlHUwPcL03jVDa
zJxqMmHIl2NABth0PdKlnvrzIBAd0U5J0gVncajpPwNXox0Qr+jwmQDxSVrzKpAWgJMUvjVJErCR
Bkd4yFPlGDiqAsG38rrBeTk6UZKrd3yo6UlSXDfvaUl2ezjBt2bD0k/h76rnVHL92sAOTGCvqTTM
fkGU/MwcSh+afZhhoC76bANF//1LZ0DG/nunCzfdBDkiPLw60/iPuj7X0ZZJFjuxijj/upssb5HP
hO90uc3CntD6fwTkPCZDHTMIkvWiHD06oqHX0Dh/cRAZxNPBeqwo7J3zi6+Ld10M+mrM6yv2Tl35
ayR53KGchI8+HlKCh7yG+553cTvFAclOtED1JOZLO0KMAwB7ZKemMSPym4eOJM0qmOIUEA5JpEG0
Hj1h2S7Tn8dICwwjIOiADqvUdJytpPPTJrIePodTmXLODLcZnSTCkDgOoDOSm9k5/HTl7vtiwI7S
/fu2/3UXY6fGYwu1X2Gg5nYlIGAL2E+KiHYtlDoiZyFxBL4z43JkG+QCgrDLz6zTagFCF99EoeGs
SvZ2u3daU0dQvYYUErOvgyPlTngZW+Q0oR7ckQqG0d79nGnxcKu3SgnLzY78WfvX4CRrK5d4eDTj
MLkfBpcdXCGsNsctKbSJEpkgr29nOmxI76U39Im/C12BGQ8zngjSe6r2e7JXDPTk5RIY38D8k3Rs
7ZptzuD+Ea9bY7sMZW8PWGgKs0sYmW3oAjClxYeLy9MaF0IxDmxNGG5BMM8S+jd1WujBLB4+dpSz
wEDcfTpmgpVrXkWEXHMKOo6HQcc2mpor4zBavGGQhoM+BukjyBmc1cH37zaqYrJukE6nBokme91J
xgvybmWWLZ7+8bZj2JtDRzxWaqFtZ3KRXAaqkI8KP23925v+aaboYjcvbor3Mr1h1JhJjLoHjl4X
7TcxY/34/5POhiFSvBkx94fTMqhUL+0h2nP88yUfUCjoPXY0/sAHfm2votd5q7FIlv9+rEwAUCPP
Hn98ZpthIbVledypS5j4mCbK0ekLbKNZgD/mGzmHjZw1lqDCv737P1lfoYSqQ/9cywfaixQvl31F
+s/O2N3S0cxvGn3ViVzZcxZXc8BSCweDaS0coPVUvwNEkWOw7VLiZ92L8R5dZAL3SvK8qx0BX4px
MVzjl5KpjUVUoa0YTE34LJO05K1Wamfwdp55EVNqtPxtTNCxLz2ycNQpr4De2SemsqqIZ5CE9rvZ
5q5rZ/wKCvV5pyXS4MuNIiUvhc7xooW5prLhsPBz5vwpELNphDNIjh7xnDAuunAqbY25JxFf59+z
8/WXylrL0VvGYWQlMjR5H+7kfBRFyIawTnZ5EKl/EWeabRJaiM1jYdzHHZDnq7HcV3vBTKHh4xv7
fxWCMhk9c90khglhhgRofcl/2ZZC4d8J0qpsoj0OeoBI//6koOepn1n6eCSW/krWhaNxugHR2zXV
WvrKoWuGWCgZ30MVUsIp4+K2pamRT6NmwWhTekABK8qUG+eh5g3jgVRrbql8yrN4SQ3LQeTRck6Q
0y650bXKQnyUY8/pZzoLlVkqlD30690LDdnKymxUv4XKYOqFtZEqb0ESNL7SBsR66g76aFB5BrJo
C5Lxfg3A6FVLV1ydKpkHx+nG6E6DdIEeqEcDb533KyYEOltP3Pn5jE4Eyr/evC61VYd+sr+93zxT
iSzvdy6jEm5r29mQ9acKTgiZMBYKTkFuGCjaRp5ZAsR8/icofZVjHohvZbh3FyuaMXFmtP4eOQFQ
quVY4niiT+RGIwbhVbYzjNEfniadKPBkWHzJ0BN5g8U4kH4Nwfrelsb2Qkn/4PN+n5TqvEG+z+ah
cSrhWz7idEs9XIoSvPu5gA8iJgSJ3qw1++6oLVCKMa0xmBfL/81Das4ySlNkoFQzKuJBxLHc5XFm
UdHZ8zGUkI894pbQBzemw4HtolV5IiByI/1hQMxvoTZ5BlZ+umlHst10YoYkRUhjnzkSrx8Qve6P
IQb8Cc+pAQGAd7IQCbQTfJlx0EJ33djK634zHlCpRCRerSupnvEFDXNz26gqlx2aAah8h29mEU6M
FM60cBK81hodM0NyhWN3h4PyVESmyYXde/4x1G/cGs5MC5DV7dZHhsM8AKDovO3pRtSBCccqgn5h
nNX9jgInxC1vQm9y/sP3rAHMTfHIQWq+heM32U6hrUUd4LZw8vf97XmRjqSr6JT9+SBmk14esRZy
LzRa+n4UOD2dcc+RAa/qgU9orY4/XsWpUm57gbmb4pC11hp01qi0WGidntu/8AsApRsKVexNcTU6
t/YJIU0aD4lX3UNTGvhoHNqG7ljGP020kRvfbruOoI7JOV3YcKHhvt8Iwn9YDqlAQoy8OKvzkNap
Qffoj7CRdFLHRS0+TwDWgGupvXDlKOo8dRBoYd8H1pI4OY5ZOv613FqLJGM/9usK4jK6xMxa0dLu
vtzht8su39aoFuUjXWiGCy4Rtlo789qGsqTaDs6M9OCKZeI5ofW9FTK36RbeM7JeY4wSuNih2iWi
/TQqcrMXXAjiCEIGM8NmVlpqzExjLI20LPbKAwy6KnJwAnJv4QS2T8zWO38hgk61/dAEqdGp9vtq
pOZ4AbF2fRGI6VsHYagtTss5KoeBeggLaCYCLrMZCfjM8+o4mjJtwmlYsR74khRFRkUUp86bFWNt
qWV0J6hX+pRQ2lTJiPeHoxK9tNmqvnBtRxylLJy0Q9n7xqkLrng6wBjwgrHVpmeYT0VWQrTKfCKY
+Zqutv+TQ5IzAGTbRYaqJDjvZpTR+u41nzcmwm2C3oMYEyysvaM1sOvFYSeskTflZUOd5fV/Jcc3
Bl7dcBnkuTROE5QtFzgWBdjCJhOh+ju388FfHRQ0KxJ1T6L1WC18b37tzmYVgRHtnvZRq+CWOyO8
L78dRTRJR87w/nDehl4qJjCZToMGe+cBGNTQbhlDevk3GbXas5nqjgCE0ooMvQYQsWPgLlnko5xV
TtR/4Zzu+yL1e23OFpx1MC2IFkwzLqc5TPdI6Z+kddHQZD7bB0lwvG6JgCyTBQeCiD64fnaSI/CS
An7ijXqq+M+S/8qe+9aab30UxRQmCQVOW837XNCjy8wuMmj5+NSgDh9GT0+xTGNxOanmuncqcxEp
3NGPfgf08XlbjcqnikufB1VNQA+NtIXAuSDoSgnn5jL1AcfqmgRClLD9nXYa+sWHDvhjPoqW5x4L
h3Rvf2JJslAeT6NBYH1nX8Y+0PcCz27210aY3fJvS3+NP+QxEs7/ZXIhHrbPW2vHKgQitYg2xdYo
WMXnDN8xwRk8rwgY7WJDVk9lKAW9uuk/vp0fmHj1mfbFxpwE+bt26WF+67XWDR9F5aZ0rzVlBLKU
2eiqpzY22LPGcCm7RAZCoXFcjkv5y8S+Id8ADTBQRz04Fyq31H/Mf1xYIpLk8O/rfnk+m8MI5DHx
oZUFajI4CEQfgAg/bAuiFcrgFoYwC1Pz7k/p1naQnKiYYdlHkn6EIgkiCmQuvuod2vQum8MK7ZRm
W9FVT4I12HzVDryJ/Ojrq1ye9M/9kwAN7B73HEEkMJhjNohlvAHFCqzSK+rRwgTXkc7lhg8DBX1G
sZO50pTn9P4GnguXezU1zyUhMdQnbJl3X44D9HHJTwxpV0B6sRGDDHpWHFKn0PkflJT1ptGo2+Gf
6jZQ6e6GcBOgxVTKkzanIZXwoxR4kL0qdyc0y2n2y/yhmt51Yv4KDm9V5kpTsGAY45okR2rYbCea
YtccodyeufEy7uOcv2LJslm9J5iamAqymL896LdBVKRlCyeqSjrw5x4GGMtIKVpp/p2qJnh4uEFC
4MRXWJDuIe9ZHW+zZMxAKitFqIx/dN0pT4Vc5syUvWtf/QsQ6tljqeVBQ2KcXLXeL+xdnRP7PDTF
nxhOcQzoWaIwobgz6kGR5cgQDc5M3Z5PmgwAkLznfdzcfw7e42ppkiVXMVDgfAU/WWetZ0vXNubU
yUtNClWMB0zvOqmL2rQCczwoBtUx0cPlTBf73I8WKopyxjgtYyhJDHpS/uV6DrTVL6moNp78ns0W
PFj7kYQHZEWbnndYa4j1GXXqXgX6UsadrPPzMse9lnqrtWAxF43otZa32iu6ZlwLP+RVtj7uxBpP
LEKtLTTjDDMhtJHTrkw+9Vsb6cfHhrVWta46xPHITvlN5PoaFeOgkMTBJGRkpnnZsLvEARX3MROl
T6M/iH6RYZmZEUiDdoG6E9ipsjkvQHhpAZMuQKmHi8jwY0kDOBup2Iy4QZjb100TMiSCLsBStcs2
zXChjYEsk8Xpvc8Jhsq251dGx06VfcbwSonpuTQT2MPH8cwvu0zu0Xn648+3CtLPqD514Jf5n+YX
8rrOlRpFCb838v/4xAWIGwuPX9LK4vrUGSwaSWmTEHXTj8EDeJzxNJaIMizA5nnP5ecMMcmsXlPs
Y0lpX2jyL0howsN3ORFRQBSF4JH2sYoNMfCDJ8qllTxfn9W/l2PMOX3XcASw/XAKqXAxrlpvbUTd
kflC0xPlVdpH1SlNltJYBX+e3Lh59qDM3TqVYVRmDiZsJ5VQ00f9NIcuNT02oigg/8/6Qhf4QqXM
nWm2+LpSjLf7dAVzv6Ffdp7GHC6Ch3F0QXEOkog2l34INpTi4ll9E1WeVlUzJuDTvM2cc2HKAzIk
h70aFugK2/rbP88HS6c2RBGeIPoySiZtRYWGWTPuFNiCIuXogk0kuXjQpDLmo5ACRFduBdHiTksT
9GE1spuEfp9Teetnd0Iw+mbdsbtwEbIBFAQf+rWowONZmqRsdu6EW8FDztY+eD4GwJFJLkueSwZy
nRTTwq89puTn5xZRC5wEx0a+fiVyFqjQyW87bwoxkThA4szzvV6VmtTOfkvvN/biOudPlPy835Ac
VWMWW9PXgS0uALkxywxOy+USLWBnGNd6ybbATEw1/CQHUlDGkHCstfLimso4TGwWtOthKaT6R96b
/+/4EOV4qc7D515NdVjFZoN+qnAjVZWLV/J020B47yzswY8Q4yDjwNxj+7Yj076ET+O4NKO+zeQr
cRfqs+Qk8aUdM9qoJ1Zw2F/0Mh+/A8Cg4w0B7nBkZAHkEs9jf+NLH8UAtHktDdbYxo4HOdtFstgU
vUJ5Dy9fYOqDprW3bDvW/l7cVfZ7qZpix4grIbbDHGgYxM0E6TeTz7Jj2wcv6JxWlZ6WH9BUblAt
SEZ1eeCIen+OHHi2E9EcY+elR4wFZaaeheKATQsxta5WslNUV61H08BdcfVRJaHt9BGmCXEL+kiQ
6Ssy8W78d+djvsyadhBexKHYRCE5qDpOVH8YFI6nGVb2N5xDPyhiTAok7sggLUprur8X3aYHTIUc
9NNBkKf95N91vMVycO2XO8Bd3Jpkk5nII058HctYBqLqrh4id90vt8xm6q8VA1lWggs+9ba0HKQp
69FGKpeNmujKdM+1Lk1HIqZoYGiopBfvWHTalQ9qg+pWt0v+K8kL4Dg10IC6yS5CjDltnhdlNp17
RSm+7pgTPzDU71Z6keUoKrRQSQva5C+MtmGNKJkdnAeJ/q+IM/mrw6Ne09ZykIADN/8655jZm0lq
wg29+XBz0s3NDG1iBDFMEGgchidi8uRYoawbnI4exCa/tAeYKiFizx4TBZV+Z0IzahrVP8ZNsToU
OxT1uORK0PuFsuq0v20a3H5LShMpuaDMgbpVjoS1fCHnujw1CPiYRhfUX3tUArmIC7mtEgCLd5RJ
+5agUXfYDdzlIiFliGG0J47mT2yu1Lwpvg8kwUjeTXGcXwk0ZA3lrfWA4SGt+6nrrrjgGCch9qq/
De1nJiEQzuFYhH93XNRXzdDtrERmuxyqN87xzxjg6PyzBCa+jPJOs2qrfC9NEzMKdIo+eNz+QfeA
4PcOOtv08GHMJvVPYXnpcaQI4s4NAJM4YRVq/luiIoda1B3QjZe99xZlWdbbH1EL6FlnO/U+tlkW
Vv+5gUW9fciLK4jR/0SjVoJhjmDeZzA0mWD0hDJT9JxjNPXitBr0rtROAaIXmW6hopPgTYO03Lh5
Tr2xKhNlZDb5o4ElNU+cRJhhBtHF9fPlI5MlQQ57exZIHRZkNSYIA7ncBRtbwu5hRP/tHrxytbnV
3qbzRV4TOyIk8AOhNLkxzu3KNBt0sKtQewNKfd3JDmmVB8pjLVUkwDRuBLFKWIpXeLCxkK2I9MNY
SQbUS1U2vdGVM5kENONZFcM4UcYwS4ls0VJQhhFPLs/mmFA+xhA89DqJ3wcyvpDS/NzZm5g3Jh3O
AG852dRPcmOODTPiqSkhbUO489SI2W91g8YddZgw5Xnuyv5+1vkO7m3bCICCdTHa+KxB7cW+z8//
Ib8FidE/JKKxZsijPDd2EkRKWFdIALBDsXiTSdL1rFTabXcUjgfYQBRQ4e0WbjovDkJen6Cs5gMc
uMvft6+YDTMd/moNSi3PNbGARwp4rOGvj3i3qFKfX8iXZBFffMM4RoeYZn2/Crmr/c9v5pU/guCg
l0z2lBKsBeWRYsF2wp8vdxWKlAxCXT8FyAWSx5wbmnSPvDxBDlLMEcyEJ3H32P/AOdq8Yr69zcEf
C7UTs4baiWOO2gCqr6j5m2OaniqcX4T/z+cHxR/WYPMpGDJ/y8QKvLZCZqQOmQPr+SS8m7JKL8C2
Edkkq15Imef8hOoALdx81g7LOPcfcmrFu3J1YLwgt51X4Ojl5aPTfOKBe4XFyOmSBffv9/tTPsDA
yc3A6R5q8OsmhG5w2t6GfaphNjc2Fpu9SPeDXxWeyh6B20dHLu5EAYrJKWnyyM+a/qDCb6XZSg4v
TZcrz9A97IbbnJ7+0q7tlzg88WvJtO4dsO85pM5YVRYIxYjSUENWAtTaWMdxzhwb3HX51tnfvIEM
8FNG3+mZ1HyKBVEP0e53x8VI1BoI9siqTrtlGLsgWsCzw/AWySUb22n5JMXP7UrY7Em9Kbuy+gqU
7AkaaRrX3WQKXca3hgY0S39nkdfxMCZJc3ZOJC7iBkwX92PnHVZOKkrCxJOgBw49purB/VpND8iG
9M6eh7j2nIcYPfAkoGhZsjEJTz11xVqnI6Jl1YDc1G7FVXh/rxg4WKWFh33nGRfXfJJwbFiVrMsO
kZ9CCYGCo7bm3yke45TwC7YWMZom7qj1FQBIMYEj6n7vE3qW4fx2yG1YNJaPOQ/NX4RnwPkVfylf
9jJZAWYnc1DTCzjYyt1n1CfwsiD50E5SJlsvt/6GD8/nwLd64Cfo61PDFHMqe8HnZxYnvAk3WQpS
C+FXLqQQQ5PU3GTMxJKSYFcQAVS8I89KRVzyZ0O3L+a9YUtzogKBwQ0hv/0X2i2/e+u4dsJB/y7c
gCU7Xs0LyQPpjppXsSfRGvHi/CZbcGQidix+y1BHOaII32V1Y390YRFv+FCBlvMynkYtW4ZiEHS1
54dLXVlHZp7E0HhVZO2/o/HqxcBPE015Yd8nWLg3rRfto8wlEmT45aakPZIQhMYbgJyD7d5GQIRA
zokuLoAQoKCtHfqZuvDVLXJCdlqhJeXM2dOv64q89/kFZfMslIe7tveC1MYx5K9EK8rSZG8pHQDT
9+RuEQDTO9Nrgdyf+hOBLwoAsga05Z3LBxHa7ZRPImPNyxadtixGC/gi4uY/Cl1Sq/uOJ8WSkrtf
y59dyUz/2fOOYe5r4aaIBORVEQZm25KGhHExvNc2kaWn/LK0+3pB1PuCftx6zSbOmZBQbCuDeYis
oIj6r7bacr4mNV0ZwVEDLkcH073cAOp8smbC90XnXd0Z5h8i8dqVeUP6p4yKcEleE5sARO9XVTVk
8D+P9wM15ar4ZF04YWqOYi8GTjwn6ayd25h698DmCOYY3b/ZvAVLaxWFSbMXNCfRS/3WXHpCQINT
1KF2r5I3DLUmbntbXyW4F+TXLkavHwM3U1DcqrFqvUFyGFKjCwE83SdiNsEJyIsJIu5+/3rWO5Qo
/81zUXanzN+j7dVwoigpTi4K3+29/mqE7dWoeiupYrU4+0RlEN0ZQtHAJ9Gw/qe5R9dCfOWQV5yt
LEcNnGDSwyonl49ml+D0m3EtYfXSM2r76KpWtkWwd9N9QzVEYlHbH18FMTL8F3nN0dX7QlNF0vjY
VAvG2ZlaBXFwnquqn9ubYuo7/TEGOvKRAchW+YfyfrEvjcxypNLkZlnhRrW58qx9JyCaiJTV+mqw
UtxTYZqbiROUQW1gv9fb4uY79/LPeUMSspBZs2O/XK84l62f4jq4G55ujNsSatwiocIwr4M7+H9E
FseqB3GbxRrt/MFNpN4lOh2UWNbjj6EAHk1lCC6wk/v4I6CzD5LuAv67uexRhxYK8W6Msz5iDGuD
LucBRI9hXGj8kRV9rvzJxAWXf+OP2ndoD1dWde/HUcvGK8n/jrWx9WI1h3zNxD4cAQN2yQuTt1Nh
CFiA4J1WbZKPlQICCMSK2ErefYISbDAiGsGtW9Kb6VjlufWt/6UG/uWX5M6GbicQlW99JebpTRkJ
LK+gQEWoVRa90+kVgo5B4w5Ogy1FIuhUqXl8+/QCIf/VwsghR3DbrmyCnibPViXf/V3jX8ZNbqJh
F+W6c6lz7MBJm1kSJY5dd8X54sJuKT29zWCDPB07tgnFF7nHwx+oTu36Pz9D3d95FcH1Ln1WLMWy
vUb41/lGpWPFSe3WhpGE7IGexsMN0K5AWiBrpu+ZnfvHToefJ/O+pnEGOQ1Ex7wwoIeKBSX/66HL
tmiBHWYuI34V1Sfpo4N5j2HM0wJkQn7HpGnUxi+LXrBozy0JvWtSNULR/TO5/wfK3zgA18J6a6KA
W6Jc/5X2nNZ0AMsWYXd3m4gAivufTYbEKyPDOpKGeL/DYZvMHBF1H/fafOXKYDWWKikLyu8YHGlX
jq14T7hvYIMpEGbko52QBo3K5HHcwoREeLWEtgWOaVDTNsRm3xQjPMLjNX01HaeLb0xx0dzdZQsq
Qf9L1hp1NjxKG/MaxLAOpseau97RMQYOKU0WAI+9DtBKGQ4H3cwf5V720YNeJiU6H6S5Q8rbUPyA
v5LEaMn/PXzSiT5S/KTa12JENj1kMzsHQCqX/M3jo45HEs8IAzDriysYUf0fp+4OtmNgsMg9xeLw
P5C+8A4I6tzr/HRYFqcUo0HwA1PTs6TU/Z/hSLobNNxVDhmTppyjJMQoz3AM/aXXvx+9GynBo/bg
j6Szokh+guOepZA1U27yvTXcjzBp6v+xtitffbcFIo/eMY5oTVm2TT8xF3UxnNZOkJQAaipazz1j
F7KZLqoD2B98VhI8bubMzZVyKckLq7nYLz568zj9volKlKicKwg52NdtE8B6JWpsPRdBvzx7NmcZ
hScv8a+mc2JUsaB+MkqCmVnhZcuWDDjFPWCN2PzIORa05pYw9I7lkh1dnR3XVhM0ou0ilYzgJMSd
ul4u1irDMQuR8Dx7lboOJYYRRyfo3gDZLFBhJjosuLIMEnMMTpKdjJnZan/VapzwCavgwP9OCuJQ
mHWY7/DgoNf3r4e+pIH1gFDSd4CX/r8aLjWSNc3cST2ANKGmbUuRjm5PHqfEfGjfv4Exe+XSXd+9
0o6XMwCcxkpM2+8vjj2153FTKbKSx01/1b95NQdgqAmqZnPJq2X5r+EdfkZBC8n2t7ltr7/VMISg
JEoyJn4EDoMKAZRD18NDBxwYnQ0zCzFXKjQ7I+xR7Q0X754iJsVzecAm6cWsm7cS8V0OrWkczRl7
eOHxDKL7HLXMic0HWq8DTn7OnDzKy0svynXvwfkX7Bfb0UQXTG1ZvA+zkFvFRRYaAlSAJEUnxJLx
Hn3dgfo9qM+Zwi9vwzTqd975s6RFaZhSFIaMr0OMlZj0WJ6GS6GyxF6wDwPrG1F9SVMFbnGwGfEq
2Je+hvDfcle2TnZ0V+mXtqDSQ+gbB68OjtbUJKRHPquRsa9CkixHSWkRQanm4wCZliaoST4hWmA5
nk88zNV2vU0unTJrdswGj/XLmhMOLMZ6i0HzPmJmhTCMY8fS3G8CReAdlP9K3Qvv9EqpKswV+BO3
fuDnPWkxBlsIF5mnymxJxuR8RKb8lfTHaiEW/4F7/YLbb1KF8CC0qkzjJ6JFhByo8yXShKqQsk7I
DM3LsWmF5LpZ48FN55TV9IoHCeC3aqe4QpGAYXuehCSiJjo8BbhXQtEfbPeQi6hu2fzxseXfR5Kw
Lr6WSivy3q/ssXNipgZJLEHXrIq2EtyQedLnheMFIAvhxglO33mgS2ump3yhFkehA3Xhwk90CdfC
XO4iBJZ4HNmfVpy4gdWL1MwR4hiQDNWceQsnYOX7W4dF59BjgoARLIPCVcQxMGpvoORDH1LPXtFe
XROw/D0T3Qu6CjmHrFRH4ITfIMfP05RLcdz6Zq/9Z8yer3XvdeG0p3KnXUsMbPV4xN+U3rOopMGP
i+A5pF2CIibJK+W0Cq5dgxN3voR04m40yCZtibjhMxpXEZApk57HeI3P/VWXULqK2Cjl56paWTK2
ksgktP6dQQ/L13cpJ5WhcV8vWsD5mC5aAKSFXnWg0bg9300vU0C+zKNzuN8w9H2sT2iLrKoe2i20
HTWQOVVTi8OkgvL+Lyf3QdgzNWgb+WegvU+je5Da4i3Ilbofk79aFvdNWx1CtCKrjHg65/1S6cwA
QiFyHFbc5L4YmiZ6auPM6UqZeUu36MWkWyfukPacSMUH2y5qusUs5z0PU5JpYBs074vVy4q7OEn6
E1OacfLJxexwX19cJ79cWZ1tqfN1oUBM2OGE5OozUoA/Wg+azYKoEOAadxs4/97DpVEPmbx54S1+
iKSaVUIg9qRinSxZmfk5M3PkGcL8/LfLeDxGAR6mOOBzxscB6fNF2Js1UbbZEwiYfWd/MdXM5Cg/
jykyFtu42Cf4YkHP7eZisR1Yw3Q/KdLSZLt93MqyBEXkTRXo63hE66JD1Y3h1fw29/pJOI2Czr/Y
WQ7/nYsElywZUn3b5KmPUUV8mndhw6+tcq0Q6z5qHOzvxUI20OWAq+iPkUr4U5CkSslNM2HknfI7
7jwVRI2/sk0aPHKwWAaAglUh/dotN5F4e4YAPwsEy2g0c71Fy68O95/tGUGikQYCc7DyytBRgUPJ
7+Bmjg3rp06uEoHwlRXsbDQ3ypdywkRoVxBb4/3F7r1ug4VfaVLLgLSlBaln95o/bWT5X4/z7u1Y
sMdC8XaBqejIpKufi8hy8jQA8pOk7bXt9bvcXtBjsi1WUeK5JZ0EUCz72y+RjpfGCPZtrqBcINgH
Z6svNj4ndSE/moX/ULqqkPS+158jpb1GjKnNkbaLAi+J0jgN2JN1akovak3LEr8Ss8v8IXnTJ/7a
QjAz84GmMhR8JoXRq1s7ITR3PtN/PT4bQPcjBhWdcSAQ2c7wq6/CU9q2A0aN2Gd89XYnJ1xHxslt
aZ7TAbuuhv7tEjrdR+SjelBod1nlUEtYL8YY86A5iBRvRjqluCpl4iICkOmR4r8czDP3auQJXhoI
eZFq7CBSaxTAXf6Syr7VY7UFmcSYWW8qh4fq3mMrKUvCPB8j/TbrqkshxMlDnZ9UYt00QVsJksSv
c/tZ6FVsABaW/M2SJGJETWpqa211J4jpH0pjD6XfNxBUwxznv0lC6d8w1k+A8z2oy9JR3IGSzxoI
mDLy2anzM7RJQBxaSOJyJSy2fwNEBOYwGsbGsdYHcMU5Nwf8wyhRdR7KUM0y0uST7roXIn+pAz0D
405i5IddAycTtCZNfEa9LLDGINcSKQbtRvgbls5ZMnC/rTxvPgyB90kW3eLYce2PEAfFfVV2KCW7
8IDHMg1pu0qMtk9/udP8Uk9dIW8g8IcUzd+2Ro1oM4W6UDj/ARvTO2r+BAZ9iWIG8ynzFJLjNXvg
gIE1nVlc2ISC6aOfR+42G2/lkX7OGQTn5rHebjgA7a20VCHGV6cvf79vFA7IwYws7e8GfmzhAeAi
CD/n86jjWMcnEvqz0jGUYvVg7sS4qdPem38NpEqDsmWrz3iLHUKRdSLklJ/u5g4oNcBwfYREiIw+
BwRrpwne27iBJtq+oWyfTNMnxs5J/iUcQ/r8Cj+N/vJMgsclHXGukCmTer9YS99X003WykaobCpj
jdJl0+XBxae7r/DhiWwCqJD6zZJqo9boqjOqW/YYrEIjLrKbDHeAVMTkr616VFcidnMbdMESM6Xz
woEQm9oOaa0q+ajPz+bo0cR00LdA3lI30pPuWGZRYvTWfkuzZfj5FXaJbXQDVVJ9sdnuqNoeJkdO
WGvSFU8ygnLUMjiM76aFiAQuqS/e65f3qpxkyP14vT/MHQRp7b4g9P62gG/bnf5pSaINZQwNzvNO
KK4e0Lr1W2VyJEh8ccajcDl2bYNjjY3kKmyvEPKZ8pDxCGq2p4WkZi+GJfhXQSb9B4ELG7Jlrs1L
kkOS71kHXl0Rcns3OOX8lklexv9UdfmFc11vySte1rsLUpaead26NC3xcO0aJbDUxzcJmtvfCrZL
2mIEPwN/i9yGw/rug7hrezx3DhA0Wgw2hOgBiwLK15sfUKZd6wFcDYuTHI7TyZo222pNJUGc8sRJ
a87TcddYYPTyk+EaLgpT1+IxNnBMsTpL3mZNLPkjVClRlbFqf504f1MiX5VrbPmsNfrVc6ZDb4+M
auYrxFkuWwfX/lLyeE7Xl2p8C7TttbQZT9H7fHKIO86KLMi1L1ms9mPZ5oD+FtVpE68N/uNQiwsx
YauRsWD9M5RQ90oKI5UjWvaJYq5vrIMiTELmnXymaBWQpta4b7pTgHcAb/chSgVdtRaKPSEaYDD7
3ZGF10s2lSsA7fhiohRbPNBE7P3LxcTQg0eOqDydCmZEku39wsNk3HSt48IPQXXZTdEk8Q2e8NPn
LDvINC1LRcaSzYjNWenXTN++BpiHshoQtjv/6KgbIwGhQslCBlp3AS8AHpLsBXi6Bsod/HqzNWpu
wiVtieQ5+tH5C8XcT4Mz4iWS+Tjx4pI/VI00zbX0bvUOuyzFt65CSyUoHBH46bPSSVmH0wZTUjmr
YCcXkNV5Y9YPvOXLzNfFKkHv+4rXhmih9JX6MfogRk9OitFthYEgN4buEpLlb/LvlTdClE06gfqA
qcKhTPQJW2/s4Iv/fISi07GGILv0iiluBzgZCDgERTBlD9iK4S4j2lC0/AiKpr3G6pR73WRGgJmY
7vYfy4LaJv2W0aFSn6SykuGFZPJ++7P/mhustmIoH11ygGTz17EOUxpVSjBS9jXwe2ot09ArUJsu
X9q7nqFV1uMGRGYN5sN86c115gzSpB7LBgeDHfT2sd0cc5jogu4leRnslp3+CBebac7Yp+afYtC6
ynPgGM7rkOybqaNmtIOy0/UmcO/J1vrvjlbDQrZqV+FtrRgDbIxKO25z8LandUAsiYpbtZMjoXK4
y5scwlnB8FIaZv+IJSwH1zJv57g9/L7r0O9GluZ0xXqPlMl/uhTQmk4WLXvNQTleCH4joKnPVsb/
vEs8oYV1kyNoblnOef0ErAG3I3jISjGeiAqroYn4hVK0Lx4eMOne4m9q0pj6Xb258xyYIQOKgXMJ
ileD3XCEgSCAx1xzb+mEEvQDg4UFqXalvrEaO+yMbfNKuCdn2K0jGcfHZ7czyNsih7VzA1NSWO7x
qwtg2+1DsGQeXJIpTxnR8JdnD6VOM2qYUeW+pfhR6zvlzRZpAEdN2/L1nCffBtZCvi9zj5NKgt5P
ta3uXMuv+e6YZtw9rtl5U0f90Emp33ijBhN84DLWEaYMyC2VJ4VWcEeXI+bK4gD/unXbB9aA48Ot
6+J6wjSaK8xyYEXl/6Ngy5P4UURULaLQxI47Xm2LhZ8IMdzzRqiwb+b/QlXQbN26aPVYg3Yzglo/
Guxi7T1QlIaIJexRojGVOU0eZpo3tFWeVqbtGgfZbv65PE4kE4qgRnVLMacDLiTWNPscbgwqfvJP
Ev3Z5X8LEwpU75NHUTl8tmdQJnZA6HJdHn0PCltoJ23bSELYDZ4DB3dR8GETg4w2UOJwcUjruCl2
/lGlk2vVibyNVUPaX0xERKxZ8uFtSxKV20LaE2SfZmPOA+/i+06p3BhEtdG4BdLzEBJ+Os2euh1/
2/ssCf8BnCG4NVANXENEjoSNaJ47oDH/T8QCmgyvRSzQt8u7VlvFFQtfFCmD+mrhLREpFn1G9urM
d3BzCiuOLSC84E/9HCK4FpD+REi9Rilk7QrTRQ3isJDdQqOabkNPleu3AucEyXfkG+R4YCnvc731
3tU2kTKiAGuUben9A0VcOunpgwiouNFoSgd04wrQCqKAhAekXywYb8FY1yCiM2O0VSET7lmFFyFL
EsnAlE1WSDuYn7eHCvJdiuKuKMwMl9Q05Rf31Xyis2XNG62xVo2uJupxGsGln64IW40NNU56z4+B
YuBX7ve9Itp6ds/AY6cylK6ZZJPAAiPADBTV8hYXrOJy27DngnWGcPN+qQwW2ZNBH3h+QbtvJcTI
Xys9Bdz8LDAJDvaa12+hXqI1mlwLM8vZZYzFLxlkLidXceIeYtqy0Xj7d5aQiXO45cY8eCcJakkZ
0AAQ5lFloO74Jt2qbfPERk8or1h+urGwou9h6+rDfMJNMOO6291Nj917CxG3N9pqqE9hz9O8kZyr
Q0RAiM4+aLgJ4qYPnQ4ZXtdZKfiOYFUjAnT4eAiISzRCwgyfmJ26jBoOtYIAi5Ji3ZGfhmFo2RKi
BosQdS/3viVREVVeD/riaFbNfFTQd1Fkeeix47oFznHruKZdnwaGVoQolsNPJw0eSOXUCwBmaK4w
Sle+CO9qktUNiLByheW1bYGP6pr1Yoo90W9cBPEqRY19x1RgwT0UNnL9NatYpfyRCIuYu0l4VaL9
Ju12Ud2hmjNf+GYgIYKv2VUOkvtpjF2akucPyE+4wXr6n0gto+xhd172K0dEDW/6yeiWQPPetnfV
DzfBHw+BOyLfZt1FQgzgNMygYxV5TAv0b/J1i/Yzcm3r/XNwelvRXkJlTXOkAWDVoM3s+QzcMtg2
Vbczze/qvOm2HfKuKihScr0+qLTaww/TnSbcxgv+dux8DePmMd9OYQT43U3hoSCweTe+uZQR+Ela
XfWXQmEs+RfCy6Jlt/E17MIadCTYqduRkb3MnY+NKGafzs4Al4eRhsDUWM6FDS4c5xAblRxODFTD
97xyo+FTDu0FyDkjOg/fKKsAGvwkMdHZbi5Tpty7RRCMqKKS+wO0I11hWbPUEdqelCXIxap4kV9g
QA8EI3H3sSnX5LH2ApAOwdHyQclGsOYdiwgHUOmU4twtPp/Tivnje896+5mkwbS01IXNNTSj8L2H
BHI2ceK88fQNs70aFoBn76bwswZHgNJ4GZJMr3ohWpXMR2e0HB/E8uM/snkStAB0F7BYfE/XXSLE
0ix7IRk1+5J+fB0NHxzprryeYbowyrNgaBT1nphTMqFqqjOAQcQIaiiU5FeDnQSEIPvcLyn9CHpf
nFGjFuBuhixLicPjVzcVesgZVTjuUdzdpDrsf/YCiVYDVzUcBoEuKUPmgDt+lqv/KSnSeapolx2p
/odIZf0TOXSiYsnQrSVIFslBLpyRTYmUP0MhgvXdqA32fPUPDL3UN8Nx6u8kL0ufQfvRWHznvv/k
r2wq9rFEv2wEGfGP/IlU5PeoZidSQy74YwewfPOhIO2fW29rszRQCk5uY8INVNcmkv0kM9Oag00h
7NJCuOObEZPJjGXIwVlOFXjLrcaYXllCFrRmO3KGzdz/6PdGSacVury0ewEHrm0iQf6yCbsBh0X8
LeDexBkRjU92fxKPDDCf2RU6/ZxKwMyvRuW1NI6fWkur6SERF9SMEt5bcTaogyfAmPnCaypk4Ps9
WZENP8Uea4/zCsbM82yNKrHsn9a83GHZeb8sxauaX3n/p0l+NmHTiCljyEOpbBCIN+AlzsX5PCPv
W/aJI5RYH+qb+Fv4yOUArc49FPGHgw8iXRXWweXbKVg3zNf7IioZczmwYmT5c7q12U5V0R278wrU
sA28WG1OQ90KDOSjH/ikyC+8HrHz6N+sKrOx3GlzRhl1A6twpr5whkJP4KJTuLvJa2ln45WpiSs9
hzOOj6d0IZxLFUOYMM3vUeVnCqACIeRzyhmMnhZs1Yim0msw2peiIQAyDeInUnXQ5LRzJWHV556O
8P5go71LGPihEuPpvp6vuIkpWNEwm/OV8+BfiksPtAm6R/Ccmju/rat9QBeJG1utkXeC51sj6dXl
XpFQbMqzrD0WeEUXFa5cNMeWyt4qt9YHqvOhgkPqjzzpwZNDYsYeme3OfliaU+kSKULvMO/fYY8U
xQiGS8uuVYMJwJgGRHDpWPBFD5dDQMkzTNCEaUqFNyN2CdHeRTZv97AzUKlhEQcqRbAoRjhZmiz+
WzZ7BOy6aZ7pIkOS2qAm0vJcsnxMnf8R7+gNKrDZZmUcVU+nqx1xfDvcbKBEaMANL2//Ng3GebBp
8KUmtWl4q6rAIGIVc5oSpQFlgByyv+txt3LMSEpu8M9EjcYinmPcllFt7xHI+gf4HDJfSXzpBqAe
BLVtJ9i3JCgceXOuXb2nPiKcGuUsYMk3VblAl1LNO6qt2xlk3jUU5TiA1XfF060jtFbL9XxnI86v
qfIay4Re1GZUrwXO8gIVL5IzPg5pHsOMl+Us+1axLwNZZPxLQWiKtFAdbHkPcVj/zfRoFpk1edhP
bWBNn7BgY4iNvppEVrO+vGg2G3gBT8d4tmC+qt4LagSa1UIXnAV9an+aJ2Hy5ltkUmjzptzk772I
AQipgtYWr4JAJQdFtCsK2LYYCBAOWn8ufCTqd7awe0n1M/lVXXaDIpZi7jImdrIZJgGG7i774I2P
D7xfSUwVl8LDOvF7ofsptUdQn/E1gAY3kptVI1N3Wk687LIH9hpHVQXAbbgnC2PgxSWX51mvlg7H
J5JbIMEcjmlG2V/lj12pTrMZxPZ/UvKzD4pF2V5j7TjAhu7zrPmFm7sPRyffhjZ8t7GmWGyOMyY6
x0g8hEpdEOlElw+KSWQmfqxAAGZUS4EPWrU7l1nROEDnA4cYBXd/b1ZnAgaQXOR4B+cCiwJgSRrU
cEN2ng+Qb1NnuktWCmDIGLrs+jZ329oxeZqezxFrvQvX7xIihGjn48mKnnWjpMn0NhOHoejBBY8e
yga9ZQLIIGDyt7jQXtXAI6i02plmQjbjlrkeD16PI760EJTv7mrfT6iV0F960cAoKN65UCsnR4Db
d/eZIoJn2geXtTD9+3e7vCp7BXKMW2xdbGQP933878W/DeuNUYDZbb3raGfxMMk0TRmrLQVC/lQa
c52bvXM95j6tP5Yz8Z835lvHRZILPmmrQHb0fftOD+W+DL6gMqlfLDXM42UaVylJerJGGwtVliTw
GiCmMTxAyisamdG0m9I3vt84AXDJTtP0N/6iwTA6X4xk7AojI2JRKzNVmGPK5PYNAEm3qXi/s2BH
Hu15uUaOdIkdfj7nAgw4RH7chgiYWl5eYvjddPP1Xv9GMLDGTRn+8kzd4mG0LHo4hZyt89KDcoc9
fdCW6OwnybPp0yNtiipd2as5/GVFWS2SUka6Bu5gzxntzDb6h3GCjkeszGApz+H3ePk7FHLu/iP8
/X9KPO+ghWzaE0AlCB2/UbH9E7tVBR2l2mge1gFnGLXW1Dh9edcgIpdzDUIHR6EuCewg+6nIPmkw
Umv2qhDwsof2BX5K9L6oQF+GHrpAIidtZEby/a6yjMQbI4rit9D9gPXS+YLySa8MPUTfdnc2KTeH
p1gKPe+R86qoOQmWQCFt7vnwaQPPAo/W1BrUFsRlEzvdc6WErBORs3dmrTT8hxp+FSx2lrRif9ZL
3rc/3M6HE6YyrZvKW2wsKxGY8WSCZ7iWxnoZCM1MciP+LvHx8/xafizuHCut1dPIE2OZoNZ/s3Bx
JcGPnrCZbzEtdR0FB+v2dRDbc6ng8o0qcfm58T72+Mq0VfvYUFJIiqpHCepeSCRagT/3DTmQBSxd
c6NRszXG+0D5aLqvn/y7g/ZNIXbQl6PvWn+OGHZdqpIBUB7saQMnye0djZZfA34irCBedpRCg113
Hn8j5LkuYKIy7LEOyq5DDJJbmIIr5gKEYqee9DZovA3FQEH43EFKO8dT907jTsvkjT+1fYR6oAhh
OR31uLbtgSOP15yJAEpEH8NXwvbTdeNTLxHll4Ns3J88qH8RTKyheSXRRMm4YgLDyaVzlvvYIwfu
5HQBlYRLUeM2t2rKR4+Q4QINnuIAsWPvw2PEq6lkrjb8Q7kjwP/1v7tfi/cJ9/AqGghCXMv8h2Sl
m5+g5MchAK+zN+NS7CXptrHTYBQK9TazOt2zrdwP6k8j2UT0Fe6BdYXCgdgYDypPL8qjhV7Q43w8
v9tc8/TYSMq4A3J6rLQThDPgOWH3o0pTTQbtSbVT1qL8E/UAuZWC7xdlQ5X0CfmoAB9Y0teGoe1g
GF6abdB6u+GedWWAjHalG+jgcEUQJJnUUY/kldehFfC3XlnwpkaVyMLK028LBgfzduigoTDfwycj
t+KO56NvZWAyIpVfQHWKcli1dxQj/xoNZ9s1dai9F4vuDXOVJ8P5I3WdHEMxaaES9YYo6zllCxCS
txetz74T4gcki+tgkpYh8tJa22kg4MhxbgQb1grM/wQNqP3ifSYSpGV4yv1Q0b1YhEXCkdDD24u/
exSnl5OnTxnAauN7QmcYPW0lWxFSykidp+cfIgbS4e6jiQCRBdou8bd61BRf1qFQynV2vRF1xesD
S7HqzzPefWmiwDmvA/rnaFOCefO2wG43pv2AY6DHUgCdLOcGoqRK/lL9Old8USOZ9BxZ56X6apRm
cZ2zoXY8aGw9gr3nxE+K10UjCoZLspfFJ/xjCVzexl32Kp2kutbvlNhtAzqNS2V4YGV5Avl7Vc03
Yudw8O63NAY3XxLP/JRd/FvBweTopWbXe+7XVDp9rMZ5jP5bGSzJzSDk+uXFuk7UENLhwepiiC8d
fXUjoZhvXfbqOktyf4/lGVEwjtQVUp0wvm4W/zVi7z2gpNGhJj0JjgNytUXzNaXH6b19jll4usg2
ytf4eG9Vb9MCd8ItWC/lG4+6mwEplmTntWi25a/3OOqXF6NBcdCyPTxwQ5N+ynNPq1fAXSKjsHw9
vEs/hKLSr12iZnQPzecVnfHzsZaZCx/yyMWUzU+c3Zk0E1kbA4fXEiMbKtRkhdIo9MDkaygsjS5P
Hz3nZswoIlghsIosBZjMIEWOGDzJ8Iw3bAugxOrgQcPYd0NQOFVj2S3sVv+16K8dAvRiaIlnTRwG
jR+gsinV9km1yDV70ngcQDex6wVI395Xp1uVsJhMd0VycMuWN3jGQgsQpJoCo6MgdCYiZGM2poZ3
C2n6qwMYA8ZdWs6/xoTu48t0NjymBcyZiQJ0Vuw/R42wvJQUtQhriZIVvjJuNoDIQ7vxtH60gztS
qgEMCqux3a9uvQ8o0+vigA7cPVg5wstQ8s7rqq8YZcYBkbEh5j2z+vQwJVjgKtHdRZk8W1LUSbil
YuB3/iCLJFF740zzokny92yrMZsoqrXY2feRwjCCIpvo5r3I1Fj6mLwtqWSmYDw77J68URlHSWzh
Sw6v5L9UxiSsfz+Eu/zOYP/n8aOSE93S0TVsLS3l731QCXGd/BCc7AwOrSL9Mji5mO5Z6ILyfjBt
qO6XyiICvLjfxk9ITCSX3E1KU5VoYw20cGn02c0ItF7A1+gG5zU7cKmUwwWV+ZiGfJ7/h33R/S71
YPWqQSUEOgpV7lVh4PK9yVLlrEOq88XbSftb+ShTvLU2QaPdEfFTl/Krt/iThpfYfYR368R+ZryW
Jt1MqlNRqyrjtO5RzhIZbrR22V41s7r1xzx908rojIIKTRZJ6fsjw2J39uPuFCOE4l+GI+wQprrB
U7R9TYzoon7eTvsMCz7eHRBeyE1mVW/E/12gID4/dpKIfmPeMNayxTJL9mbtbRKYsVlEhAL5yotX
5ddmKtE7s7RT8I+bxHDkt4FX40Qh1KQe844A3Is69nFvYlE3DLCzF4/u4XmEaUWKLp2GVtm+vS6r
Asy8wkDyyU7Ey8izo8o1YvmR1+qA525NTXayjJ1M+GUyxuhRpP7jxz1GP97xwNWi+g1SM3qJiOAj
XVyXx9iof6kvR58PA019WQGMCu0wAnk5Db1vTMHIaZAugoIQjLU3TF9uVIcdVPloF9qq5WpSptKB
jbF4cowgXyS3izKdAET7hkywc1bPagINWg8/pNJea3WsgeZnK4Nz1E16j+iEVyZerb5Vwg/WSrlU
Q6mQaO1146Sc6UmQCgbEALr76Kk9L3vYHNfuhH3ew1q2ieYXVkN6wy7BPwiI68ZibIeujwgCPHyR
ii/i7Wj3hFG3+ch254yWTGtz1xLlri5NpUnhb5J7GY8sa5Q2r/Gy8ngPJOqyOLbQjAoIgVp5UPIw
nxIq/O8DkSr11dV8BxBGk32WRjbC8m8vRGD6+/GboPqH1LMGLMaeWbccQsnpcYI0WmZXfVZ/Dpzu
YVSpj2u6wQM5KnEF7Ecz6tVewXncGf/3yzrYX2uJ02RoivYjoB7P8LzVNW11LQO3buMNQd98wpov
ykmRAGyLOJpkxSF+3JPv8hSrOEvQ/bs2X0ji0Eun+DzKX01Gd8fzVOfZ0/VdyjYWVQLU+ehfOlcR
fcX4zKx3kR7T0TyryH8vz6HvSaDJ7+TaeQUVk/QRJlrP1CZiKjfQ41SRyp7D9QH7hFnR3vLP6JIq
YrMV3zoNk+wchhYwp7G9sl62LdxFCNn8iaaOfZDfNdik1Uo/Q+Y9U2N3OnW87IfERzqDXWZPjqVq
era4gHywDJsAHoSZSsvT5y1G6MLM8aBQT0z87e1JCNQhPy4kW6UfpwscjQ+ewLdSQvtBQUh+GDad
zmK7YJBPLCXC0XC24IHRLvyf+yUB/V7rrc/TnCsRptrTfQD7oNmNEBP6Y5cpK8HJThxRcSIFCP2L
NjNrxUEuxwbUFIiB5dy8M1h+D9trRBZvMNqdoAWC1Mx3rbnGjQTFpkLiczQ6BiRjeLKvBuu2go++
Kwoz5N6KUZIV7J2SJoHj6O9UKFkKMRKK55LadM2e5N6yRmen7fqDb/AtvTilIg1gyUH0AMbl0wKD
cuj3jHFPKfXAOjgjMdHZOMXNzLdDgXk3VDRGQ8qacNJ5UeivtjMxObAumDQ/GWXjKHuoXvVFy9Nu
fO8Syns1Tjgd0q1TfShq5aehwPySJ7Qn1Jepb9XJawCmEdN+NO0FSs5zptta9ZGXWteGv3cAM3OG
Hg9dmZ+nzH/lX+wuj/Jd0l2CXkrXTeHoTlS2J2p/SYCpDFTFemA4QP1zJ3JVngbW1IxR1tEjpCyc
MA7gSVyyQhd/mGpuSHGtHsiYMm/hedRO0VQsgI5aIv5D37zpA9qZJRvJfRbVmidJI4fVPZw6qD7h
UPrtwZyXiqyOqTZEWh49DP92ks8o0/HR+VpOMRz9DsS8rpwJmPwqk4teImqBMwZbK2qIVLQUkTzs
Ltw3j7spsk20tGB40h7fBbSfYlXo1+OyiUlDhNC9qb1G/UfJcBHiu39gKh3j1bOAdDj5wQXYDYoA
NPvwCEakni8fEsFu2m25WdvVM8ifitXPYdczYXhIDxO5XJfaw/ThYI79qC1EZ56TpMGhjjaB2goY
jwqM5a7Smysca27Dsp5QmrkNgXTvKqcrIHgFVqNit5+tf+wCyBwhLbo27lP29WXhLLrsjFENU7FI
UyKFC46aN3y6SMpERdRVn8XqwcLMuHD/PU3tkMuZbjk2k8OMN5K9MwUwduM2nf4YC0yEIbTRYfJN
wNJHmpJbhlnp5uewPsPA305SyJkH9ZF/SnO0BBqPaMYAcJjyODn5Qy90RB/9IWTy6dlqx5jCKHRW
yIBGRr5jm4LimKz2Y0sk3kROxvv7M5uQE1jlkYcmvG9eNOXeCvW5ipMOVt9rPHivgCt8gxZX2QwN
K90eqMfjbPW3QvQv1xrX9O1pxbQkC+NgTHoxgWlvXnn6IE8zVqRannBNS94qsGAADiCkHQAQ1qAi
JbAka+z2YkxhTUdEen6sp3icslIDNSZRqAhmkJy440nvDc+jzE+Znk4vZ1rxkVXD/ZFtTa0uWPHj
BT/fq66En3DcvKd9ShuGM1b+HM/83y1IDcTV+wrjkXC6ckxsiK0NFGE+cFZH/BSkrvUkCDlcmXJn
ytJJaPE4tvSps7VhFh8jNbyB4yaK2dUVoRrysVHoEatZYvlhc5zh4Y+8WZaHmSkXKNnmQglkvqcV
kk6xQqeCsynDeawtipjjvED6CRF06cOZMcQN7Yzw+AbRmh8EKaIe58EWG5Y/0xksAUIESrEk7bcf
CRt64wdt/H1ZdSPEtOzTx+xMiNprDY/GGsRBsd7vQXn7aEjQQE6RapuaTky60nqHWnrbM4LrJexm
7E9yVwGMX0v2Ddf3Y4Ls1pS7juzfJyVLASwT1Oy6uJVJr8Sh3VPiRtFm1r7RkfDFllWrIIzEKYwd
mHVoR0S+YqTIt056amVmbYWwbN9AAkQAFSIGoQe6chaDmoj+ztewZlmEz3gbNwBVW4OZvQBlyLoZ
tJ6zbhBeZL4oHFdvpllD2AX1Z67LNyo/oytdYD0go4msXm1wUDMIvuZ98nOPNHAVIe9BOOdI8VCZ
EImcewrnfZnXxDh0JW/hr3j7Sy6vaL4roCOKuTzimg9gTRT0FxausM8nMV95TElvnqVdzoUOU0nt
tAtuB2BmYSTnXeUtktCofi7FHJoCrcAwtRuyfWGG8WFQLZs3oDCbczPXupFEYQfWBVZleezcWrMf
XC1BdCpDB2hx6rnwr4TiRqEf+m2aH8wYvq5VeYiP2w4bobJuu80Nw5H+0ISd96Gs9pkZIL7SCamw
cxfhjO0qnsY/rf3Moyf/ozVX/4cGStlnD9JFXiFnnu/rdYqThm3fN0WWJtdLjKmIRNRlsK0xxrPn
9+xjhE2gRnv8DLbogwmV1GOQHIBcJ+e8DwQhaRxb9kqRVTDe8lhXGBgapEQlec+u0ALz+Gp6aRq1
ylbTD9Intu2Y/+DxRFGngrgrRWrB2aP9bijI9DuQdOTDR/FSugW9pe+J373SedlpjpQGeIW1TFgC
IncDDXdhLcgj8djZ7ULXv+Rog2jGHh5B0jyk32sWVJLIQ7ZYI4seTSk1p5u/ti+DWNI29ozsnqvF
Rm9WOclDmYweM16LIvGAWzNKfkyUk6tScPnzO5dmhQmMpimrfs8pZQki+3Vf/vHFjuIVExfYnk+J
w7ItTbZrTVU6PwCUX/ntdOMctCgKrRJUFyDSK2OOc2apQkaiwViD0EgzXEtboMw+9Wr4OoIe/L27
jahEF9AERjgdPxB/hlm84rcuClfutjVkiMXvMSFlc8hxwhXF4/gH8BziZhwB+u7pP4e/+Me+4i/j
4dACfRoeKwqReBJ+L8FEXk1yMGNAKokfd2eo3PmQVk38hHuja8QajuzYYOTwzq76MDG1jB9j206W
9mXjx90lyk+0W3ecENwVGkZOQ8+TtClWsmng6h84ayKpFAVAPHz2fwVMFMCupw3FunJ+1lwGCAka
rUhCCLOlNyQELxLn+/Nf0EYN24/WyUw8P5v3iXKElqEpuy4QEvDuWLCph513M0LXAt1J6t4TgOvS
ScrTLizY5npocXwjN8GiKlyTARveqVk9dih4DlpZjkVugZsY4lconkZJt0YdxpTC3BVpHZx7lzuz
dIjsjdrEuj0F02qdlhNHMbbk5UiswWEUEycG4HIl8GIjoXFvQY84h0baMhqyrvbMno0fSJSHJaPd
tw9bWo2godo4cxOS6MaOozUVjaosJ/EAShQe2VsCDXefsfWMz/uOGjz0XhmLybLSzg5zd9VShxm1
2xKuVPl8AzuU4GFLthc/elz1PM0g3oO8TckmK02woRPZSMS4P9Axs7UO1Vg9dTiWKohyUPq1zEyn
kuL1SGG/DeuboYbKCZMDjSsYaRSQ5uO6k9eMwM3Fka8VqMoWqWBEFzWus50lQmE3Xc6FsOEIAgdQ
H3fVcCJ0DdcFEsv/y/3VGg5DctDpv2/GEb8B5qqx8OFbK1KSh18Ugmx7KK3Z2/UHjNa1ylG8ygvh
SOaBCYdrdvFcv9JFw4yugMzdJfx0iK4Dujl2sUVk97K8pCZDHH/MQQZkFattbshhhGQ4Er36O7AO
JL7gAmqf2uFRChwirJVgGN6jjt/P4zzoDVgMzUbMcVVl0rjXw7zvAYsSudLqdeY6uSt7qCat6zbg
ryuLDmFGMuFn2NxhgNlF+K3XEGrTKL4Fl9hsHczJHG0boIrSqZIyk9dhur7zHRwgcg8jVxs0gp5R
bXX+2q0/il99EGv29X4mUT5s6SuJoDk7QXQ8QOtWvJDWZ5JsVBlqFhhWdewu2W7WZIQG90fzdBs5
/+O4hMy83Zk0eXgGScfEb4reg/XcghRQuWvKMvgDcYfDCu7Mn+iB/u8Vb4fNkbLwrPV8KIMoKDiC
hREZx3jwj13+nS/HzLxDM94XcqA5ZMGNmdLIj8tRepxsu3lrtrrsztpKapyEfFnyoLPp8CFFx4nf
B4xgEYPElY5mP3ZSPle7sgkNu8taiUb2weF9JmmYjQO1aUskC0pKCIxCsQFnlVFYf2mQmibj7cDT
rzpl5YRoSlthlorv3DEV6Y4/CQGFBZ9Jr0ei4d3vMwSwx3A6a4WIv5e7L+visf2GyQhVGqyCbMI7
nqxSZMo0Ym2eq16tMX/r4aBbATZAlMGAy5YfaqF5sxAywAyhsiqbDh2SXvFPXvXu8mLlq84McB0v
zjUqWwXCfnNrtmkO8vVkKtCNc80ScOTQRTP0bdgHlP+Z3h2jQdatN7D6tMmPk89TOFK0ImAbKJSd
DXHWQOOZRntbF2wwepKqr2NAkts8hkqingy8+633TXqshNf4CdSTGHkepLTvAZ86kJyPxCiePljh
FNaRmp5NIYSZHlZ1jc8umaAPOYiHm0BjTgVnzWazZskra1ozIPEPTIlzdHL8tqtHblYnnmzjOelM
MsLrmrZtMmS20YKSL69v0kGifsHIGXbFAjrZN1o11K+RwyCoE8XcRa8apxABiDVp44B9lfd83jQE
9LChyqDAVpdTa4UJ64NF0kuOflAqBARWSMkGxdvItMBTiIGbyVU+TbliFK8JnWX4IRu6epsJuwMP
8lh6XF6B/sgFk6JqjFcVNb+bufpY+Mw2XsjPoa5ftAS4b8oABc0ck5zZcsrmcoaBw6tYlWfAFqJe
n5sszyEVVdFx6GJYp4IQ1XkMWAcaIib6CXk8lKPwGq6ElkINKUfFeYR2c/LQ9m8gqAGJV08S4I59
01jpYvljtH2zwQw6+Q0ZpNcFtdDsKdAXnRZfB8LjMy7rCrZGiiDMYM1UfZNbBseRRzifxHYDBQZx
XnwQf6GWJYbXSt0ng/DS/DiLIXgJJ273gxEyidKKGGuM9KrXltrBIuQGpHCfOQ2aSjx+TDAgwcwo
TErgTr6xseUANVW7onFat9QY8cy7ifzHlHlyH17hDDhQ7v6o5b+A8NJNBzEAOeidMAw2fLXHvw8b
Kk7KkSsa54OOIWdRda78DVb7KrzENl4btTTfGaRI3TTZNXEpE0lQHwYZ/bDHjyJA7AqUKg20l26G
7Lu7zz7AJ7D6H9T2vOrb2YV86eYQUtWW/x02w1HXdWe5wjcDqaqdGtJ5uNvDTSodteozHi/iI/Uz
n/wv7YeyOjatT839gbnFcdAtavc/DxWg5sEljTyt78vNK54xf3LJ7Qp+XYzj/FDP9OmeBb+EI2sj
0Gc76D7LznajQ+qiiihnRBOlo+4m+VBaSNmwfVYnA/ClAcNBhxt7gl2rfoQXP5bVd3+9oXLeZTng
u980edlUsMSQ1n2oDNw9XVPKvnhuGw37Hm08q8EoDMvoDljqjP0Y0qfIdSjiZmNw/pLj98/LG0v+
uSjlHM9WD6cdTNNMUfl4A5ySH2PIyxD55iJj2OLXlihyCrTpPsRq0lDgMk9nbFzmHOiSAzL6PCLN
VP/qHsszEAd1iJ/kDhd/fff3fDrBJ2TyGvVRwSjqn3xfzgkmGHp3lN1Ymteg63ZXGmHvkf0td+uX
/WQs6KIvmmPDhc/GmYeZzHKLBF5WGMlVp8uqE7WaAdKgPamtcKJ8RLpkOmECIGxf+iyY8xFAxr33
uS7oZ8XLCRRJ4uFQ09PIGyrbvQcKdh+KCt0gNdgiHxU0HHpnbTj+JMUqRA3VA8/lAgeb022GwKhU
cy95/ib5BCCQrM61VmUhVblmNfYCIHGbbT7kyHAqZ5DMD8hd42IlEpObECCB1Y3BVohqIhUoeanS
bsJtOeSLiwU+UAhKbUlQZwwsfljdVna1VRGaVmw9D+IdMxVtJIEpk5r+9Yl3NCJ9LjRzBGl5Sobt
ioClygVjnVy5LuICkEv05ctLr5tLJf95ah7ogsJJkakXU8B0Kb4h7n6WKG/bkuPONuaLUKyOY/L4
eQPWEpHntH2Q5JrSFlr/1WXEAdHpzXT2KzZXsx9iqt71upHzzdlH8rZcfQlin7C86WXApQc1ArbF
sf+6br0vTuAYSf1X0VSKA5izpNeWPCyf/MUi+ssz9V4lomFsZ87UsBjhxGCdNf/k1OD5TmeH1mIR
B8iICAev7Jj/p9K24CY22u4Pc1tT40iUESYQwqDagQ/kq0SNHNdXzS0/gejE6CAbUX951GD+Cu8t
Kejkiycz0pBmIRoQCy9B7l3xew4RTwYOH847XH892geUqUL4n8df7XOxGBbsYFhhDiqykP828Zzr
kQEJ9bXYm2JMbR0JMrJyTa803obunjtHbQoCgZ4vF5LklnOMOrmPWsvDREGQkuwfdcSvm/dzW6js
vuO+glkxw7ReuckC1njSG7q1pU1Xn8HqtFQo834Y0tS6NpS7by4IvJfa0CzNbi+GpdA9FAvNs5Co
pEyyd1Ro+qvYAtAcH3WD0/FIpiYWagPTWNTUfbiieCRx2rqVvE/LXiLyyQhT4j9FV/UtsCPZYb4a
n2/F0dq2Yg6Wbb/2bjKu2V7j+DzK6qcEtEXrK+fPQgZRPGh5ljbVX7sizLfVD37DTFnHOh/b+gBK
gE+V04INpoIhCTNgSU/2SVvS416eUk++AynaxnCjrsMENOCn1EWJhymUHso5CDTnljFnPT16l2HU
NphsJh8MWfwyeyHzs/AFCCggLarFunxHe38Kl7y08BeK8oN1k3p+sLc2wIRP/yPJ3jqoDb2Xukle
fwP/hApHgeBZ0vteLNTexIuDUgvjEJKevI7gXoDtblTAXNIU5UkvZ4IGOC2yIPdnZFGJEH7OmByL
vbWb0T1/suKLhcu8wOfZ26CSx9xryJ1SB/f8BtvPsWxEN6bWi8tBWuDOfEfLYdK7EDHMMu7GqKW6
0+fyjJdWKM7onolPoxMyz4UYXr5uj1otiVLqxexjTCwgEJQye+GZP+mYfAfe7tVCiv0HhXZUFYOh
8DXlFVCyj/JhiTryR6z8nSeR5m4qh7bjfrENRlfE4POxJP9YBpzqjxa7YOSxIN/mym999AW0bAmh
2JW4HL1lbUAVc5xXWfqqEXdamdE61UZPpNPgOgafFMdvo+fcsCS3ARsxzQW4NWds2HL+8FyC/+YZ
jnBwMOUMIchFFaFCKtOCxmK5uErXceKbTjCCTjDV6PKoQfMHrfXqJYGQbNPqrCyjHWUqJ3Bcr6h8
7g1htnFvKku4tCTfD82YJp3wLRzS/jfZVoDFGh/IAKbU1TInPejaL38574xyR706pdSjlGj9p2k5
cE9j59Gj2mV7bCbWd1FRS8dU3F2ibp6rGyo51PW7Q3wQ2izFD4HV6bChMXXf62ZgVANSlITYvYai
sgNVfWkBalFj0YXjFfxxnCg+rvmGcHBu7L3nEhoaDMqnw7pHsB76O2wD3rNCNvTt/zZ7QVoSn+7Q
RNgDHsE/pHNGISzxtT0iMuobDUWsc46GevhlrVae0sNnXJi99RB5t5DKTd+Kk/jXVHHMEoUJTY5X
4IY2E2inbnZ6/JEQRJdMBiAD0kp3sfSKy4anhfYwjSlmC7V+qan/B+TOKZ/b3T7rwYTnDJ6N+xRd
qxGf8WDa/MMaVNbZ1UnxnbnInI49Nt9FpKQIWdVWDZe3+rBfk2M5BnHl3jYKV4n7vAaSmIpoftO0
MRnbQDKEfuidDIzKGfdA1agUVHunTVWTeLPEVrl1F0zTx6s2qkeZv6RdmlaJzZb3jCrkglRBvBDG
8VzRyV82GcDqSquT3YaLaK/hv636lKzR+d97eQJ5ANthV2mC/bnqLfmTVAkn4vsurVxP6jMo+WeD
Spu9WLyNJv2JbmIZsGULlMzTjItCa0968Z2PmRVra4XvsD2WiHuVdztXPNn5lkwKi9IoGk9Zbkzn
w4EobKxot1vVBHxNWJJT1nton8x/btcLWGiEHoi8JF9W9OOqnGgsUwnoz0Q1wSWnrc3CpCRXtIS5
FYfPpxMIhRQiZTSFNhP1x/3ZH8NU0nnBRjZ0d2atrg+C7GKW9o5tbj004vB7L1wj5561QeTLl4YX
EwnFyZrdr8YYM8RMWCg1tisJh4QXQMQLPLu8Hiqm8hrgtm34MzrziDda8b9Qk+c6bNs27Ui/4l8b
9jrYse4eovHvoUsPTo51p4I5F66D3+06Ek9kcWTUAjhq9y1aYw3FOCIZIet6QK1HO7pnDjN9YZyS
wcAHOS0Zrdw+YDYvhnw0Yt05c4X5fbvowjN4UrhDRdGQqXgpdyUpXi8nqMbVIUwcXnahvMzazfCH
jBdxfbp0TCjJKbA2uORy6j7aH5c956a97VtfDXyTfqVm8OGWSJCjIEBk2MH3BNYKs+J6QrTAoya+
gRVMa6EP5puCk9WOoSL3Ilr0WvOJ9juYDqoLkUuYQovuTLL3q8MMhPv+m3c6zodfbxp1MCkcALEU
l8hlS9P/L5nPEIlFf20rb8chFyumx3r46dntjDh3rVAYcJ+ZGSMw7qfdVUPKMs7YuikgQ31TQJpP
CxnYMoiOv0jT/IfGquNcvR5Dp2T5AiWHP94ctCzG6Dclvyd2dpqX4RFEhSH1Wk7dgbjWiY5fQyiK
KJbLHXoADvw=
`protect end_protected

