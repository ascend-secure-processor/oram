

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b+s9TIKQ2srU66ga6NqYLlMsutHIlYRsOft2wKFSwgy+hRJWLRvGZpcDPDE9HCUcI3iRhzzHED7m
IGmkFXOWBA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jh0mDLMUl62CltYrgOjVvK/Dm60IX4TBPyDuNbBqv+aCEb6AGGfkf3B8KT/avKj4QPCAyg5bEu6a
ybQnHxeozporhivIIXNWT/tSp8Qkl4zUcxyBz3m986uvhHvrh6YxdmQV3GIgIU3JH69+lqz/UXh+
vGDjcYJ/uY7meuec+PI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vqxEYsq6p9EAmQc2kuZjDeW3B9tQUGIsu2NkoxbRF7EyXuIW4zNp82Sollimgs0aaJ1UDYFhE1lb
G7jRxzcWwy2lVXLgyWRU+SZEk07A1A8UWxzy8LRHo2nV4zjjZiN2T9YonDQHwvz4+JGThtvn/1Z2
J1m0x6dGKYjwaGz6Umt5W0+7F0FhnUVLXRr62UOkysYvx8kHcvMb01Z79h8Lx6r4sMZQsXE+4mjR
Tdh1Xt3567k6snII59t3CsHCMQRKr2HRdChoOMycGgkIuJGDfVqv1jo94UNRTmMVdzpFb+sK4qSc
mveF3yg1OLoewEciYJww1G/ZCuNgpIFcBzdleQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cgEX7tRynX4YnZ3YQk7Zx6jt5Gu/tC4qB62ah30hHuPXs8mHuPEDfzYuv7cwLxBi0a17QcUb3a+u
Epa5sSS8qcjiRKgABTWcD3fLI63hQJ/YytIIsWOG08tOtiY6tKR7F5e6pui2hTTQHo26AGxSJCmf
mMzTQu6fMq7N0Y/npKU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eaTYamZQgmxqe5CtPyiSozNXyLvRADly0AtlzXghyxIqWtTNoj3DlFB8CAASGoBeuf0vmlnA8bP8
YaL3tPNBA4wJw+VFgbKf6+hWLMWOi1HsnQCfPANgZBm9CoKrLlpvajTSCXp2fzTWkNA9FLIuUU4g
atTwqPn4dw8tpsxzmrm4MXziAHYAJ5IfEfgYK2OmU7PSTvPPp/RlXqjdUL4j8VylSqHsHl+9VDYe
KegnahnVOw1DnD2bde1Qsvedo1cjp0TcWJDmEfhidGc2QCw3llz0z0H64O9351v44hdtby96vxF/
txX3T1VA+a36mRPYBykxbe1HXOs2KNfz8psxVw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4704)
`protect data_block
bYBCc482z0ynHwI3xcT/lqRPUGIUHDMya+44fWTXkhX8sEhJrNbv+oTpBpnNGuqbmhLTG5HZ7GZx
kEeeB95dwnZui5096Z6zDzPKOADmPfiWAvnyLqhDbg3LQdVjHVvJf3blqemOY7OfmeKH/YES8CzU
45ylpMwTwul9cZi2OvQ5kSTE4GartvLl7HR6guWM1vgXYAp8uLTJT1gjQWW94+Iue5WBYXW7HZMd
Uc6LXZlbDkXX8ZGIb1DQw+eHeqplqrsm+4IhWA0c30wBzt1f1DrgBHkE4PvvMpc/tzs/St6jCFpU
r8jeX0SfaBUCNtrC+WsF5bULG8IhJHfTE2PCG/jv5trsqvOm9ZprHaG3yuUJXMYz4mhoRkFfcMpF
KGVpxRyc16A4mNAXZdijD4ZUWXSCGXVubfUC0ItTdWQny7PXWJpVjm6V7t+KgaEC+OU6kNDwFQHh
kv9ALVYEBwWAGIdKeziZlaNHyCnleDNRQ+/CbFrxJ8J6oH5yQWvUJnVEKQcUlsDC3Pt8ZQgcrYfa
kof2KgUn4a6f5NJgbhM4mu7p4FydMrh5XvLhfjDwSvnUfuId6Z6p3XT3q1oOUeyuwskM0tBVkI4B
gMcr2SW3zxy8Et+mz0EuQiEXtGYqIsz3clUQCRkpz172zuG0WVXdHJNLdIgZd72cAF49DvTyewYA
//5uzxY5Mlu3SMjxzLeneU/wmozpi78xWNpo4Wrj6IVQj+3hPsuO3p6flXlc4wm276ES6PVxzRXn
zbmRoe84HfC1RlNaa8RJ9UQBd4KdG99a2ysSuFSiUHPL7/64FuMtYZozj/JS1kCg2t7mlgB1zw0D
utN/d52BwSMP0ZfDfaa0evQnTQ+NwjexSBhfDpVV2oi3lY2DSuBdPVYcJN2BLA7q/PrWNQRWSu3N
mPxlbvnRqxXUtaFriKaT4lsOWBOFfGY+AH7sBHUdeeg1NNeVvZA0P0TRgqhZEg13BlCrYhx/3pU5
lOF2NB64JU5SKJsnFt9sOT/XIkDyNH1/Z9OMO9bo3jcDP6ry8FWIBUM1BeUHwvtArFJpa/6LY28Q
jvzmJJ4wTN7Zc7c3kRkZzw6gpsMt0T+JMb/j7XEhVGjoNf/+qBAsBBbxMm8XIVKvM0dibpyazDkM
ShCt8+Nclmmo06UWPyGG4YT6BQVBs8FsyLbqJTO/ZO5SczNRXihI0W4Rn83513AstNFJPmSpe4rn
n5+pUjkKVJ6/AOP/xdnHNr9gjSiSi5jir28LLEdkVgz3UgiLT2oySAeJ64xrAyx8d2FiwIr9/Rh9
sgI43T74id2sW3zvBJjHp8QxJbg6k0/JUqA5IcSKvzbr8C9UQiYRoZ1vFKubyle7GqAyUZKm9Rso
u5BOKpULavZfdn3y21FXdI5G4M+9+c0Tze03NPQxEvhG6bcuvLMROFf6q7egwQQiHS8G4s28cHph
Dit+j9MbaJWbSj1YeiR+TnOsw5lx9NE3JfoDiIO3NaNdmphce/ULIjvBVsadIbXKrDW7RuPFWNH8
FYoErPyRZDveNQJWkVXK4yut256GQ4upwqJ96zi4D8BkfPmwso/xXnzP/9Pz0Ix+Xgm9xmMOjk1g
Hq2QteAV4pP0vc/j2Oeo5KkjAh3cjvyrDzmY96t4V23mUEWds1C9WihVMR8H3aHeHbc576fReQ1z
O4n0uJhXuuJKT9lE9ecM3f67W40iPnTKFY0VPAMiTLfPnclh1RZyPNjAy8b+fXOf68eRhtLPvoLS
XFjHFkEkF8kyUSagVWyNqdrSACdk4eqfnCxN+I2TEDtwiL/3+tmjOi/VHwWVyHPaWTgVwFuFzXvy
Ex35OZWP9C1jmWZL2a+LA7rYOYH4Bn4hqkkWIo/rcORSWAemzuU46tza9ITu4ACEt0AYw8KZ9qKN
hNTaIOxgCNs0qXqZjS317ywWRaR3Z0ivqw5Ws7Su1YUYj9if/3JzBEvvmnpjNUbWhyFdXk+57IMT
H9WATvesiSVMIWpI3t835/gb90kekWytnTlUetRLEnvTf45Q8SDVM1PQ18ucXQV625F2bmuZYmtJ
un6pVz1WrHb20SXQ1ywvGk4exFYz5QWYPmbtVQ8fj/e+0j11sOmEc5RP07/Y21xjewdSz0JDuVDr
hIle32pwOETAdlOPdAeEpSvUbyA7uYgqHYPpcjcaEeOHsIkp4GMjFGSqzUlxqblvG44OSsXXPIfA
VvWp2k3T3YQ2BjlNgJZsWZht/Bzh3vn4VdQpI0k7HJKoSGdjO7+tTu1XykJHLu2hiVGZkuRGVYAi
4n76DohfCsbeQXPjl1ebjdmqqIyfoVQfVrm9Vi/a4GqpEBgVq69c5w564BZtEfccAzGYQqSQWL00
h6iJpoMnJwOAGkTpzifnDY02LXsjl4MxTss0vq2JZf4JCztCtjfi2hnUP+tsJe3puDXfSKHEEhbr
fX9m1A9t9Lw6oN1ChzIcw6ql5IxZhwJdf30xAdm/LmNxl6+AQBBmotHuy0LH2fz94MK91rod7a39
md8HS8DfCu+3DxzibHORhB1zCH6BptU4Uy8Gfoiq9yCXUfw8yb4IUNBRcCNEtRPI4zNKK8XW+tjb
cEZ0cDGk8rNX3uW8PqBX6k8h/1or3Y8772CxT3UzzMu7Totf5KKoDQ7KQQzqIWjcJohojcJ7LGCs
LQXU1yIvHM7q/xz3c5V6+OU6mkwQ1zWghMim2KUU+NmaITxkrYRMud+idomBfI8yB79fgzcxEqg8
rKpudigsVQ/RXt++LGL9fSE9youi2FFfrpWgNi+t9+SJF9L/OrW4oHPBgsJe/GyWhBZg8I45RiAc
51uO5N6HEISYEUr1NUafjPwmZ8NB/1umiUPau2Bn54AUzDyEwp0CZwoc+9+F4MaewHFaw19Cayg1
NwDtfhN3zNqOlLYMpiDiQx4pI8iBAdJizOUORIIsmr8R41RVWbOrhKtDsTqr/A26r1Ctl60h5xYE
B2FpumeCxQNZr7bXCHbjy7G3y6aXEwZI7RuvjWSwwgd2lTsZcdItl6804VVcNDKLB/k3oZZNPLMo
ntXD/UOZBGnydQQzA+WBr4QK5ltOb4tMelsmO9J81C5TTZxEEsFPFkCvGvFEPBkgqVb9pFog6VZ3
Yknjlc4TuFCAvwE+jjr56tXaPgoxAh2v7h9WA50jn8VODAqVrbys82hmCLk45ynmW/Nuin7CAOk/
yMJuZYOS8Tx/sOugTaNZixQc2syVSj0DMcAplxN6S+/mTXorWPiL1FCEBGX5eB+ttFY+CWM6U/gj
OOR8JztGU9EL33KedBa6OO8SBp0U+ikw0aDuebKudom5DoyR5eW8Ze2jkPtkjU0XhwhXYc3o5EU6
EZXzHRdJJ/dHH+A92t4AOQO6VZ3rgXuIxEYOd91PJpQmQWoxRBUbzsmRGeK3TM3DkLLniKxXpqnh
WYeIoFMDvUKHlSAAEY4vT4QLYOzm8Hpa183qU2EhM/p1abX0U8DdJ+zA4paq724VsAbykrpNoRme
NVPxMMkc5Ccj/12ok96qaLXUlRLeniVKMyiKpLYnq48PDHF94+6ixOhQ0AaFBntsqt6IWAefyt1/
EZbYkMbg4mMZdTmq4fMwIWPMJ4Bh02kXTCMQavb/ZpQFPqk6Nw9fgqrSVBbRMkOgqwhfXF/tOO5g
12cblr2Z9oC7icsDVm17mNnNukZtJn33nHPobEBTeadr1oGWBz9QOXr61nB6qaYHKiWijpj0DwF8
xW3Dv0ZmbcMDqxLbGtVjPHMnUYH4/OWV05ZqTzqEMBXN0QiFUw0WuByWGZlfV+gjhqEDjjC8btJm
Qx3YD1nW0mVtJKhjFcHeE6yxdQJCvl/6jgvJS5NS89YEL6qJ+CeaEGqTlJn/Gg2XCrjQyavwPQMJ
evktbaDinHcLvx3wXUQpQrrOlySRXw6vPL5uchrgbr7kfgWdzu7FcDMkmnwKfLYJA8RQnlsGwGR7
IcZNL7Bac1rxmRzHGhRvmY5WWQuaK9G4ePCYPozKWgzGUnmVze9IyUpNd+uOmTflVFty3P2M9XZp
xnvl1vbj7XUnaD/WKV3f7hKsjKPwMEQWu9wdvqq2AkSzwMZ4rVKYbOst4/gIvPIts78hLZIf5Q0X
lKhViMuSN2Fh4YcnUIKcbKKtdIkfacdiiT1uXaKi46V9WOO/IMRfBlA6zkAmUPCwkbk0sF6UnKct
3fih7vOu3z6gu0xaq0EJRYPCtxoHpGCOdarpKTCrBYd5e16m6H7I+f5MiCq9lQYbbgckAeouS4sQ
97BxDsa7oqL81Dh8J0fuNvNvnvYRRjqhKpnPeeMmJdnPdAoyRAGcGIvfOyUEwehm+BV3RmaLImeu
vTIZ/erefJfuLC16112PF0skDKV0EgtNcLF9yzGPT7YFrZPYGvxjqVYK2tDEkaWHrk6+kts0RVsw
iGYd4bmliHX9dRgBWrbmnJY6LOA+vGUTv35E2FkfvoQkAD8NrTQDNmphgrjv6z5uj8ON1ClnhVxJ
pc+L9i66pEnDY5KG2TulOuTI+BIGWseD74ONmwKCDwLND2+Ha6VHivSCohx9+4nOt5NNHfFK1ecG
hxuLDi0cEJ5jruoMzY7lyRu5EB63WXyINuoJLTr70UAEFVIxFRW95s3wEL0pz++GDVyf7yyxFyi5
IBdmff3ixSg+67BxPe7s61HQC8dt8Z3Yz7xZVVvf7Mx8Tw8bSo7J6snPKgOCdHLqZc9x9WWejWC7
4UCmveUbuwspg2TJeNCoWGdFnRle7WfNIKS3Rki+8YzudUFWSgz8lw2GS5vaqaglSPJUNoOEwVB1
fGorYN0fsvwjIUXOnYlcIywbSTw31pYWF8Jymz+9PiDSG4ybw8Sve7Xx4GLhzUvGqvKJAXnT5WRO
plRxk0zi94alSBRk86ZvyHtpkDMSL9JikeEZkJusSFvxjfcbO+sORN64W9pqw7NpKsSbJ3yxibk9
0/57u/vQBUi1Fp5achspK+Q0UtcDHDVkL9Y3WHUvvzgg1jzaEiBXS6YQxUvpr0N2CgpM69H0DkyA
WeLAm3bExUUFIbILI8A8imOOeJ6qXZ6ux0klLwi10OMcyGQMeNV5lINou/EIu7RCcnwD6mpfE73g
Z1gP4jL0qAir/3Na68lt2fV1H4+nB5pgxbn8mjk0h5nCzxldKusNUbyrDhSGyEC3wXuuSHnjZWNX
cmWQ6VBxhPSZp++H75cGN4Opt4+lFeR7ftA/yhlEkoWjERGr+dM4Ic0p38wTIKIOV2MelWCnRSPZ
QewQEOyYke3O+oADiTVWYQaw+ye9rZBsydSGylxLahBqrkOe3oP1hvstfoPtmCsARrrkbq7tBDTS
tR9u1HoRr5uYie+XqHdTY5DxpDNQv8XRv72z4BTz1wlP9X2fc2lM9M1/uL8y5rQyOjfprNcFs+NB
5D/EDe4SdEZvCi2XixZqmEwdG0mJm6BHosuWgG7UGhV1R+oJfHa0z9U9/5Mkva4HHMq+ZG/YRNuv
gAtEc/wHXvNBm+LfYeqRpL6M0R8DBLlYzL9ZlzxRufAwHrKUsm4wVHtOGyn2L7nugcu7rTIod6Vg
QTr5HVnrZOOVIwByD4BjCmEYPK8xkCfL4zbuDRqlOOwZryaRS+YIRU0RA1yIIs812f6yfRCMQZAY
5TliARXOu2FFe7DJk+LwQO1N3sWT90Lp3QNvuaUkprvAcXYwDMtdZTYvMV6srYUalhjl6XIYnrgJ
SeEF3mWt5RAkJuE3PXMik9vbVh2hla9zk0VzEmxh0kKp3hUeuTMGJIO+Ie//gwqBRSaLXjQs+3iP
y11SgOjBBJ6yGwdkydp5JnQta0gNdSW0txvXgDSfJq6C32t62Cr5TMDnetpJFT2FZGWzlS4ccLc+
iAoMYZtGE8kcGVyGKpcfnAY/fMLjuJkHbGNna3xf74mQXirAH6NgxQcTa1f+EfAEiC8ddqw5Nnq+
owHCvbHUDqdNljr9cQwE5SEoI/2puCnbBFI73vD5eM6hIxy1AsGZ2+7tFPJN4FcajdxcdhXVuCop
CU2p0xMsWq/ddVvHa5/3e6Qp5qS2GseUxN3FxQ7r6/vSTbXWcxX/jjk1bna3ek/2BMLNL+hAyUtu
wpu0Ask0ldmX4GedfsF9KsADYNxZ9buwEFwHSRe9ykWfb0bIFMpy4L5Zhoetul9Omu8j4cy12AHk
lLd8iayijkiojNwOtZVxLdNcmX2WxXYGVBO/M1ON5Qh6BFf542pkyzEEmCIRJnwqsSQzVbsCDEru
p/1VBgMvyAr+WBnmNQGKS+T+/hCGsLX0B2/Z4mNv
`protect end_protected

