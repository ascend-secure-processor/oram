    parameter   NumValidBlock = 1024,
                Recursion = 3,
                MaxLogRecursion = 4   
