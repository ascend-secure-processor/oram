

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IqsJ/aBz35K24t9LZwiyL+Wn5yoWfTFIEuxs9EhFvCxLyL1ISGvv4JoZej8cTbfJJ8xMt0gqm5c6
/ScCZ3Ek5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Krm7WZRF+mn4/RNLJOSefxQ66KzZ8dXriLS4R6+PVBwn7glFcM5csAM29K4x04+ZJ9arg9+FCoXj
hOM2Die39eDxmaqjn5enU2ENA33CDB6OF3Cy83BxLmdqpLNGbeiuOr6MocsM5a3j94X05fQ0LxsX
8/EZ/stZDMew2exXSXI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ckKFZ2pg+rP+jJSuNGYaQBLJy4rnXh1i0CUulzPO0+hlcYLZZfsQV42SzdRIkwP9HPkH0XLQ7PIK
FmYZreryk65+4YEQOfngxF+uXbGat51HhMyq6XYqnVuHOo97ynPUdFzfsz+CeCOQYQ9m3r4Rkgq5
dC/mSZfTvYuTwPcvu0CdadIV7AC+V8C6GIxn5RYNwT6lAS8w1DHLOfwLJrXDd7x2VL6czZhaXriD
loNoUA2T1oIOFhzsP3HtbhuENHrRWI5yODiPpQxSEXe6oOQSb52J5JUrqYWl5nwrf7EoqKKkNM2i
FaJF5ZS8kxC9ORr013bOtdA2rRz5sv6l0YaHPw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CjHaz/2VemQNS2RAIhpRvzp2G7t67gEPCT3XVBn8mFuIYm42wqeB1b0mTBRnM8IGt8/FCk01OQfP
V1q/HI3J7pJIAFvKrC3ixpK4X+PErkFp24AovdqHg3im8mtqqnz3C6pKRTuQ0v1eyxhMlpZeRWoj
g1IY3e/3Knf5rrK8Ias=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Barjj702+mUlW9Wk75+WrM3JMyhH4Dwsk9sMnNWciixsDZmeu4KhuyQVO8UeV0aMmwq3CAC1kxY2
j6/W025m2yW2I4FqMPnPBDzp3tds+GhrpVjVAszsZhyjjKHdGw2ESGgMXINL7BZG2COhKxhMTeT/
auMHzSoY8eG6DdP/lCA+Bir4lYJZNnfopUkZ5bN5YksJZNQAXnxQ5k4CbSQQXEp7R6NVOS10yPMf
gsnCgUSXUHusBaqHhyP0omZEtpfVa/mBiSOrIty8lH4J3jLwsV5lInMF7ztDXkGFrtuy4Wcd/fOQ
uk0jXt9/UvxABBPZYQzfVmcOw3xOiXWJDmktyw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
aKDyvw9jTNvQFJy2UdatjUrXCg9ut1edCBBd5Y6DmQHOZrE8M8Bk3r/4ey98eb+89T0jgeCddi8L
QmrFLCiYGeTNj9jdqhXvXyYwvYWE8NL/aZDLSdWXw1QALVoGkYrWLZpwhLr3AL75gnjctccWEji+
vRbr3nVgT/dyX+ERJDmnbC8tKvXT7vqopsq3QmqQYBOTQHeToRGSWNATfcVegkJoSiCY4EzjkiyR
RFdQG09jUcRX8uuU0lrs1brwLfUvuZ9xqkzbMsfgCWmDwtb8dmmeNIoX+OOZwt0p8MtJV6Pm2tex
/GwGlMN2Fgvq+ZwIVREZoAze1iM+dKeKqvAs5/L2ZHsQHm+tYDTunyrulUlnUS3tsePi7sqlwzPS
xYsrosnzRJlTqV4vCZY6T91xUdQpHqbnVIyVkpgBT0a0kd97Na8oCGcPTL6mi0N/4OezaD1ZwvQ/
BBy44fC531qsJSZt37LI7w0D5y4Gx7++QNRkHOCAjY8WIjiCkV25cPu2CR3Jxm1Dtl9uB41qL16F
Mn0HPoYI/KHSMGAKwiLB3h1UzTyIjiLyA4Xjq2i+4n5n3grIhnjAp+P9Tqeg9mPctSj2IZSAsRek
Guhmxf+3N36WcUo3t0tCJYO6oYL5l9fN6elAK9DT+clybFDQDezIuujDTYdy/bnSlzJZ9emKS1gB
WPjS+WqxZCP212T7az8VLEY1D4hLqHvA2tokK3v/W7qZ+hkg17salF04RV46HtYHDkUy3SBp6Foq
TIbsYW/uWN94TPcgup8CPitrNJndo1Uae3XDnYf3Jmn6w4jrN9ZUJDdR54KcQRmLwL2Y1NUkkTbD
MYgLVFxvyWg+lMqJbI0kJmDZGjAikETAV95wZili9AHho8K0vGZC3ItGsDUVb8rGazTqU3naf9WT
0vsIz9JjTmLwuTNxbuNjxs3xDRx/EfnBNM2ZN0C40fn6iKUc5+OpxLgzZzQJrj+yb9mgy3FlaNDQ
Ba4jGtNrgYGtg+rv/lW1TdJ9RqOpc6uhiLdA1YKx4zwoIYRG1tVYswhsIdR5+ezNxGntePYy8yhq
DUnzL8Pircu9CyxZqCXy5qQ51R9BdsTISnGvEUzdb4uXl+s8yB+Er8+JHhtXZsqztxnT8WA67p78
nJMBh/3M/gkfxcQL/wDvpLZmvPHxXyht7HjgRbBCdXWZZTABvOm341WniLmlhjG4AYiJE1hB7BIW
OGPa9jYQfGhQSaoQIAk0Nn+IVS/OhFog96EsJkRejiXdXBSUIBJdm0ZJBcIaqoOsG/44h5txsVS5
22oSSa9UM35wxAD2OVCtG9Ih0C2AeMzHip6y17gU+CFL3AVtfTzLkAsaPvaIGp8GhOQZHdYtl0qC
JRdj3eeTXA7EE5emIIJns64sI3EBt75B5baqagYqIX3G2cNLhobw81u6LeOQVYKtPhiwHYXxmMfd
tQ9tvMkj/OCyzXs1LVCz4591gZbqiS+G7OF0pFzwqwgzOzL7A1cERV+G5KFOgCVbDWF6dhjXqDsY
1u8ToKPGBhF0pUDIsGmt4dwhzzf+2jLEVevXzpz1FuvpkqD/Q8k41nR0tUAiKG8nnEfdlAiXdeX3
TgqRNfQXYI55s7LelDZANLjnkHXHXiK2woSg1EFsNwYRoSWDztepPKBr0f0L7+0m662pborfyQtZ
npk9i8TBMJHkS8IChKLH38RiedUfUbKnHFrZSLDg2gH3x8T5RXMp8j1AcuX9SAu0To0QIC0zkDwp
NX1rfzQUxf816EaGyydOR02iwFiYYwKUptjxtMgFrAmWUTmHBO69ns8RhuvlNEkAnDBlKgYuGhJx
9g0Vn2RInwD34SM0HbMIEx/SCg6OMZ1vMLdUk0eFeZwZO4752m/KTYKF9WiZx8+msdl680SFcqRz
4Yy3qaEWtE7O1dz/O3LuaRcZFC34aQ+bByZtFvsmnOZtQCjGWAjZmkc+jOANOsJnoY2SP91uOYot
ZhcwPWQfJW2+ue6oJlkE/HypsSwRwIhajTCwvsJzzTJAFA9mY+ELepju1KsGfObHqj73aoXUXzjh
YxUmIFaVUvC8ZJzNn1JbzKoRNxARIhy+pciaPiNojWLrb0BauE6R0Whkw0t9nn03AUBtZEfIZOFT
Uv04+UeGboO+VqGRz7k5NoUcxfJaLPwR7FJQ8X2R67ol2Ht/qRrRUBThV2SlhtjW6b/aewrweQ/m
4Jft0uGoA+SimuUxjlsqquqpqm2/S1FJyUtF95YTavLPnWy5zZ7U8tgRM7+EpJZQ2ijcdt8vD3PL
9hU9sXNb4DZXTMrMLtfOInCVUfFipHANBFbBWV3DCnc+gteSJefRgpeRHmllwBxY1zt22SUFC9ae
QhPbmlSqAcdWcnX8dQqtXHt1IpSArQ9xnCbwZhmlsy2Z2Tw4iVCdvModmyM9QPF7g6HMX/I7gRwG
fioaEqFLt6ve6JJ+WCQMGDHOTfAMOnh5MskeE6Su0zMNgHnOjF4hQRLO83/3wKuxdnH69kejiIn1
VfVHTfUIrMtqI+82NESXZyize98gTGxvm72usmrZ5wXm8I81CkYHxI5AnuhFdTE/+tFzGynJPtVa
9J+DfuJjcwXSQIcuftCju/bAPaH0u6seEUBrgHRCCNIuChbW4BP1UOTVxIYwkGyzTJDjRD/v4//C
JabT53bInRYvzpe37ViERoQ+ptwo1XhAgLvGz135YvWwlm1UQyPhO6XwXRGlLklsdsOQxJTa890Q
9uPB9M3UHZ3rX7rjeyI2vZBEOaQwBU9EmR/P/IpyEdmfsYjLutxGSFAo8a70t9gJ3E8jC8xEV7Tq
0T07D0PS84uAm3FrOrnnW1wmurJMT1bQXJQBMyg9j2c6nCbF1/yGwsetcaWzQnCEsBH3DMSAfr4Y
leaGKDWIDYBp7PKIX8DYUxgnDYLDP8J7jOCBsCTEZ50qaMPECMm8l7Qu1JN59Hr74uwXTH9Nk8JU
KMZ/N7iVjqtvDSK08TuB4dLhWjXqexrAjbu8aGcBmM3PlHx90+jeqsDzGa/RQY6BnVnkEJ1FpJej
wRuSpeMVip0oMkQfkYwLQbe7/4csnu47WDSZ8aQfVkTV4AlG4ZLwzZk8G4oGTrabGA9kEVAv+U8V
Ss8lTI3yiQDK+1uAAg0J5XO0ajh+9d18/b1kmXuj5EN3elmMmGY2UcuiD6PoIWVR/6hS9S67S0bq
fIM6FobNXMKt26S21GAu0lRGVGPHUiWNoSaICAkf1WNInDh4U3Z7hBiYepDYjJIX9jXSzyh/Pq1H
bB25rkmQtRdO+SfDI/T+W+mZbQtQQYgfBGk303Id5nqIg5YtWxn5inyRPJfHY+p3HI+LjULog2GH
XiL/DSauOHqj1r5DABFlyu/PT7Q9MTUWos5492ppwv40oN87CZrp4anVYH8R5h62zXroNI0Go7Lz
S7jg+xrJYkAp8AKBZ3DbahzGdDTLLYfQW7gqwSRN9xRR1dIF4xkp4RwJQ5LA0Ey3/jEYVJhIdltn
Zpu073G7hqaYTfOwCGhPCm8qeun2RTVXKylmDivSd7OQRDGAlUnQ8Z/wmC4+44PnGwm1YLWS90L7
uek21Y6zW0ngUXFy31WnRA6sn6HsqVVDYXrMre5AVWe5E0PugftcHsOk3Mjj8hhFC90f2TXtABT6
pazn69PMal+UmTQYzGP1fPRvjGMEu6bQ/rieu13h1BTHIIRpkXjmfIlEZKfmya9W5l/o4of8YHjO
HjQ7IFNM4P32Pxrr2ErDhpDdsdeJrhahSBroNOB9FAkA03w/120gDrgy0c7SQw4ZxfnG/BsH0NoZ
y3wzdp8yWQhMwhBCTnsYBMeT2enySEzsHSEFllu+gQB5FXRviiD8OAbTzBDzX6pobSOZ2He6g8Ok
pyzzD93xamqS4CcReiWNNZ6Qy1tr89wdvHfzvZL+e+F7icPz7yToTt/bB42bqEMVmh8jh5rkcxEy
3DyRGpEMmALTy0zZmXV+cz8l1u/TQ6p2LPLzOcQmFcq9t3/SwRMknkzDja7/WrsGITaOazPsE8Le
z+5vK8CXLDl/gnFT28k+4Ri7MphGlhXb9B2twjAaebpPJhLp693q+ZEM6PoUn57qN9Gtq/NthFND
MkNXYEMGQDcDb8BpVIJEi+vv4AWEOU8Dy01ShCmh+m/D40iFa2+KdaTHZ4yI1U6nWG1zmtoLpdRL
Sgzy/Sl4kst4LFfEybB97nF2FILTKpY9lA1JPiKJ/6Yt2fllG8vcitH2T2jCubFb6/5o5PS3VV7F
PU5iUqX2465Bwe39KLvfiM8HBrZrlwRhDNTfZvEARHlborkdDFAkAE4NWRZYWQ329XqfmTc5sL6l
yxYXTLtWblXPZNTn8bFbqNM5dPS0BkrHqMLsCabT7DeC9ptlwGhIU8CQwQaJVOyzEfFVg2lCF9cf
xeDvusE/JYxE53LFVr6qbmAYyXXSlcnjNpMu6Ox56D/TOd4qoGCsz3CbBEcXDHffkO1yq5keBWht
jrD93e6vO0NY4EQVO2rqDs6FZDhMvk909Lt4G1gA0nr/wB/dkbftn0PB0bVzE4f92Eipxm6KZAHp
ehDah/tI4SkFQqiNxSWB+17J3CO9/faIZEFCJNdjlr5huL9SWXn1fNYC5aMb1Z+yYKZJIvuM+CNv
kw0zX6gn5DA1T9OhfMf5JmzbwPRMmWx49uZgg5EgqAEEIQJqZ1wTeQxXvSkA2wnSqkSjsJK93zhN
F692JIkGJL1vnFdjRpEMAvUgwxqSl+dB9vmvUcaKYp7vNzKQOVS6jGVojOAhEJ1s9ywGARFUKS0j
tE3adfsWzLRIYABVuGDNQIN6e2y+5sXaw7Y+pVd1oD6rlCggodEm1BgQEagMbFHMazVbH7oZQxym
kN34pStg7sYfX754z6Zweg==
`protect end_protected

