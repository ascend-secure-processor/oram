

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OP+KjfVRZreasQPIncWQPmPZCt5JFWhIIy4VHjaZxj7Y6wr2qKvywHjbF/yXodNxHFYOy9sR3vAp
hH71X9VK2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mnsLcCIynG9TEe1wotjZ45CdHCA1MBFRwPegXXONgrzk1QXBupO65Vnscm84UpyxWv/E/UOw/Z6m
Pf/FhWz7L7LOInTR4LTQqP4jjMtGlWEJjxFg204XylszXVmXu1lCXqzI7XU8izUjYa6qEci/pTrG
uy1jgMWAZ8rCB0EyheI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B5honffKRyTCPFgC8h5SSIyg+TXvDcf1J7FUQ5Ne2IA/vtxwp9NMLD1BefZzHdX1uf4H0Jx23ELj
NIE8A0Vhe37jzCRHQHxRJABSQ3WJUfLKT3Mre2wQAv3wS+SWBv7ZJtJXWfdqc20Gytb1eEt3UYn2
fJtMIxzNxRY9eMascdgF+pRnoc82jad1+ACEnvp8o5T8cn4yQtJq39geJdlD9sU9sBGuGOmyIPEv
RzBNT81HUvqAzS+oO3VRVNBiKBgyX99Z8iKJv0LV6Rs3VWCHucNnme56IChiJgaKkU/pn1u7LhHE
zv/4JuzIspwJd0ZBm9BIe9lqyOqr/VS5Pj8Kdg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z4vWmjiUJM8lPsUoPX9Iz69piUYkVaeKiIlUTC6Po0g81y1+/kdSwHoTICqOsOlrho+30wlQeUcc
lOOj30uypDyt9vQGTZboHLtPXag8c5Wfi9gwTtEJ62w5iMRDhXWRz2TXUBWIBvLP/Z2N98pnK5nT
SR+MY+xMYUxhO4PyvRk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zc3yAKfp8yBwKOmxWwVMJBBil1Ug0keq1tMd6HBvZAzoX+aBLSZRbz2cRmFNvxCsvfdeJ0zUP/PR
z6600GLE6sfXpPGrueSjV9GuJLKHitvDxOICOmHYDias+BlzwEWLU4FScw51eam1o5P0Ku5Es0w9
ZdxTDAjr9Rov6kEgFq9Xjw+oK6nMOwBdgqCpoGcx0m2WFgKBhVvP5ftOp+x9TdF+wxihznDgsxwf
AKRNiMxg5/MiOWUSL04whxGZ7V9IkjqeeJBSByNQrfsmVecOp3PNGoScSJV/M3xLwf8fl1yqf5PU
3SFUExMzKuJasmUTXlk0r9p28So4NLOZpltxkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
LkOD41KNqyBRoQ2uhcITU6umJ767MadLYrWwvjPhr4mfakN7oQ5Ty2JPZGXKgSbjwe+NqUez/XL9
Cvr5286ATArBcu0MPScBKgoR0IMxs4lUIgrGCO3T+MIvajO2G32N/3NbyxTm0ooJSxzF3HuNQq8t
Wh7ywAX3C0+ro1kbomNTlXtSl9dHWgXHGgst9b88uZIdKAmgVGLdJwKD7+kBBpg2J81+mLHzfedg
lqiJ18OHRwXi8aw1jIO2bnYwXHowbAS0cdcY/sx57TtKozqoq+hIZK6IfKQKj/jfSXIPBlUxqbsx
uA9X89xUBHjNfAH6tdolW0FuR6mCe1oNg3f5T+PsGv7W2F2CXo5gJ6HezAMqYZxeTnSeqUS0ZC6A
GgVQMH6NA9bVj0dnukA9jXFzu2iO1Ej3IPhP4dmJdvyrTaWVmjXWWw2Qsv+ER/uJgb+dFGBBWEM7
727dpX21KrmGKgofx7ocI2L7OLM5V68W8XfcJfyvlo5Aa4j1bovMGLiN23B+NdeIc3h7+ezMV2LD
dYoqz4ybv0D+mcB/TqbFdZTQCVQL3oYeqMp0TK3VFsr5Sh8Dxx7G1aVWmUkKIvVrofH4wU4UaDp1
dUV8I1mCL6x1HNia7IzTkRHyq+jmMp0Y3WJi8rXddvSy3YFV+yY0xeXEPu3lGRp3o2RF10izi5KE
GXo3HV1mDlnG1ZpIH8pvupsVlQDsRFxKTMtqxShubc0sCrwwIT7yha/r9bdLvsP1Ksc8MUoSeIhF
8tiMikh7g0PyDRBKjst+zm4O7s62TOyIQOPGa9hm8Q7bQM5aBNzSkkQERkkiCL80YLtSsbxD3w1Q
DDt4hx/pZgBaeu/LY2wZf1W53JSuU33VEcYCuy4R0ESBJLRl5lm2l8zrOrrOcCzkkVKEeAEdlmYE
TAKRKRulFjtG4b4yacgEM5Vq/TIpPur8OTnoKCkJvlA7FUyVYjXMY3RuCFlfaAQAtW2dvC6fszgP
HJ/rZtLcICCkvfj5AvUIuhdeRCOy1xN+g5HbddOK0atgksMX2ckYu6trzBLN3OBovK0DGPTmR564
9p6eauCfDXUn/SJgten4qykSlvVq+XPEy7gpa2/DT5ds9GBO9bDNz+dMSO+mYZc2EE8NwCsWl76r
pheh0ydZuffne8CML48UX3raGPAX9U+TBWidNXwJaPxuJG/iZn76MVRIKvNXISqm0VTC91RBj2sv
iHFvAu6DCK8lWp15gM1lsOWmjB3/1ikqwIUYAjrji97qVyM/UKwwJfFJZ9n54jp1bTn4Us+LS9XV
0fx8F1JoDtCZ9Mzq1O+Y43niYFxHrWV1b4Plb4/eXaB2+EKzLLOSO7JJ1mgxR8arYh/yd53iVroS
vJ6chqAyyYHnunsD6EgTcwXY6Ixo/1RzzMm5OZdZ5W/kUi5OO5m4zir5T6TfJARA3nnGl3hVHOSZ
rOqozaysNzQ8+zKc2XmubLRNw8Pvl0C7iVh1UQWUo6y0q2sAvTjmVhJx4ac42K0LcmhIg0z94Hdo
r7WlM2A6yZjEG2LvZBMwLbY3XDV2xZ7tWqxVo7RYr6xCGLc50TSxNQ1RS9TkEPHzXTduzTiceYqi
f4vn2FAc9dc895e1owshb67qMhtwyYb6LWDS+V5fgmkVyRNqGei7ErjCu0JK1Q7ikxbGLOaMJvun
KyeJHLMFvEtAdhNzTzmqOe+fYHFyl333yP71Ha2+VMP2XxyTdHy52owbEGBLOri5pOqHadMsOnKq
DlVroEqsdjxtyUlg+lS64SzuYTaUyxc5WfVyTWyxUomDRhRniuCar+4/rDROo9GGsSEwPvZkUElR
rwAJ+83xCz+4CngyNdarTL3VAnY0wBaY2jufNS4uIftm7ksSB6qnoIBFgTbKEGJVHsFaFf7VGUsH
zcn2+VxxaHFU+ZcensVSeXJtZ7AxKfsLuMu6Nev42ac8hV7b5ZN9XZYTZsdh6XOsP+B/YUsccaV0
n0HvlS97L+yLX2heT21sJ0PnHXUvpqXYokfMfV0G76igxu4e64ornSbSKzRca8rpntdFa8g4Vgt4
xo3LGkg2ZcelNOFawKd/p6l2viBA7mO6t4Z5pk5IqW1rNBEKM5/m5s0C/jpYQHLldiOfprm20z4r
d2k/awQCvYADRhexWdILREJvDdJ2QkpwyG8GUU3utISh8CDZXJ9K7C6l3ZTOa465evxs383bfQ4n
Wk5qC3WmMiG5lXIXETGq4qIE22cnO/XHrrYuPsqMKSEquYyydUYqlRR+GSaS9AU+IXUOjzzPvTD0
2v6f6KMIrHtAYrIf94n/WC/m/MPEzbP1WloNhc6Ri90Tj3gdDOBA/5n6gKcxdOH2hH4BrlcggIhH
Wo13A3NnjEwE4hjYPM+/KK4Gx2oDiNc9zhEx+hc3W01QOBp3w3hVuR1wpYl3Lpj+AZ+5vErTVsdF
RwsfKeDlvb4nIgLk1MXx9Wiv5WMX6oTFbvfJ4cdppcX7TAsThNOMddH/I2OLKIczBrp/xRnSTXgB
m/uK7QPE7YkDnHVnk+5nbHukwwgZt0PA2jLRIfOYjfQpjRMGNt+M/fRD1Gowyqalp7ES5GOBJWME
NLheyotTVZQlkQwF+zxoMKM+H+1nibDZfYbgC6TwuiRxeVDRMmIyBQc6rt0rGIeo8fhOhZSezLkl
OJtjcxlND7gyL8dKZ5wOrSzQrOa8Ghzf7y6D1eTbQhNAeMuE5HwjVoiucT0MFnJtC61BEPwPGmri
H96pPCR2fBvqb0s9MgjjlrVZdcIw7ccBkckNNGw0hJbkNHuVGHUyZkwB4tFcCqG5R4JdFsfCBs9y
9Vih7pYkhkRNSlJuryLEYeXOxlNL/efHK+QMhV0Ju/3WrTsfqFt7d/nPiqWHes0i39mqfdr/d+2a
jaN/yr5Z8VqTVWi4n/THYZ2vt1/IEPBO1YHs3u8AI7vlue3yv5O6AIHaDhVUJVm2bo8cZY+j9jPT
koLyEPSReWsu5wTsrTYTiLS1IEgWLXMQ2jYpvAzNkddqRRZ71gL3b3/0xJrK/5ROsGBDCFHPcZDc
+FgpPM+R5U5ODalSWd2xebXmzgdNY0UuZ2mGI4yY/kRGsXOYgTRcZOpEaSVxXc+Y1NKTehlEdrN/
t3xipbE/9xNZ/qpRddj18zgog8gJQWTAmgaUb3VmHE/ZREhEIrSVTB7GqDRe9odyZMXlg8qw5gem
V6mDPC1WlwC085lfdW0cos2eEH9mw/6XyALvseIiTxCthX7ze+8E/AEtLmfyfE9iIDtdyfWOTDxj
tvx6Tu590ZsM9ILb+qNXOMQ62OILihPSH3Jzt7ABjw0p++ZLfaTcM5RhRzRN6UGnHNphbpef1aEf
qBz1BWLLSioNlc1jlCuk56l0yz+0xjmxKPm247Rnls8oSpIWKtqmp+nzh+RAaCnI2w/39z7bQsKJ
FtRDL3GT34zUDQTdxr5j5dD2NocgtjpndnivFm8B7K3wyNuDanhgewNaQiWQMB3ct64EDsqiVSQe
Or4DXnof5EGf4WeGjAT8WdGnAboT45cyCWpcfxnqszU3mEqPjFZDntdo/8fnWxDT1P0HD607uvhb
4fBJZNWZ2hQplaqFsbflaB3WzWpYO8i1Ck7oAD+NvT2G35VTBhHzglWVs/0c6xZJ8hn+XgvbksiN
UNW54TgDpl8OqHD+eTvuKDqDWeqs1rd/NMEb+nfjrjgFPYJJomt6i79meeMgGX41Q6wsLdS8jvxV
OirjYlZOk/9PHkJ8+XtvNslhNgM16IKCUr3TyKcXbE0YXkn2G66CmFJJ2JappJfVa5vyoJEX6RZr
XNkn7rG/vYbs+8pfmmtcuE0Z8BUt2BCPWkk6TmCEKarRFGSUReJopkZCd8pprWofNIEEAbCb7+fe
xLOSvK5B46M4baj5YiWC3uRauJ2YNu1xLFp4NaNAO7jb5aMl26tKSrY68r9CocscstIy2GVSdDmX
WUw0VHJoovZYSIQI0SXCMxZf0D8tDehG6k4FzfclLTFt4MocbrFppEQwnjzxMpmHkcAREQ2b+ooD
vJtCyZeftpiB0pH2uVPm8NJCCMCauj3nyHCvhyzk6vLKxollxj/Uln+NYQlKwf1zeiDV44I0pR9t
HtxdLBiDxT7FR0+yO5Ec+3thCaYc3zIfAQXGBigvSr8f6tPACoeGxyyj/H5GdULeksbKaAAGoxOA
fwKdgAGqJRXcnc3Xz4PzdT+Q5ZLJzfLpeYqHBVScDLfB2f8aVAsuEmtm204i+Z2Zu0Rv/Ns3rHFS
dAn9M4W2bq/tEVLCXhbRZPFczOlUlMzlzloo9Mhz/Pis8WCOLwG5kOyD93J0EC1MhHxs6RKxfeoq
b1u740DS237aRVDCAnuPa8eCvsE/KDE5GIGs1agvYInoquAk0UUOE1d69Y2nJZWZAndKuq4Sj2qZ
eaO02bTOEDJxzwrjgOyqU1eXtvpIkI6mWBjeReVk9iFQCam8JwPnj3ufzUDcA89B8bW+WSrCo35j
TBdk72e9Shp2QmdYypYW3av6cyA6XbL+I0Y8X9IE+QdmYsJSfNdcBzu40TauJqhUT5X5pRSyuGCe
18ocjj6bIG1AOUDdDwCrIY+2xB6aVh0IgIP6ZJ/M05m/pXmHh0U/DPVyRI1BuzKNpbK//xe/Lpof
tQTcIrk3b+e9U9RZHIwOE5JWpZ5/qOQCKPw5dfU/1/91Nl/JTcKW1S8Mtxt+Q7I4EpsgbCmYPMc5
WogzcRZELmONz456Xw1fcjSGtsrVr8+9LC6pf7cXvDIZS8UIUKn2BxgKEDSKPG7GqetR/rXFAj4D
xv+F6cwyEZAW0ffQg+stYThdVadbdHK01dXMXrQjeMGaC+CPaYj+MzNzGjmV0eteil6aSacmK9Xs
7thA/NKjOXzHb59DPIEOtBkXihtCpyIyjB6376EWCAkUHbHHboX12AudYl91bCgsUuTQopj/TOAq
o88o8Ejfki1pINxkIyQ6/LoZU9W/griMm7nhTBhjmeVE8uHrG/uBemvbqtXc7OQxkFbrcLD5GOVk
NXvJB3on3xLiTgis23V3yUTWwTFjU+832rs9l1QsamjJP09i7ovX4gd6IRnGxIBbVne5RQQPAABk
j4nzOezhWjyDBRhCEMVbRwyDFXJ6LEaKHbxLc763LNQCT5nC6y2ZRm5AprwP3jU/AI9wnHIEUf0w
oL70/7+Yc6JhiIMhQJ4Luli6mPpc4nf5j/xU4pXC3WsFRe4CNwu0SY2r3wDQcbfwTk5srRZp+hT+
l9TG5jmNtLjYCdUSghwMFkp+nYB2rY25Yt1CXP0AyYJJSQYUg3BEvNnTw8OoxgoJzTsMnXykfxKc
RQJpnsPe2BMc3PlFeRV3NRJSRn4R9+NYjBubZA34wOp2H5Y8VwbiE4F6pIKL9E6Ifw/QzMFaFVCW
iaOs7DBn8ZvR5ODyodUnXAaztH2R7z4W28sGw3HkdhsCyeaDB8Tl0DCuQGzcalRkaT6DOyQKmi+H
0l4SS+0IC4esCcJb22U2YlYnPCxK/oCEbHgTz2nxUCAR5bma6qILZBaxUPBlMxkguzgAamhrl6ns
MNqt3dfdJEJxu3eJ5JMwJauS/yLw5KZV+DVsjNt7d6QJIydXYOLzgqSoXy3ZjM5+jDshHOtAs5hP
68bOMsBwZdZReuQYgo1/gNtPCqdGBGadw7pZnAhkQW6EhCGQXeygej8u0m4nsihMI+T5IZ1pl/tr
CbzuFeDtCFm0suYLWmq7xI/Yi/m2oMla4vXBvonvjw9Bt+mB4EA2zPW1OJRvTqYnj4sWtV7zXyPM
t0PwCt5r8osL2uEJNG21KnD8PPmkpP0YqcEFOi2Xgc0H6CTYImyZcsDQ8QhIlCWExCdrUrCoPGG8
Uj2WZBPWr8HD12AZl4PkchOsqkkFuzHa6vYqoP1PF7ESqBNWw2T1Coi8CddYVTu2XOcPb6+VtuV3
AXK8WR/oibpFEH/hvORkCKepa8gI/Wacb8/CT6FH3PQpk60dzJ9qTucGPygKtnXdU3V2cuk6FPE1
v2xmRJCuG5hyFn5tv/ixWr0tnk/eZ5+4iiIapEmkXnlMS6a7C5idKyi4nTExj39ViXJ5UEe7l1v0
EHG8xAD4uJWMvMOqpIsRIetfb5Nl4SW6uaQRdGg1TAhQh5UmQYFr7AIap/ZlaBa3micf2gAOq2KD
gnvhxnUg5u+mkrkKLe74tcx03RGDug2maevK9DI1R1ExGzeYitklj0VtMWv4MWGswO34a4o9c91o
8Aw1mnpNbzWvtD9kwvzKjyDMB5Ybxmaq/+FHD7H/26GL2ueoIzKwlyQTYY/WvzYSc8F3p9gDdEG3
n9SWQ0kzc7AiBZMInWE/EkaggKvPRfq44RtumJ5W0AOMQWi86+eDzaI7/pBlCvyTA6lS07DoIBLK
AGUM6bZENJ8zlW+tn+k6l4tYbvdZHSmy5JsiOad0EFgwv4Nhu0lFi9e82ulTGZrDiojyIrOsbpQ+
XqmnV2rtLSdQePistR1xmdsmn0f0zQBYMNp8RiWxjwFYGo/ieMyL4tdEF6ep5F3KEUGG/6ctWIcL
Y3shYlhgwavM9ORXv0Ebmzid1B1yhfwpWbgji5RLdaSS1fhzSrn+d3RDQZGRz690ijD/VCGDCHRi
YIyjdBrjQQ47aghamOufzWuevNii67RlSSPkfbmw5NbfByGZ1jbt1QCNzqccdUIOcFas+F2rNluG
WAkJku49TOANR45ExaR6IA2TJZ2PldIrVnG5ySltLjgMAf+QpnL1scTBqb4U7OMjVslExaTvQFAy
K5JLXyv8JXrhFfxFJFHn0ha83WyXs5QGNuB7O4YJLc//h5dMiLGcHJUTk52+dzSDxwtaJTFHCJHR
CU17nnSVif0JDG8aDzud+phBo2VeoK3O9TPvf8rlL7GBnAEGokBjaf7AEtyLP1MV0HA0Tv47DOCR
JUN3LoU0MuKnjzQPkCsPk28JLl9F9UjyUshjOq1gCTTwj5p67HbZMOQtchyxINiwtR6qzI77abid
jI7BOYOxMA6GMHtUbsBtAD2lY/IG2tcp/vWNF3KcMzeymdknwHWY4hq4wGLB42jh8AUHnyy5QVr/
5wj6zNJnrbeMfMk73tDnmm9n7DXI4T+xGxRo0og9K5X5LJfN7B2iOcJn3BmafBXY6s9bw+xqrBQC
93rlKMx+sIcWyIwhWHUFl89hXW4u0Nj+TIcNfMMhnPPV3PNSLE0L2j1HppS5T6ZpmnWvw85tevnR
uTH7apjyNxBKDK6IVhr6Lt2ECYqOoDkybr2fmla5i16RnQwoSo1zdi6jZ4NJZoA60BL3ER95bCCX
hu0W/nDkHO3vD6sVWzcCMfzGs20PyT7yFfe78YLr9+OKe8IWiZUgNuu8nf+qNI1jVM4O1zlLIW1K
ZKp8Fk1WBLrii4GCZ8+uncwyn3NzQYzyzZu0ZS8pIF4Gz7dYgponLzLulZJgUmuph31ik0vUjyZl
1K6/Ho1d59XZItRcSWFC1z7N740ZSSyalP8+yfrMLhGpOgmJ65IhsjCR9v8zbpdjh57BMS0fxiJj
ZYsA0NJ6mBH9M7LlUR5y2Z2AiqRURp5sOwjM27uc/LFbWOJwtN9jHc6/p37K2Hl3gSWvNzp0foPO
4UfOC8JXqvnGZGsEPePRIAEdb8+v5vx5yELPtHZFTgPQFNaUl271likMWT0nur6bptryq/374P0a
oxq8GwjGrotcWSsbKmdFvxTimk0zJsr2f4X7kFvpq/yWHghOb2vOP/MB6RKwr2Fu62U8NozessVC
+O2C5wLGfGWBHvrzdJPYtJUFmOTEJ2zGxqUDjYAtW9MTAuzxpOY6rGGDeZLueOvE6T802clcmDDo
LDdOcMpwqF7KqneFKXm0v4Dc9JoKHZmarRcct9v/hQxtrbpFLcSdEs6iDFO312gYwu8IasGtD5NN
48YzNCY73wL3Fa5TDNjBi5v97n/v5oaC/tcpBgz6bkJSvPyRvLmybUWJ5VANym7z9CUDiQ4NlktL
4ZF07M2kGs6Eg8Tv7cc8FaStI8jmeFo1VCHciCzUrbUVSSchvOKRvqlRcrtzAIZBMg7lNGhLiPc5
1olg0U3RTfAHK+BJDwt+FbjopTaOgVlHHVE4cFuFKdGbpPviGum56TkPAbtZF4DNvh8l7qC4TpCo
GXs3cZVHgD5+6b+0aMwk0RdboGt/LvKr8KRHqBJP+UNnH0tKi9ANoOgJe4y9edkSrT5THnUPZ8KX
nSk0n9zhr+1KErxeYHarozJZTxAZP5GKsOvRQx+AWDPGyTRYIP12UdLO937O8EHiNb2lHODNf0jY
8gaNJYZsv0aRpjwFnCXwHEHG3cPEIblK80GULFvKAz+wGeI7BmsBmlo2ePFvolgXM7mPoKD55WiB
6rhBi0FZIN0LPFJuy6ugMikuo2/1osQ5tqCUw0yoyOlJfaBH5pdEqaUMBswFxP21rOI5IZwdLbbE
dxMgPW0zkaVEU8ecqq/Jn//urM264k0MvvuvuKYt/97VTq66hMlJn5JcTWeH54iy3Jswypy874E+
yY2s/6w3sTP8jz0nw5LGGZJv/13IBhwwBEdExkviHaDFT9ALGtHfCz4b4uodwRGvOnJitzkzEsFL
RubyfnagFIMkm3qy8RdYrfSdnbIom2VPvm77J9tORMbKzyILSckj/ELzdMOmotVdJgp2lf+ks7Gi
DajqcrtYHrNC6BExcRRETl5eTvicIxvVhQCfBCMBqP/I5VakqHkukjAGpx19kTxaUSCN8PP3aJpV
Rj/WvtDJrLM8X5iV1odk3dOocxcHkXTK1YOQOP6kk7TpviUBfSNo2T29AUhOBSjBjGgbwl7mOwS6
g4+goJJ95q80phL+rdkiU4gjeWOly3N3NZoIE9tBGqz7Fu4YHutVnJtBZ4OCJYebZYnNroVpQgDa
1jZRKOidXo4nimZdWotHu5Vej8/CDfx2xCYTF+nnFDro6CM=
`protect end_protected

