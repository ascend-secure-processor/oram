    parameter   LeafWidth = 32,         // in bits       
                PLBCapacity = 8192     // in bits