

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
a4nthpZCOKcSwlnR9B6aIvcbDt7FTlz4C2Gv3lkG836dWTDn/Ho90y+zGPFQRLjhFpeGZwLoot0T
Kzhco3bhqw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q6OYzyT/gdlqiVeb105Jy2yZIW4HUqSj/gQHnrG5Lh7sQmHO+iVfnWZfbtel+ZXNtO8qWS/3HaC+
trNKZWLdd4EBLfjGU5ABsgXiEwpc/RMnH5WEdD4PgYEqaO2I/kIiD3BrwovLrJYLz5j53n4tAPw7
FAXAfS1ErzOj/rp7U4w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nkBAGl28lO+TwxQ/k8h36d0GNjBwmBr+jUY4EvVjE1ykNnal5fXfD9NEGEH512COvLCvOTS3IsFl
HgVAVq2g9KXSEKIzbdpCmTGkWV0ijzgtsoga9IUc/kUZEfy5C/WiEfg+6RH6pgYWk0pV6OITE7Rz
fJDvCuPWEiy56uxmQWW0jHRlLO8/ZaJapNiOfn2gHb15pZyTgBbObpG912y1huS/Q9a3Rr3D6bXX
ZNx7FG1rUjPnyNOK/9ysm1gtTrpJ/PI0oyxOwhfzKe5VpcaZvLRj5P1cDx7fAT428WRvOONe4+Wr
JQpyZj8VXEHtuKPkbCf/CdfhK9ORwfJtnV3gNg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3Jb3rNUI5dNWwV3arF0xZcEX7KDiro77QCmkaDtoqIMF3stES6jPVixbg4FyByzgFAOye/NjCTaL
F25rXIM1erZW2B0ND6IkQmKVxfP6ISoi//lF0fgVb7IyX2KdGOGMdY6OqDW7iQltLKJ8TY64JnEp
GwsCZCn3RMjk8UX38wg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lNxjSpOKcHsvKMv+3u+x6GBJzt0oItT8as0KaSKZY5/f5wKIIjNNuehFuuTQ3Mgy67m3ZZ5NH3kH
cvgfNE2WfTFK/HOv1iWzZecvG3QR4ksXD8YNiY/ewtN3LNu11E/6X/zOeAujYErz01ZILkxEaQpn
3DyeRx1TuqR56BnTg5dFh7mhyn1xFnBqKJAVGu4PciCgJ7JVwcRy7RTkIDPh8lvwlp241QTrFinu
A+t5u9KGhJk4tbSDH9YwK23vMMbJzEwVW1bDRLrhse6ImVDBBM5XPJJIX1hmx9R9Bk3LsRhJKCri
Y8w1FqTnRgHRzUaRTjYT3dgmry9AUtI4FwwUnQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77520)
`protect data_block
r1rMZ7kgxEBp9Emm8WscC8gduI7VDEM9Q90mhrlLuMhX0uHEg+TK7oszEHy5Gox6g6PsscPlRg4j
ZTOxyubKHTFunpaB4BxiATgp/kzfXSbMhtOcGpfWhhNIrSR37zgtH9AqyMCUwCi/NIHgHQrX8Fxx
dE8qk0poAmm6jvMkY1SrpbWkWWb2XkDQAU5GxMZcOsTWw/kXqWfJ46OknTDPK/olYtmzXMmsD70o
1IHNO97gfyJ/f2ooiLvpNyM4Xq4eY7wrbhCOfnDe4cpegof9TQZ6xTdIZVk9QNaeUEsKylqCwJ4o
mRtynFSrwJhdsFsjFxsOc0PHMRzpwqrq8P7Icu410w/wfA2oXlxDq1nozRq6K7NHRKsc5kuNUmdk
RmUe5ZMpWdAjSpWUqrsrdKoz2v3ehwHDEhaLsZPoKdGkakYOv9tXPoF4GwY66F5u6P+LjqwUTT5Q
fYtTq576vrHiCQljesvg5se00CzUwaFaB2CvQyPLCYQ9kcnJ2h0qff0YMDMG9nesepJ9pBwfNu23
BH+ZOumR4s+BU/PKZCPN7g5Od6d6UVyU8mvUp2KfRj7E58YoDACtdgz48NTAUOw/r2I4+eusjEwU
h/GtAiPP6SvukHEqqKi7/Oq9ZnS5ywm43wJne/fHUJWtefCM9Addzx8q8LxfmYqsj58fDUOBFPR2
tSQi2C1hn7pKc6ztHB+/JpSD3H3MvWPhJ4nrYdJMcRFX8iEHl1OmrWeBOLrKSJ6zo/hwSNfX1hBm
73ildHH5yT7/0IIR0xD5oLXsCJO9rRgcRHzLo0gwiMx+IX67nC7e48G0WAWvo8hRjT8yzGDl6k+n
MaMgngdLoeuGmD0DLPp6uSFfsIGDXYmsg6UYqlMuLK0eJjW0U5JKfjGkqAx8qheq9TWXmLVAhkgr
yfu0yhlkk9rWCcCiwqjsDpvoz1lPElOWNWMJwMvlTz9Ab3zLCwbI8R55tl6TqwYOfKF/BhC7uqLy
glnfeiM9kkovjLuUA01Er8qYnAM35ccAdxhT3z6IKp+h0bG0FP7elVPwIBvpMxvellrHiYe8VTlQ
I+RJKf9fNuDupzp7FptXWn1oKtF6KruI1ueflYCJeSZ0lkHYIzbRaWMtOMcwzDWTBPIyV+YjchL4
r/YC3Nl3jV4pryHlTzH36qjDXJu6e90foLUGzxdctUzNM5dUjG0KLVyoKUdXaSrMuPw/l246/dnl
CnXd5MQ4Y9f2y4owycZhXMMPCB5bspQc3iietPKIPW3PwxZKoFhcHXYqTR9dOrKJiTnvhCw04Et0
yJ6SqChnIgzgPmWFhXOoCee78eCRoYPNK+KkICqFWmtQKpKlQoLBDQ6Azt8P0NvpWYl+0PDJnxmJ
d55+6/IC3V8nS44vu7mcn8vbrBBGZnxbZBR/W6cv2474PqdGIQhrb8GMAx9mZ5OPO1E5Zbpa/egd
XWjS+AoNp57p79QcQImVZ7YoMmzudoVBM6uf3QOBlK/XNr7nx1SIepzUrnoc2FOa5gZJAhPMmMPY
gJ49m84+Gg/f0BsDcGnE6UhgOys3y3Ov5VjCDuLw1mwc9j989k0wtJmsbIrOQP1ZvkJv0rtCXLas
UlVG8FZ2JSZ8a3YW2/yzyS5+bdE+UaiZ2F4BexmjqW/s7w9tvGaKOzvm+7Cel+BDzpntpi1AqGMb
qnTUaopHHR7d11mIXEy55ZYakC5yqP8vamC0MUW9IepBrZmOuC7ZXMhBIBUhh938GUeuxoBBgeAs
g8IRK4L0DaUlYjckcaUwMfsctJAp2meLptOl0MftHjfmrxiNrG5r/5wW91+vuFyb/IluxXnL1nHm
oiKLlR7CcoC4UzC1v46jdmTC19qshr9qWhaitogCDWCTkChj40VQ6QixRUI04JWyqfhdUyZRUfoi
dbdRytYi3YO9Xa/VjKWzag5TI5cQ8nk8KLRObhqczpok5G/pFJL/GQDCLn/v5DVk40QBinfMimZA
jCII+iZOWA8jNMOPJrNC6YEir6UQZEAZlT2al7OEVxHCB2k00osFYNZUQ74+/eCPWK+LaN6iWKz3
k4W+dptc4BJS6AuiVjJayF2sDtFXx0rbfoJm6B5Z3hsCQnkvOAEDwKC9PleIww+8e6EgfOM5CSZI
OpR9dPrQld6qWaJk8V6Y1tLJEh072npqMLmkmJcokSM1Z1Nca/HzrKt8bRrmKQEDIWrmU+VGkxSb
VpNaje7Ss77wKuijmBIhuw5hLJGLaCByxp1zhf/VmCelDz6chHYNJdsA456Y9pdoUm88NJq5dPYG
q0xDdV8gwYFs27UxttxlbGvLIlA7A/6aLIq1Vxm6kjYOYn3UDekRpNJ8v+dldB9A+db9qoZZN/jq
OSoAKgY+t/caXopX6+Y3jFvOiWV2aiI5GLdhZcG920UsUM6SsjJldNazaP+aJ5yHneYeCKXVJQb/
d/mZPaYopstDdZtBPAZQ7Z3Bw5VCMAg2uWxW1PfSyBoUMZHETxxeGJpZVfeQQQn46maqtQOgXeXw
IEQQcKio0GOaaJ83kbr0HTo/CnUwYFjkV8G8PgdrMcNcWGdq+7x3YZhKb4tRTMMVPLskO8by+CZV
oWsibwCWZy7o/ucSiFwbpZbYCrH3yDARaW8nep8o3FQRGZ6P0zZApyC1WgskEC1Zmaq56Ruq6iWT
yLUShwrfvWd5RTEjpzZX26vIb+/PZNHG5aVi6qr+GcSlQhVar2whoXxRW2ZXSOq3UmIoOHvBIiAi
mQjJ15006YagMOkZkT8SFDj16hD4y2aklQoDXDVlsid9WwGeaMgk+LAZHf3uDnS6yVq0M1wfmGbZ
vvW+Tz87503Tq57xolYZDZVJqwI82X3rzjcn6NRZf91PgbafJF1uNBfzGL01jWBti8B0KnuoktBp
jblGuai6Sg9E8H+5NxIGZy7YcY9Ro9rp7acZ7QKmyFjXH7c5FFT2EcDydqf87vCdTTGEfD35YtEv
gL33AtfM6c9VXQ9+ml5XvvejuNGbql9/p1s/JIXvcbZrCGohUoRWEX3f7hfWx6ZvXXfFOSJgkcbY
KNYW6ucwtJ+GbBv6/HNgj1U6jFAvocB2Z+C17Y6nUImfmkmGNtuo4glKPadPHLaDqTNBb1dH9MOE
2EriYhHcVczEgoOc7UcIyDc06CllRxe2mMOQWFc6NEcWlFCzKexpzQjTDsZrRAk7yTDJb7EHJ4Cy
xMQYt6TsPOryOWT99O89cXV/Qi97z0e45z7WBd0d0E5vqJFseV5fiWE0o+q7fHdpZdA+pOYv5XsM
GUmbaQma1koZfW9/4AIZa2MKjdddRcJXokv8H5rsxqbD1t579nYldzI27EH7ldDgprB9BNT8xW/q
tvQ1EeVHrGOzvFwFoVPQ/9fZGzqaJmv1gqZL/1ksonh/RJ8QOBTMItRHX8Fhf3nc4xI9MiM4ZGPW
Mj62yMR/etsOWOnLeL/ERDWC1Q8mdHTaVfHzAljiVl+tfb1qR2wg/qjogwJuI3JgH1RBOQ7pJZix
PMRreSK0Bok5Qx2ufLay4tFPC7L115hdBUWp8Tvlu4/gHdW2DqZ75vstrhDefwzWtiD36kaS+itX
Vdo4j7hru0TdLVQn2nHqyIFts69NgyEGZPnx5OCCUFN0tMRxj2D/C7Akv5nn32ieQAyQi+Dc4Mad
cIFwhfN3MtXu5t5Z7Hy4TnQfjuTSSsGcGiCAYxxmW19AHAVjVmHV9XE+ELlXhQ8ofTk5McFkTghQ
Qh2LSoCB8vMFKssIpzebVvYM4YvdMOz/ve+SgVrF4yoPpj+2WnVY5BxzcSz8ktbGQaFSudcBXjUb
ikVcfdG6EcBBONToReJRYS9HDQGHDYLGos/Ea8KJltDqfv3ew4nPuk4npHW2tQa4boP3RDivtV+P
TRdjrf7V3aeeW4AOTw1jRc0gUtuaEJy4D+nIvit/koLiLhCy5oleRJq0Z8Wc2YRRjbbYEwXVsSGP
dWzSQiG0oFoZUTo3g7thbKEinjVol4g5QmfKJv2vK71k9Q3CLiGYTaUVoKT9a9XammKa9KoqoB8d
LxImJqKzQKuYSKebdJP6xCdyLYIH65eSPKtVY1es2Kf9CZ2I6G9hn6Zj1wxHP6Iv2SxkAfVWtfLV
JXDTkVz4gEBLJlep21LNFHxyXnE0v8oU9rsj7CuKj0W4JEwFTdkvQVHljSQLs8BpicVhdtwXCsgD
rIlkmw7Ffan3VPjJj1HLDzrVZUN3HHY6tBstn0fg9IYb2KtkEDdRyJgcB4F2X4nbEPfin4EpxBp+
Gx5/L+EBgsMEqiQnSGPtiUMGSnu0w4cjC8Qq3yHqA/jKAqi4muyAY7F9vMx938MPhV/sV6rDVWsv
/zlg9AF+PLCqvfnDTxTVKrA6ZDahG7AiEyqy1J+PvmP0K9dBRmV2O/Ht895+YRHxiX1fNm6XjqCY
zjGRnMQNX0QEaTJeqEvZo3EiLLByOCLDUOFesuFUq8H9gGYcG1XF3bWU1GTO8cuR5zpzR28PBG3m
CD/FpHmlH0Z8BL4zBS4hLdCQ1JOpNrLd9PSPJ5s8+wKsf9cQnw31FlibJVMmXa2Sc09qXtnn6Ehq
5XUrZdTb87UonZT+3N8PyAUGb2rKq+Ub/0fSyJqvdxAmTVQLMileIJnQm/yMKyXGrMtdvAaLAXdn
5vklD6ZQqZjsNd9mcZaE06RtWGoaUFX5mE8KMZN02oMSWngDAkbRgLRNgMp9B01925t48lg+rXyW
NOjy+LHOQLPr+xCTFQeNe/UBkkr9nS1Y1ADe8ph21BKopJdzeqCmPY61/s0XAEEjI/UY7juiLIFD
TmiTYU8e9YI0lWuvJtKIcrP5h8Ba8N7kgv5/4ps+OFMvD/RAZpCSapBwvGKl8OnsAJWD9H+DXSPF
X7/uzAjRkbj1dWJ0ZlSprKt7rNjZ8dfyQMKIKrUyD8Zni6j9KJMdgf9FhZyMHbfJner0OjDG1RzB
3JgbQ/3zsw6R1T0TecFDNlQxXf6pjy0H6337YbEPbRqwas7bWyyQ3YePr3e1qOa7ng190xEvRDQJ
/wplAaOBLjCmCuF7AJ8/4pyVqUQiU4XLP2vXYeGupLNy1GbOuvi5D1mG1u3e5pvkWY5fP7xc30e+
ecvMbwUPcyks2ZHcUuqT9fELhcCTDCRNd1ncpbtEHE/TC9OAVOa4ATAot2vO8GZZNnt9126rtgbe
DNGFo/7rLyYMedwCDqEXqJw1nWDMgz1S6+PbBDI2LubbBkL9QrCblK13NpzmrMniqWmjQXhEf6iW
iD5HOyvN6UjcJc9cRI/nX662/J4ypDv/FsaDbIrOWh90qYWH9N7fV2nbHUd8fsUG8cQKZ2g83g7c
+SYaDRXR+83DjfG2GHH+ziwC0dVRljMcySSTGm6G7lXy97hytFDtwaAcyBwWLqrCqRqWdv5HAvVY
tgcXUTM0ut2hB97bEPO44nQl2GljVyin7AT/JcVKXu9eKp3Sb83U40XYl3jenPwNXNa3I0MFwnjA
rycAQMLkKsxSwYUKyrF/NnZmgdYlfLsRpivQ5MdUbfsFg/NI/NyaNmmtiMPM34qka9ENMrIww0bB
EORbCiA1Qgr0zZ1/bhu2K46awpRqEuKpbLBS34MDITzfqT32b9otTcMBEBYU5wrQ2/cmbkWihy7e
xZNZtHdGxUyy/5ST0bpXWv9LKHKTWT1BkDosjbLZJ6TU7B4MiFyWaoCgAhzxv27T6ZLV9gG5mLsg
FrV6n7pAdrNnh7O0pAy9N+stzM5o3Thwq2LqfrEuILf1evoztrhppEeQ6pdWB0yB+jJKdvRvHFEk
J3PfSIBZBgb3dI6W4YIq0G32nF5Qlskw/j6pf0c2260rtHIfMGnpZHg+xINJoHwpUEiIcUeg0YPY
gjNj96v8v0ZEX8eek2vJ8mI1qKrqkT31Wqhqxrfvn/cUpGXVSExI4Gn/jRk5ACGCSP25Tr/e1M6n
cuRYiXOXLRoLE1FrhPXPWEDJ6A7kpDe78FqM40tIAUndd60khbTeXobDsjoYljxWo5eWZgbmKW5h
8Zc81uZFdNnhNdKSW2pbDHXkBk9MjCvC5Ln2fGT02wVEtin81rLhOAsU5ASckEi2vOyx3GvDNcGO
Ks4psiZxfJI3aBmobKQtTGvPVJqTTDKoYy1I6vv+NdSVjATKDZ6r3eltN+cK7Cur1YxlNxuDiaSQ
mQ2RNnzNK6zknciof/pNpBKodrRhXSakmqUcURylvGSVvxZfX15BbzM+8IHmtjo4F54s8zijQLCZ
gt7kBEPhZ0JCGBePoOTa1bIhlIuyES0DGhxadRFqLU9EOoONL1BLBxTmvTlNzp1dV8ybnyfBqTBL
gSC52+vQcz2j32qeTQ6VwctBNfcsZDtJoWbJVGdrdFm+4ur+FvVuaAp4gqkMGkxVCCchyJtn9Oe7
M+QHjk3T5NIACOD1NbhNgzcIFAtEiKID/FAkIt8obFQ5IeWiI4oca0kAkYC4nNMqpeHAibE/n6si
EtLfXMOeDFVWHiT+a/MBVp/SENW8B+3DQXwjZj1ZyrmWhxJ2J6XcgtyVw+JZgBGb1y0p0/hjVnwV
vsgdyP6Tqy9nKhacC8dIdEaAgKuFV8Y1++K/SCfK4HiNYkYxEelOZ+s8GWTgRAQSqbldIFr2oHf7
xOvjJRZ6AmNnJABezyS2tGiQzCPACWCVsjYBTmTKqN10dlMM49y8HPYyB1XTDYGzD+c3Lr2sqEFf
z9PZnFlPayB0Wc93+Qwf7tw+SSLt3tc3YBrNaUVRj+KGA+Iocvf8useMcJF18Z+1WmxRMF04dlcC
Svk29ZZ+GE5uKMgk/aJlJ8fcPcwOpnb/PKBlirmOLFmmK4oi1MjrEzkSieAqj5UdicfzDrtWHQJY
zdplfkHIAB1qYNn5ses3TPvv4hwl+lM7V1OFUYE42gmBU/hKx3N5w063YAsw2TeguPMT69SbTSt4
UDHVcoz1GbCpf1O1ORVXf+rY/aXbCXqsBjKLW2rt8gO8LK46UQeSWOfIJUQO97CHmmKJaGnoImQT
731udtI/iVXhhylirclOESc1LNUBzvyUf6EPKwl+dseoVo+bIqQKj0P76aAclJJfTPfAD9HejUCe
p1YVif7+3ovqeg9Fblzk2iMQk5mCcX2wQllWMKgFMv3ChQnsmGAXuU2GHgWriv9UdKMrkFf4xcsI
9Vf+k+h1H+PaOUmhe3fHaKslPNC870wb4kOBLU0aM1P8AFmnsLjfBNisZZIyuykIW6mMvt18FpWY
sVniikhIStHzR/X+0Tz8Ez4mht6ZZcsjuZDRtFJjFriDo42AjCO1KSP7jairmlkdQPAKj37YBQoo
TuNZUW2rrSJV+WHXHrfNn4dPhOtO624s1aWZEkQbDb+wUMWAzgYiuouMrZmcJ5pP8QMshUIFJ4a4
7YhnzFOULDdAewqlQT9uEKZOl08RiKFHuH4PBMhf12R77FzyUdPJhQTXismmqwGAp4ncIVJQ8Q6V
UacCHX1xMHMx1sdCy8Cw0gGl4VtTDc5GLBGKuQzn6fIuG7RsEm4gYIGNOZDxrQfEd/ojc6B8K0sQ
T73uaNodn9aXqHMkftcq2jth4BnQ7Tz32waSEXLwHCB5bo4c+aMxX6NG04kccFm9dj/77jCkMYRK
h5zb3L/WU50M6osHN5g/V6mpQtorpwCVQ0CLsUkbMemAbAprPRbLco+d3O5LTmJ63XOeT+mFFDCU
a3doRKew+9TD/X9B4WhBJn3nYWfwtRPG7eXKpycBbN/G1FW0u6e+AQiOldr7lemcK6Ir7BREHD9L
cf+P3PHmmmR0iOCSfubXXTDhYNfVhH05j152s2A3ckYEwCpgobel9/V9r4bgto18MdUDPYPLlsif
SoPU6epwOwSTGUbLx2Tp4Je/P6kqdLvLm+iSCoIp9j6mehdu7W9UVylGLIo/Ys1wwwweBFb4e9Vs
4n41EnvRfexS/4POt0uZ8gvY21tGHUyzSNJvrQluHjiGXqitLGj4f7yfxm9IUqZ/q2NsNbkCavU0
k8kKrB0JJm2ffGXMi9NcV8zU1yo1Dhw+Go1o45hh0ke7huq0+pp7Vwd7nCfprJYCdEPRlv/daRlL
LCYTFs0RLVYQGmtV6/VU3rBEQtPo+5ZBZWCZe2sTotVDUtQLyKwXVV9XQMR3jrkMr0K4hn1IGpzD
ZrDXZVOIKleyVyqhxV58DR1NFdbLesbzb4pH3LxsW7EROAtBekew/HU6Jo6yoPEGcAsf25IuHIso
m2/PXkruPuOaTV4SaxT47gB62wZ/8L73nJnJM6xuL2rRBLePGvQ+xjhs3w6XhZmVV48vZFLnBK86
1WB83cGVfm/4YyJ9cMVb5k+n+AKVBfGSDQAKYoTGKrsMVLCrI7Um48vcytLMG9kb7/OeZ2ieRz+U
imNwQtMzxJuj38GIWyNi0ff2Tug94oKqhE3SG5xGjU8u1URWXDYz1Hps/OoEmhyROorBktOn2YtF
9qYSbKwRNTf5mowoaervB2shh4ECCBEgAvpqYlkxc1nCV/YoBG1HkmKY5Gl/uGvfotjukrHqYWee
Al1/3TjgVlhIMTna06E1fUS08c3U66RNDwM9ix+URwdsVnh4IAzM7CATu9Zfh/i3a/xrklNfgiX7
aeH1Y0twzG+EYQTseEnYIxjnSFNtahudM39I0E1j5ULt+KZDB/JjUHMg8xsH4KCW4drS3SYeSbW+
40RfGeFs5m/0UC1/2/LtJkgsr3AU2H5ajUOo5qDFZLu2jITb/IWBW7Z2m/C//UA7quttgAORJS/g
53r+o5UUSGptvkRLY+noR/4VTjwilqhsKbN0UE6fuS78LvWoBwK0Pd8qeekg5NG7jkBYseSF0eSA
NgEcKtpEuxAMRY90mBNF8lexic/zgHYjjdzCenXc5Jk7bx+w6+uwY0li0bat0313kKbpSggcrLhI
SaruTvpsSelU5RxpsWDbXNnb9zNsfPszuGkbYldzKmH0tV3AbldP672U87jDZbe9wgKEqcYDFUEf
XSlFXYDbBbU0JkWOOLo34tFUPhd31/PtoGYP5bH2JVOG7CUsDRABUJzU+9ccsrZqFDeGm/mUOtC2
O7NN0/Hvy4Ukm/8X+391qRoNIZb59kyZAghyZTuc4cguO/SZRT2dAoyj2h4QN3mntlwCko9szFUz
RXkcLCgOuzltVtSb5vCz7zAcrOvkSLyeZcxdUnm7l93QPliRBZ3boEgWyJy69Cs0+dNPIKKoZdqk
D7o5h2ja4PSg7Asa+pv1gFa6zdCafjE3ZFGqOprMSqjuHq0YfaPSERRT3Ah1lE4uhM66bHlzm+vx
HAYg8lyTvkAH1KRJ8R5BXePcC0RdCG9a3B8myf+yqHQf6iHX2CDvYFnkBK1HFZZP0uH5knIJOE3G
+SfC7AvGPIQY5IIEPbJjZnq84VI6TKybb0kB3Fnbkdr5issX8lJC+eyW9zwyxABSmpYG+45fpAVy
lnV+nxuz9skn0lhcQmcza4U3x2jaDCeRHEmVpI93bjsugB5R+fVx61OnCPfttJb8tQNuD+ebcfK7
aubTGUq1XqcztdfyzqHBQi2GbBO7lURSji5eMNTQnnFBImUwq5PQy3XIq5A/TVF8Ldaf3FwyQLma
yrwH4RFpXX9eJT2J5s+5z9KQfWczelHhHz/RhuJdHvztWJsoZ8Rd20dfVDEnkNu5UyYH48hTgUK9
wVNL1qxAsdBGYCGLa7EA163azfbNP0Y0S7rru8kzaoUOYRCM3EqJCkAHDitIJe95Tp9RVdZKPcHd
Zu67BpZrsYjhxwmgWcK56sV7TDJ0m78cpXjKOAtbrOSpw1L8AIGBLIWF8rS3GdX1sUD4m3ei+EJn
mG528YHlS5J+DUYJ6w1z2ez0ccgI1/4XBWOQabkzi6LTfnfGhdZEetw5KaJIRXD6g3xNxUOqqXcI
qwGOVqcCayfghFuXMmU3W2bMETHv6m+A1DAfR/C99WgI12ZWqNfCWpbXCDwWnTvRyjAu9+a2Aj72
eLIjBw2U8gj0gN1Zd3V7iJS5HG1EBwAOMkYvZiaCRzsPMen98IFev5/k8fdV+Nsp7hIqX1bR08i+
vs8o0IkP6UQB9Bzy6Fq/K8KDOOVRDVFA4AbV9kPXjRUs1DU26v2MV4UY5Id591xvThkgLQkqi5tz
dXaO3ro8m9nehNS79m4xU76KZmKJVPylwudC/AZFo7niTX/W5JIo2uPXkfvdqsQ6HIWpOHaOqCsC
0SKK2HQ0XMQL4ChcP7XeCQ/a4EyXzo6mnI+Z5eyMeymy1Z4AB+GfX1jFcpY4+BoXqxZCLHYOJBsn
ZxCP5FMBUHZagReQJUnWhee5lOes3CLlK6uAhI2gTuZ/zNlrne0CuToGCj35OViEJYGbbZH2rC22
Ts6FDsPfjGbbJkJlsvY4TOpFWV3/1b1R6wZPlvSSO6bXjwPO0UhFJd6S5RrTDhPm7Wek/3xZCRcd
ai9pDD1tJZM8EZb391rGKi1A2NXfSGOipDc1jHoKYqRHmbEuUKmrzF99+59Speu6q2I3uijFSwYb
M0r2Yldri/M0VnrAQlB+xXV9RwK57u24YfoY170dXfphmB1zjq0KmLngi1xfHQtCudBPJ3QHaoaq
BmlUzcdknW+zeGg2YOeOW37jQoa3CZgPUOnE9iTLjkFxE7xRlvx/34g5C4CFeP9FqRnFGEL1Bb64
5jPXYyBGqhvai4IZ8AnstQ9adVpdlxmS73XgynZp9wi6wzMJMulKu0MEN2MMJOFnk6XV4QHvKOL6
O+UWGp1XS3ygV0rwQpduye6XKzfT1zCmyoNp/wl2I9hEKKunhvmxETVGJu+InacbNB5FWKc5mFqf
8JzRIr3yHZQqATr8DrRfLKdKKBXwbYsRfcTj/Yl+MX5psJVHQDoGQigaHoeBRg0WFCj73Ml8MPVk
8dD8j4mBauHwd5a+OcH/0cRaNYFaB3imMAn22jT6HGl/D7w8Fk7R8yuEg0pDvPGRCijoYhI6/8ef
Sesjt7HI3+JeHcFkVsLPs2SOgh9DtQLTO2+Cu1GHzIgSl/cOw7FDQLvylKmFPdO6O6MlmbsFtFlY
QaOqUm5o6ldr83IgQ7YPz3gOJjOoVN1wN/0ND9kqXEaPzrrSoxMxJF+D5AuDI9hV0cILNYQ3Vpgy
+EZbxBzz+tdlRqyaoCx8NaSdqjC64ZNCXIV5PLlUwnCNkAaKP0tMxVmHKXYSyhjEzjNTzKAtpTrO
kPWKhdJ29abJmzmOw77cTPJn2h6n1CEAdk96+CRqFpMV0hgpLpX6zkdSse0jhfMfHDp2jGD6NKi/
6s/ET5OTwh6rlQSGLdt+WXGNgzpgmqzZ5aKBdFPu3Tt/JAmZHOfcFSXv05IIwVu3QCL91h81P3s0
QMjOr5F90X0mpcRv6hQp5sC5Wq3+jcnuZtkxvK7bLJrwPs1Hs9G+XvuvmepckVmK6s70NxZe6tJq
+CWZmBauvH63Dd9ZZtN0PtFgmw1pIwXPCK6yTm4mTBRWvCA2acQXCdfNk9FLkFbln6pK+raABqzL
sOzpp1ROyhRDaprYpIlndVrRlelLEHft4DVR9rKMQ4QDXYBEVuBlslDpwqqXpKFFn5DMAMLNB1w6
PLQQZ4Jr3rjpgTSd8Fxx04b/HUDOELPJyvbIBJlDnwSZwq2x1G7X7jHpaekvq+YSnjBbxgxUUqVm
UXgJjbyLhHEziBYe1FMo99tsJQN0A8GwIliu7/olRa6lcpwZSPD5x1zRQ3nvDP+2aDCvsa+Lh+7Y
z4uH6Ryame6O75D+qhvkdNDRZukBrMHI8v0ZaxRf7peXpMiI6ZBG1mfbTTOyePtTUp6Pe3bxP7gz
zfli+rytOt297zU0yToQdpDjXIU2YCXNUoAJcUqkz5R1nZXv9WCQygwVdtUGnxKt4TBzzoQDeN5k
yRSAS1Kw6/53zYAQDxM0FjNCvyWn2oq238airfB4kvNyo0q5q+LbvL8xC/LHFrmbDp2aINwn8gky
MKSM/lc+j/26TbB8JInbUW6dgsThXfvXUe9yjB878AoawgQnXBeqrJ1/FpMbCX4l3FatiTbYNwAH
oQal7X2iZ+Z5pjJAP+H2hR/kYmM8A65660pl42mOrumsEc805tW+SCUyQ7k3CegS9DOjE9vQl3kG
JvXJ94r0nF0l1x7op+ZbQCJOloouPi0mkNPrbiJhhpFx1zjqMX29L+YMyLb9dCdXdIij4TdmYrXU
8Dyqzl3Yao+neC+ilMXrjKINvD9e66ZwbPS5XidEEud7RME9dOG6peIk/UNuxos4fV9RCbkBDKy/
gnlVwErmnYhz51V9XGZnP07OUcmxQ+eIqCjr8yvrXbe+E6pdkz1Cv4t+3Flj5d2JaepJQib+58O3
5P+f7oDoYBMRonTweaphHebQn/TDjOWhMAlqwnXptn8KtHk0hg4NtAeKJYyl8s3e6097/5FY3WH+
auBavXXUwROPYzNkvW9e5F7Dk/oDK2UkSJ3PdVZULrndPrEoFovC6bVMcruLqmJGQim1toIFa1OQ
YGTzVEWIos4sWRwGfmkYijDDhAOM4oI0mdHBWr7Oaey2u6lftWUhphQ4zJEnd4+r3Eo3xKWKZskx
XHBl2hLb0T2CX6GiY/V9Zp4hpKThwOMZCrsZ93K7VPuWNUAJ9MakWvCatLtovWAOwWXbHOwg/K9n
cElHBK82uBMzhV1nTJAuFAxgtxE7Ci6bwNlWhggBJvVZGHwwWa02GUu4mhT8tlvyCYJwhfsMvjoo
zRF/SbCmp/Z69YIMfzqQh85kMSz9F0qHTxo+xE8IV0Gt50dw//Ru8+jBOfz2PnuJ0xE1j5tur/21
a6nDMvzDQefwYM7lh9plDCDj9a8LVkxZ/mRNaU+x2t4x10mOJ+8pxHQZeZc3LG1Uj5AGckz3Ab4S
qoTl7mK/VVqdhPoIGXacJdKejClyhNrOSDNTB89w1NgvZVkKuCnX2GZJkR9otXqd4CS+6VeN17Tr
he2U3EX3QavUKM0IuNADfGPtAixA6bOedKZTsVibKmDQ2BYN9pted/Z+dM7wc17wNDxpp/WkhWVe
OL76pBRbpZe9F9OUJVmebxnTJ1bKMOXMBHw2Cs/q3xV4rEOyVIpHylKLNG8gS7jFRxtpfy8r0WZW
hym+O93URnh+lNeLA+CgwaWgdH5Hts8/zHP2zogY3iUpsVcFWvywN0Pf+J+jhh+gBXs+XXSgl0D7
RqUR3rIv/LF84lBUwyF3eL2anlGf2SwL70d8Ho4XfEIb0XVML35BiPZQkAak7YnTa3JiVsz2ahmK
afQv9xHO9ryQlGbSLnng3vxxNe8nNXOPqSzDYHF1twuXDuhX+1Bb2uBzw8rQdaOzM26Si9YdnxL0
YOSdkDgrig17pXCEUjYuItydmd5PqnlFrNxLGa7Ub9wOglBJZFODcxx8JlMy8gJ5xEuVLQD2ROdc
FRfkwlr3G4g1r46NzsAacSFRJyieei9OcAbgBB8XArBY/4LKmJ9373XvoBj10rmw8Ls8JH9jDAEP
MR8GOulv8MCo74cKZ/sQeobv32JzBeOF4/MZ+PLhUqK9kwodqjUiAQDvba303jsDcA3taEB60tNV
MfeW5wI3PKKO87i6OEad1ZBc+2EDRR1xpxbZTiR5eeWuc/q+RINVZG/23wjyX+7b//z3GjMcSgZm
/H3M1glaNL7j8dxNXCsN6dKpIZS4T8EMMuckoltx8o3lc9o9G24xBY8nhGr2mjkzPWR/ywSRgGZV
VGrMajykFemdsxY67t9sG/D7Wdx9iXyzv85zM7xF0OJnPpbWkFS9lG7ZXrdFdb+iJPy4fJn0aE5c
4yxeh9IhAmBSpcRgW2mD4/HrxChzWrvZSjywJh98xBAxGpAPvINJitTK5RbFNhi34QKaD1/P8TTl
Nbq5x1tH/cEbSiRz8r0vJu19tI4XqVBzPwDbmBb/oIsNyaUo1oL2wQHeig7A0GitfwsCr247sor6
ohvFtGdna231sGRHaiovQ8QnORp9hch21+jwYM+vI57jmNLPI6qTULvrYOhkLBtydrtMQjZyPe9t
I+6eWspJfpo/PHODiVAxkILp0CPtWhQYd1bJxwPuY4wkdDxnzrzlQ4FMNkiDXWco4Njqj4/69B2/
ASS6jeg3gJxv/Jv/pk0C0Cz14fngaadLEq/sTCqSDMFFp+PX7oHhuNmJEs3t6om4/ZrSm3JQO9dO
Ur3Q9P44pbsTN0j/kjbruNnBRB1C+qnfApR8u4wFYA1WOv9xNgf8zLuAubCwTVhANiXMYaG91s83
efvdLsZmBR4IGjKxbSELTDjMq62rwzmxQy8vIHoXzMkJP7/ZqoiDuSzPKVFzPWaLfVfd28Dulfg5
XWaa/coMKFyEh302e7bn0Hjp+6hWZcNPwkozpI36sCSGUHj7C8hnv1cD1l4EYQy+lFJMNd+3FfcE
RbCQavXl/V3hRiIqsr0wvs7O7QS4g4ePfjqT464ik+/hw83xyGvG0qX5CaKQErsPtdaBLiWY0QeF
JYJYTuIigm05j0Oalg13cN34E2UHcF3tZUKlzC9M6TZCrbynPdbU98C3miO/rSbqntfBHQWy2qtb
OSO7jwVsVTFSR1stAK5A0uEMpf8XMcrVMhtSHIzwgyRjZtv81s79ARX9icew4nFIf4qFwPZZRp2R
fvw9bIL90SY3vr6aA/JIAnWtyPTz/6e3192nNn2aioNFDYTQTT43jsU1UxTNIPn/jHKLzPTAIvSP
PBk96cJylqRyYBiLd8NpJJCCcotPRzuQIH6R64zfbGibz66OVTKfzI4Ikr37AzfdxLxu647rT3G1
V516LxFpZsgEh3UtJuSfzYEHd1MyKmp4VcF+EMWqgrU/or+zCB1dgXciNBzhxw/o93S9aNvKMN9O
fx52EW9mA6mOc/uZyTEXqHNY+cT9mQZ+1Wooc1Xxyrjhd6+0PVJVvng7OsFRqZE9Mn2eC5YPoEbi
CQ7Gexr+1RqgIY/OxqwTJEYlYu0ASvSf4QMezRRzzU086eDMfhwQon6tRoHIeb/AgzJJaI0nv0k+
6ZNcIdfQQhtuyYQCsxfa/8h2YW6vCqR2tngP3k5/5gWrl7m5VcnKUZ0QsW6Uii3f4JgiS7zxoVyB
uDDSwc82VaimZ8C7HRrLxiUzSKbDOrpyOuIHEDun8DjneoHrIbwUGZsqo9rRRQqa1dFhMUZCwr7c
j3Uu28YuAATZrD+G1IG3KZwcT7wLl9c2NLiwZ1rODb1XINS9XkGYPvn9qw7RsbPd52ox56D0wU5w
fr4cHua62ogu4KfSckF5wQHPhHaUlJnVl+qw85pqvvdH+U7ADvt2Cdl+Xvw+Qzu/LPMgY+kupchN
jDVW0n0AdCExhedQ8jQ/sj85gP9ij56eUfNW4fVn8a6V5KyMj6XXT7+XMh11QnwSLV3WH1Slir85
85nX4PnapxcC09z7ux9o88hhzkUpn77YvzGSnwHt6+Jk9prqqHTsRR52uc9tB+meh8+T8aygPkiO
7OTria7c0tF0oDx0G2NzKxB5N1DzvL9VtLeftqmSZukhAKdVclwDn91pG+ETvh5j48xmYGwzOhCF
A8Yg/Er1LTRF+oshSgwRCI7AXv6oQmN7fx2q3dFFE7Q8pZ0MghE7jS2PfWTITIhffMt7U7QeV6zb
09/5y4k7BkJgSm5HKLaO62yTUDsU+SIAQ+3vE3Y+JYpGHA5tfs5BeTJKw8GSQpAeVvcS732VI0lO
R2IaVHg6DYfTQPWUXInt7cApluviq7u3ovNRpH0HO8mBi4X+KSprCvo4ttP/jWyUz2sqo6a4SNFX
CY9NuoxItU6I1NsWH8gp40HPRi8FJwXYTXLdMaX9Rc7GIfSO1cetfGjJi6Vdps8F0LdoBI9+29E4
BhP6GnVnJW9J0XEPbz7bULFCfH8bZhZFtGg+exK4YX4+NawopqsOVhFN5Ybtg91OghSMbMuyF5PQ
iVEEJTber455o6NOtBxMf6eyAt9AIJoFYgIAZ6hk2R9WbFALb/w3O98R7OWnk7q8RPAZEeLDLHJ7
6x5izCBwETBjFMrjMCC2CLiEWL2OLJZH8MaCIQmP+OJEUV8QEVXN4dmYAOAc5ikM4Lj+GlzrvEUE
Xjgbc1Sox++O3Utfs7cwUl+TrqHerTKQehMFyOarhRKey2WRtyzfLVV5yXMh+o/53UPbD+GZww0C
4bmfaagyNehAjgiR7WE2UrmnDl+7XAc2+E+Lvvbg0enQDMpJwi9QhDJk9RsPebOeTIXD2uXPlm77
m0eICzLBIBgO6HkD+nGhgTRhFXlrGewQ4VgVjKy6hntZJ7ZNFFDoHmGL5L1pePnXm7m92jEFbLJ3
/gwHyX1ilEi4PimvRF2aEefeYD5scU+NqL99EtcqrbKUeUinkPJG8U0UQ5Fb7nnpDYk7uscBLDdP
/46gbpw6FuvIFxlmfP2CepFAdRIRydlyXPrA+Wp+dADScsKqfv9B774MH6dAXBbq+QZ9qK04DAuu
efzQ0JwBrmdST7ki5LdgBkdNqOUE+hrFiroEL5747wXVVePU2j3DAEMsku4H4hv9ZOUXCqKYi7L9
sDv0nLTaAXmkUX9DoNabxkY25ak6ivwGRD9abpz1PKHvVA/oMROu6pP+RPtFQR33h4Zi2cWaUpWd
CZLu1Dyl837y1KabGRC8tjUqvgDChwQsQMR4zbSasDsyIgnpiNOEg7MrZu/p7ZcLLnt0PGJ1BzdE
7RQXxWplGcAmFcMxtkHb8y6grMyn2S+S8awu5CO7Q1x7gAibHTgx1mclWPKtLcuSxjY3aRuCGrpz
icakJMkVufhI/2kx792MSfZGsomsdvThSACa55rAloNwk+c9pndPoEf9q9he9pVHlppV62BUwbcv
Xk7e3T+tjRiaMVhiiGKqiUvxXRnA5q1bB0z1R0u06ACW89q3dHyXzSszzb/RsMpcyqMuVNSHP1VR
Nzl+2vkP055uL+u7eC4D7irR7pXfAt/uuoUhdNb+zXyJexdNivqdA+NDd9ogDn7zcx/ozNuuzHqw
uKVHuZrZgJOQNR2GC55aR7BcvWfTP72nI3byBdnctgZKcQtJxfmCBw3kmd8xG6PrRElbY94ZwcfO
O5XKVmtY3FFYzQ/pLVJtI8BukZnG0V6wwPHAzkaEyUs7B1PtcilsASgmhKqvaSxsMMNZ2vtxSsd0
LMvFoSbokiUwWbGnTnBYJuT47CQnrGcVJgZL8G4LFrjP8vqB2CLQrpTy+TwsnMkqklqJOJzr6zum
sLeWwntJBFOkN08tYZOP+/goDQGSZR4my09JzGQqhF3oI8OCmlv/bCtrMPOqHF6mQgqdH3XG5fSU
QT4S8uoGxu7ElS7wi+vTM52Zs0FNiizwvh+2dmUlJNJRwfmHp5CCxLnlD0v+XwnzR/B//LJUDIvn
CE4gNDXChTtDHJRTBs9qFLFz4de8YkPSYw2hvaj1kS4BYkemZbJEt46wdveKiLigC89IStp/Nw5X
J/8ID583e7N+RrPrlQfCyrtGd7HUfQ66/FwOeghGPphysmIAparYM6CXS8h+2n5wqfOYpaDWOLZi
J/5foTGkEfGA0tHb65KyOYjuRDWDFmNGbIYP7wl6qSJkBwC5BdVovJFI5y/ab6tWTKaJm1wG8LIp
i8gkeF6N1sm9T0FKR1Hoc0zojHqAFVySo5AjluLfHanNg3Nw+n/u7a+ViB6GPGRkyzJUYJUydz5B
bMmwr8a+yZdcEDJm0IOLIC7zErfUyVkkSFqVSkXNNlREVc+aLE3szNA2WsGHFYDTSlMHOf85wYG1
O8W0nzlY+GONdj7PosB9Ncvc+v8HEpyG0l5w6skBkE81o/O0cJvrNC/UzoTqGl+V6pfQaGo5MDaB
s0AThjXe0Nzd6o41+DDroWuncgJIHgO4lpB9REM0HR2G8SUN5qzAVYKSANzXACH/Ina6ICNO1ESB
HDGAcGv6+o94Ge0tDa0fSFwVsWJ4yfKOWTy7P9fyhwk6Xj0tV5Re5bPDs+9QdD3kEhgtPKArNXqc
2bd0JweNDUCkvzdyO02FQb7UDz7RxHudu4jaOfhNBHIZ1ms38fOWDOY8Hy4y6WASJ4oIZuci2ss5
aMtLRG0eTih6MzIqtKpUZ1SrlFXVV8wO4TPgg+87MFzXcL5uBFioTS0wuBA+osFWtBAzy3S8or4E
pyqWtxOplcU6eUDB6OwXTuU8W7tQEUjgmrj+XipPpBp3bjbj5TRFSAMRaAHzS168YjnIpDiTor/w
dFi4DWG5tWgMQMMhtyv/nP+JUrgqgluX8WMm0eVkYw+UWB4n5Xan8VlVUfM4mZqcepmybT+h6y9w
Wmwg9rzuE6sxUDssnj44NwaH73MKFVeTi46XzbMa0rlKfFoOli8+VwNjU7etzKt0ckOU5cux6BpJ
wWCTxL73Z11qQBtS4PU5PrnNuj9a9QfaG6QSnygm785+gisXjTM+sYs7u5SKB1GLCzNrd+9vAoFR
BHFlq47rRB4MMpTm8HvZGrbWr81EuV0QwkkKtKWYF7d5+JsR7LVS1CJ6Uu3Ta/iFVlBspK30Oxeo
gkrk5vXjBQFmae3+khlxcMxBIrgqQ7lhrFMTbmDqXp6XQVT9PKOZ/oR/zDWirg+YI39J5eNM6Um4
6Ef2wiRE3ADeuxBXrXHCOHCTkeP8BKFo4yxyy2OShh5V5Ku8e56VhCPnLa66G2dsTl8yWuT0xACf
p7wA3J5Ztn4ZHALicp1IihU+8+AGboMHutIHPLRFjTAgtzf7+N1/I4+oHvvL+MYTNI7TMJubeW7R
ll/Cj1Jnlr5Vx/zCd5+On7Gmdh+drZdWFDzEGZN7MqxF97gpmMPvNAowUrKiIMe66V9mJ/O4nLPy
2uoZyRgC0SGqIifVaPuRY/WBiLUZ0I14eFgwj28SQw4x1eIJv9TfXc7R05RMthGuirU1H1x9ta0I
QFnmsCWNimaF/4VZRr+p7ALVosfjSZjXWJsLVCSkGNDWVGhs2qjHeZNM0zHSz8Bm/PPUa0l5joTx
SnxhiOOZdCHtKVs3ZneE461uNsSrymtdqeH4rHYgAyXtw2W/N0arCcEK7WzPFQ4Z+BpJMiT0LGA2
hmYJ4tL7DYMiaq9q57lisiUnUbLo+t+Jb6CqIhfGvfveun6+PAT4k4wIPDC7co94xKgX/FqiDnHc
bxJZ4UK4+46FL2454D/4banR1qq8eKqk+pFxvHwEcE8kmlj6ywyikE3PpgaZuZS/ban+SpGmBabi
XbZGKXXUcHoXvQs4zoKeU1MWmRGUMqFrW4oMoEKyDsXvAs428rhFHN93/QbFLlMo6BeKbrwQuXTf
qsBcjdsu9V/l0fWN15X325E5om4ZYsvDT3sCTOtaBPmNibznzsuEOeyBtNEUJzvuh88NhLsJdqzW
48x5sZl22Rm/lNB38jot07p7rWzYgZEIcVKrmR5H8vqmNcRxCxuZY4NStp4ArjFMSjdC/YCJqAgJ
Mr2msiNbY8H4iMwEFSmuOnuNbNBchEEQ5c08erefUw31asjEBWEAAnhskc36rGkhj6vX3sfn5JqW
7tUXKLka0b+fDtKgKHQ8cOwH25/c30CdZkawja1cT1xNoSYDkeFyq5Pu+rWagztbm1TqpvfG2Vfe
9kPXUN/Bv0fgpMFsVpEQh0Bb698QGi+rJykZlbqL7diC08PE+6Sc6Ic9X9VY68KOKWHsEex3TbyF
+lixGxBURmbhN3FZPV+lY0EXdoJpCJ/upQpGDTxcLcJbKpKec+06JsFJi+cCncXnnzWbvkl0FQ47
8hKx9FI333AWx+yS03Y6Y6KwSsf97um7gA2PGUtll/oG0wXFFxZJUzmkmYisTuR8nfowcuNul8G8
W32pagVxkiLjh8OYrcFna9kzKMLTHcI9BHV2C98vH2w6iw9UAcTQe10X41XaMfmY5NX5vEf7uHYI
MGKjWiGmO22AdbDe/5IKqGFdxOOKgpNiAHGxx+/9hYm6Vh6+D1bFbdpO7wN0vxV+O1A16nmfe5ub
YPe0A3egAaM+LdAPNQcnPOEv3D1VEBZO9/7O2E2UwY5wF9aQq/cd2aCyLJgGEOuW2S5nMh2q4di1
YEcTU+qTBJgP5mvMIljdu1DSbroa+dEBcfbBwAz3wiOWg6JEEJGFbx262MiPGrV9jI9e3SFyqxDx
vBj3V6S0vvP17uI3EBRXDr5qIBNTOMJ9vLkJYacNjCcP0QfI4itFpwTyNFv23GZvFOrKOai0Nm5x
B8Vv3Oin/HSySgKlwsorIay8VZspFHWDflV+4OGe1oMS+9qk4um4+/DVxakAsqmJbwZZKCDvDtWO
5WDFsYAmsBBdJSyzSDqF1RZ1rJSt3O3RxJun6NjEmxNMKfiJrpMcDylAq5rLIvcqPivHfjUFgazg
/myJjDggOd7HvVf4KbNU1y+8zxeJdPjYwSqLdbUNoDG+zNuA6eKiaktYAMAEbDMVfaq7ptGR1Px1
qKkRVRJrtSeZzQDtx2mIHuHBSDO0UdnSe36cLy+b/tMk1AcL46uvlT0/Arq6eECDKPTnK7lrO6EH
Kj4EjwPNBAL7yKJ5m5VLid6FpZZPH5EaVXCQtDiNdF6MT0yhZhUkbp+zu+k1uCfTQH+itbs0Gn4u
BVrlQ82UtR7IvifHBP8Erk0nmcyUVwGu+N32byJM/KoryDiTTzILNMqo8f2LNpT4/gn86dswhwDj
uakLj1twLiBPWZ+nJOYqcbulOfKWsLEOazYgGG5TjiB6Y2f9oYeh5Arf+FwJkfG7gTy8UEqhKqtX
dfV00NvnuH8bSrGnfMhyzMX5oEtbCGNcimJKL3RsS1rRZf4zgyx/21MaVqq2rqY0Gu2ju+PL3go5
wtA3X9A3HuuWIK7KIgA9rzpmKabKLYnT9ZY8MsEK6B9SmhUl/66Y6LrJ/AwCLcUYflV515Biee/7
lsdaX46JGoVueK53yg7eFZPgb0x1kkXO/ujHTLiJfOGYgd3Vh6qLENGAi2b3dMxYSuUnr0qCbNCo
+v/xqZzdmdZwV96XnZ5cVmei/4IB6r4n64avcrFXiqtJJIZdBEG6O2E76lt691UanUcliCj7h6Qe
arT3OJ6EE2I0Qcrruexe/KucPoLCB+poREc7ugmmFebxq0T9E07SKJkYzwaiJBgor6yu5Ow6yGBX
AIw5TgcJHgTTYfYR7Inq6zHKYqiqV5qkzoMDHDpQQIdUV84MoMQykTZvKvwABT3JCyIlTQUPiiag
n+YJ0bawey0ZzpVFZ989CaWLkR9BWRc1/WJLhRWIb1DlZJjjiePNgq0jTLxz8AFD+jASmvZMIdud
NCLDA3ZTNL+Mn6cyLgX3qaJxdz5mMpojJ6oLt062ouBa4B7wdI+9qlgAbsrv26FbJs+2/jftuyh9
NimligZZeapEQEFCSiFLB8Vij4g8FsuIIdalpAk/e/8A2UDxafAREehxZAVtlOpMj8X1Smd5BT5N
+x6DnZ0yt+57kJHsdQqgplbZYfK1A/vucVoRHjSOXgTbeEWnRVCGZVJEt1lHRq0o9pE6HrhzTHa7
8Jz5V45XKLPDs2lfADDkzJbL1FCuzk+M0nhLojrSIRH0qRGYE2Z7OP1RBWdDsxWxPDeGwvDAn672
oExzXF69Dr7LRJ1hRHRN6kbZQsJ0GnLGHWNDvWJv8aoKWMCPT54mLhyPbd6qyDLxl09V1O9+sF4x
WjSOt5syd6iaR1mMIPzBPFKDo5bEXw+/2grWIJkKqkb0WIoUeuftJpMYp2vy623mzldsI54+3DYI
iG/YiR7yV0abOF7KitUd99xGGSEIP6F0qvaBe2P+NsAStFjpb/jJ76HhQc3vYTehOeZaZZEEQcyi
GS7HbHpXeKjLZ6i0BRyeq31acsSHHsBls10vaRfKmu4/QJwVxoZqSXPvxNq35Sm9FBWaYoDFPMm+
BHOEH/kdIQ+GZ+XWx0uX98RTb6AEsES3FW2/gLmDnY/dLbrII6VmKIudCkuJhSj5Nf59TSytLtmz
xy0rEuvsGAk0mdYjjfih+WpbEaqhMcPx60YCV9Dw1FYGHXF5Krguzeh2aMcHs0fYkYFKmVQxAe7H
xDhU2wPPnuFwmey2eoL1x/TKgwl5Ve8bVDQl3mjBMizPC7iWp2iML9Orwk6gaSwHcgrJKXhjiTXR
M4w9pHY25ACKfXLWgC8WUIRgD2u8DSyPGhoF6OwIJtKi5/7bqVRF8mSfiXSqjsT8dchQ0czW3qV9
7nnLvV+Zi9QnUXvRoQFs83P/PzPolI2nRRjsZQE3qfGiGfJuMQc4b1CAh2hROICXK5pNoL7zaEDw
J6VAYclFe1uo3PLrKYzqApcQj3EjDkY2Wz2eBXUwwvJ/rFhMhppeKSgpt3vQdpp3zj+UbsHFloRv
HUjDzY6vtnyrzWK2AAAX2iBUGBZcukX3SIwDY0lRM9NYExn40LDUEdEKC/ySAplBuRKhkeQtYO93
FpLBMAHtGuAejebnkhfbt/Z+oQ+3CLUeYwRui1ZCG4WYmC1mOQuhA9hf6DRawK9arGa9RZXmk6iS
UkZP4fnjyErcWPpjj3We52P8R7AGsFV6Cg7HCqoAphLLrMD4Tn/v4omZnrx31vLjZPAmMiM4NFwC
txNfD11TZeL3nf3jad8oiCyZ593r4y9LdZUqW7TWJ/HuAAO8JK6xukjNWv8emqkAAeE2oIcctquB
HAoWq6bNpzUECSRwB11kmYws9dT66CvjG271Sc0l5P4HUH1qGcZJ/KYeXQTW68/emgzAz8+DzUPb
OHa3x1pCM3EfIgiI2/McCaAHIkPVaOzxVkeD2aGotiRHYHThrMSeDJmJOw884Fjo7kq58ZC63IIo
5BIhFpUYX8tfoQWcZPH5pw/V2agyG8u/Z/At0FIHwQwT24HdUE7TzkaOb+OmY/ynAg8AKzJCQduH
uJkHmgFoaL6W9UNmij4Xuzbnz5yBGlu34zv6p8uKYJwXBVzo0gHj3j/6fI2ixcPb0/YQH4FjW4z/
LOy+yqdgGHNmwrtYoGinUUQBpwLE99AKrbFnXsrrslWhDE9UqnSfdcr07h9bB7wA2JFfamGiiQ3I
fvpUlP5NLkUeEIcHyegfJABTdsvbtcStg2cxvYR+Cq0oR14/36BrVkAlJ+vd4OvINmyZhcc3hIDm
Js5gHu3QjezgBMtwZpGgEdnR3Zl+hwy5jSuN+cDrW83YldjMUu9saPi0fs8EDPfwTixtW6QY3mr8
0Wt2tUjC6Jyn6+b9GmBQPGepsFwaaV6cyxMN+gvI5QqC5Bdt3DC0OazZO8qxI2BO4pvZIGdZT3hU
m80qL1uswN1OUtuUR1FDS8dTCdTqRJGs3W3NfH0wROHcp+T/b0pTPY1JIUFcfx6qQIoe/qZPtDsT
qho3oeXLjUEk6z+Vza/3+MsRDjZlO0wZD1bNs7Q2QqX94QjdqKyfxk8ndM9bQpdcSM8haQEdkV3B
Ob0qVkHxO4347EHae4Jry+ZDZ/4TMC3Vfsc4IoEzGAC2Lri5Hbd3Y5hPw+HtAxDsIW7WEVq8UEyt
fJKMLMWQaoi+8ngx3u0szrmy8w34pEsy6ConUDpYq4eWPefyO5iC+jCyXVi+vFyQ7lpZHCicg5do
Adpxai3v4Td/nNjZyjG+zMyWtXQwo88Z9Lrfi1ykc8m17akSOTeXy0MZ3VY8yUjQOrax6uHC8PYw
myhhfyyLhiwC0ZkRlgzRWOb5lPTkUOtGAjbdOPvDGy3IZBw4frMu4hn1LbXqkkv7zfQEJGUQ0G1L
GZpo5Yvow4UZ1nWbuNXxnZJJYyvB58HPy8PSQEA+ddSvB15NFaJnvfx8COj1uY1Q/hhL7Nt6wWO1
rttYjncN+XZVf65n+c+O4+YeFI67LAzxiLA/JhUXuKUuKpw1LzrousqJ3GazZjY+UT27gpP2+nFN
Vc2vPxiDc+7BI7pzXLKO6tJ57QfAH+6gNCWxcEhE/53zTuaXH3jZP5setlkxvxouDUahzgEzXZN8
PMHeVy90UCWTI6nESHd8wXHwNG3/Z767aj7LewsSBscqlJ4/SnOuJpiE+lVJ6VoPaz58dKIFlGfu
rUAjwX2r5KPfyvLZfJNrfCY6YeQlXawIFQ9hrw+6e/iwCwQJHch4yfos9+RrVSgJb0KQuKSgalZJ
mwv5kdFTFnNxWNfzIS472+FJRmvKiU4w/CUkJR4ynQuIRy5xlRXf0L8nQBTp4YJNxvBSJwb5LzRv
HjFkM1YuhWhpyTeAL99rgTBQ1yhNojJPJMXz9uOq5vd5JeqanrSKXR0BPOSNIMR4DsGcjMVNUDNb
7fb7uF6NL+oG/MdqbHqsoyAaThwC7tIqEGABKcZiWsSLyR56Y0QrLn/DGMdluRKwUrRDBUZF/sy7
6kw4UB+rQSYMYykJ2WcTpS0WqAO28SQC65IgbsQhHoA2n40Ej0k5V7Zy8AsdZnhqmtv8fGDk/NJX
gUlXinklOvbYLK0kFoxpxgW1kBoW9N3TUNKokYiXSOGwtKhQoHMijusH2nMC18TyjQavjzli6Pgr
yJ9hgKf9M3m+ACqgjaanntFYHRocKxD3AYgkO8/8SygW/pALb1hPLwEqFwQRRRv2SPp+o0vRAd6b
Dw9JFBgKLsHccquLx6devcHx5BJuJbC0GZo1TJOCxCgumi+6wzXN76+22FLJKvrrV2pSTB8hwY5h
ORJjIgFGCOPzKDjrcPlnTEYYtA+cLv2TyLxt6jAVh+WkXSHtALt9ESiszbR7a7eLtzc/wngaAYAt
eHo6ercZwI94Sb1EVe4A9sZXOiURVCS7GpgF5r3KmDI7UojTT1Uv3d1o0nX0XG0KTJTGSAfL5nqs
aRmi9ZpXLeuCFKmwxiP/oJaaPkjtYYR3mUKTlnS/Mm1Amf/FsPIpWk1XvEYI0h1uMuY64S62VNz2
MoeJgkdfukrz7QeSp53eQACP6g7MR0+KXRqOhH6LQ3LkDxervWAhF8DdZVcLG8XeefUYArvbsWNx
gApF7+vAoIX5/BS8LKP7NJopMtH4IsC9Xh0Q0XyLaIPniQobfOW1CZj82eTaLOTS7fKRa3hZ7lMZ
PEMo7TxYEfeDrYLxHlNIIIJ3qxgUL1jj0yg4WqV2zVPmo2pOl2A4EY9hlsr70++yrJHa3fA894PS
GXfDHkYtfNj0oVZ6RHr44Cq2GprQbNttaz3dblkeY/yvX0Bx16oPpfItPY3LYL9o+uO0KaDW9zpY
ZHP6EKEk8qMx543LZ1kx6xyLaoiNUI04guV+PZM7Qp8Y62y1vZ9gQxn3zZH+ETfSVzs3Q76XcGtn
vlKOXn6ycGaH5txaGcg7kKY+kX4PzLGh4IoiexFZnBAzlhGuZbZT+bL+/aguHdcLSDa1RgPjhmd/
Izrl3+SPBG1KrZ4BubFWiwQ8Y13Ax6gH0E+g/U4M4we7fXG16DxPa2Fzk+xcnAUtx/XUm7QrshL+
dpV+k2R0p9Cq3bXaWge6YoWl3yhhxzp/+jDrlCm8DMykJVTiEMTOwlU1YJxH8nFkSxaoGcylLqsv
Q4gOcN9mTq2z//K9nDPWUqRYCjdKl1X9Kk2eA3VVxD6QrbBAsi29OPUc+1jdhToPru1tQoVRYBQV
dL9jD3R1Erkde1xKawNaA9Gpe5nrM8j0nGhlSMeNgjkx1YdJV66Oo+/kZ32p9r5Jy24DmiuWiatc
vQAh4EKCgsSvjCvcwDZlzzKPmuNX18KOvfU93Xyync/rw3eQGnDoYGGBgpfuBRaZctBn+JFDG7Zo
3jiKfVZFsMh6paoZFIewnqE7iT2kel7bB+04cpcHb1LuaY1QuiKkYoVOxNCUJGsjWh7G7G4RPx5Y
uGQSGwL/4HwS3ncCh/FiqCvwpi6G27ruanlXomdoBiHRbgIKuZ33rxe7bmPXDSJu44ss6EjtCR7y
BZVx/9KrOWrhNLt3+84MGCF0eVaGNzFnPFlCORRfsTXnOXnZ37Cd8566zd8UhSfxF1kG2Twv0ohX
mHkfOwOr66yd3JEa7FaJs4n8ipn9c3FkoaMgO3FuZpl+CUQENo57xZ/AWlBYLlkr2zVpcPrkr17S
z0E33EkWRzNzO54vWOHsqGIGWKTT0LzduTZdMRt8as1HCSABVaeE3Ury1iD0HYY9VTpaxGT5QPGc
vpIGx7Ih9haOSJ2Jh3KO15McJh4vQP5lE3KL/Dbllmf5JKsVbY/V8aPtJodA47R8pgQlL3JwHZfe
VA+gljWhoqZOk8sjfZ2Xy2dX96Cio5eKlWsauXLuNHP7DcN+nPwB03gXhwCU/Kt5eewXQ7222l4o
b5rAwWwTfKhBu9OXFN5QdjEb5eiEvd2+LpVYRrm0IzhGSihhZ1v6iF+A1q5J3BwjsXj8CkZ+/4wE
7JJTg6gdekOx0lRbSPYQyfvWlbilMRz++nd1R9LDykGl5aZD6gqQ+454vhuuyGtZi8FMSGYbP6Yl
dKGx43RXPcgwbUaYT3O9nHXHwwsVkrsWp5SReTIANVKwsoq1VK/BFEH8Z4GbvdLwAr/OvzAJeFJB
QNeWAJTHUMaT9ol+n0CLygkLR2bYsNlWu7G9Q9G3YZDUqC6q8zC0qwOMM8JyJwGesqyrxfNRZ/mw
ns5LiW7OXPBK1G7IU3J0dup5Sy/V8LQNGBKn9nwtD62Lvz05/dw2mDxC07JGlCuxmbQXcbawknfV
7koIikPk5yCiH0Wxl+KcJSJxS/7EoEFMGXkM0sgExrLFbc33NYHwA8QeaMEtXYDF4KezsQUWIA+m
XQMzpJDZJMlJzrwol90xHKo/gOgShJ7guBGlA2H1dlNQpa8L/DNFuHHsfHNWJXypBYcWuiJcuqRd
nyqtdUN/Wo3NVieyJA2/qfSGKsDdDcUQAkmMLfwtFov6pOEKCXAOkO08zitq5Bf7hlyGjXTuC++G
LV7agTxquPi8iernCpDLsIyaOU/hRSE0ukRdtIS2XzRuKtckvtQwxFRbKDDTYedWSt8LjRDDN9KB
e97lG05YhMKk3T6btD6L7hsphD5hyxgCCfzJstd32Pv1Zl7QEBgOjicVhB0QkgLSdxFlyHF+pozA
Tr62Px9ARwENcQ+LzeAEiJOOvqpu/HQbma/LkSu/yYoU1gB0nc6apab51B8tFSrWX6TVBsZJkh+0
PWyD1T/h8QB+TqolAB31Wg52uAYc8pICSQkTNfel8M3gx1uN1GJPTNEP+AL1G1IwlBBPtDpUpQ/i
NJu47R3T6gOtNzTcjKjS81NwWHgkbXcq5D/P5c05njFq6+YHFBB4wGbuZLYcOzyreyJeMjVIYVrP
l+IRGSs9UPsHZ0YA0bJpY26JMqObN2MRtkmWvkmtBuCJsxLANOtAp8vt8719UkOIw/Y0Ul7BsANJ
mJwPLo3FsUjv1dFaSDonrBGeZVEpI0KmsC3/vV546CnHW/M9KuCW21vBiSlmUClBkUZkyO9GEri6
FYThI7T4cIlBk9EM2yj0gaqq4fJONFnR+sjAaGSaVJObHw3Zz/jfZGkgDyE9cV+YtCnCR8ad3cjq
Ft923wUAXCZzmqSxC40dwIE1SjHhzQtNAnN3OOfzjmI5YzI6LuTNEP4HG9ZVrj1+6bwhLG0wj0Wk
uywQUuBqxaCcgzoYwsbi960uAdWYP6GBgCYU31oGbYKLfcgHRhDVE+ijeRHe05EnUqJ6ur5rMpS/
u4eSZUz7Jo5yl6VOLvrvpXZzxMMfDKkEs2Z7V9ll5kLoC8D6YgozG0SRrgX+kBHQgBUTgH92VC0W
eL686GNLeWnlaKT6bX1ZjXgxF/iXsD/5qEcJcSsyOqjcEVv3H5Uy8KxTcB/rBG2nCvqAfuMMu5q8
obE/V3gohm/xeWCTUpav7GhM0ZkYcaaM3rMubgR/pwtlOACsU/7Zx49MMTFoWyWn4Xs0HuuAC/QY
lke8BFk6GqYBq5i3ii3+WlezbNdDmWVhJWNLqahYbaJoj8tY7ELqA5qw8Umq++Co7RWxNDd1nTEl
cHiiOzMrFpb/iN6FQTK9dNN1I89RibwfGpMASVmkpI86bis2NysmVeZGrTy4DLC40+tUol+r2/FC
DNIUaN5AMFHtfoIfrVDSXWG03IQZfEcTA0+tQZBdIQpQDr8Ni0I5ZqI86E7dSnNWTtxQmSgqA2FW
Po6SI1lJvnGU3MOQYhypRMg2rzp7TntYgcXY+vSah4vPXhJQyBYubX7/lf4DLt9Wr+NOS3PccssP
C6nmxXIM3S8js2xX3btkx9mKbbujR9BNsa4/HayBlpE+pr2QGyr8yzyFnU0jk5NeupIFJ8LWmKND
+tDowNGBwGsAf6CohbDoGjQC5FMqln47m96SSgATBa8p5ug92UjmiAkONOf9vfa3kbv+6h9tnV7q
JHjZ9fXy1AJHp6Oe5dOMQxXBNPTbiPXTFWZ/XXJQvedEE8XosEIRl1UfK7gK8vb+04xLXYx3zJ5v
wsZzMs0HYoEvDpDtamChDhASeceuPYZZpSOtwdde5JgnghKSeKcVUcmL6yfu0NMe1JDsTOV02SL1
ptx2U9KAS2exsJvMbPQWSonvZM++cBdH+E2CNKMJJeFfGg5qXtVus6396zZThD9HsvRyj3BBXkzo
0jVXyJLWVTnRTHZ9zCbYY0c7SeRoyEEHaOF8fcDteZGnVMkAM0JLzVyj157b0yFljeiANxa8oWBA
NT6Mu/SKrX2IvYLMo+7CKJY+WqNFhpYzAe6L9OR4G2u7TwN5A4JNRAoncgDE9Jox2Tw92elMJqoy
HSogfDU/5GzFDIu1RXPsox5yvXhfBFXoNIsUUTfbcF79YB5s6HZmOlr7UdDrem9QnEUqppZqB4TP
dlHtkc6OBctT+o18EGr85zehHq5AXqNrSQzH2/MI6EXo79XGNTWFgpsOLqO0x4Sbnu7AlJn/JWWZ
yC5kGtjMaluHA3hAOxiPkRp0qY+9spe207CZX/OxdquzlyZcC0MVFT8rVQwNzoqAglkoqk1XtG9+
XiPxsVNapT3RG0ioTDV5la+F9CC37dk2hNmUVK6LsfYhENtcdbDoxB6+R7Db00UV1xUOallBwbXp
fnYkpnCCZ9U+ydzXe4QkOaRk+tkwhvfiV2hIRO80xnmtWFY6/+0rZxbiCjh6EF9lkbWEJ/ERehfD
iORmHdZXZBzb3UPDB1a+0njIVE/yhqFCHvQVoCH0HocRaignr4IpZFtSXXcCixy/ZmJhTjLLwqdv
OLdzxsYyOQvsERq1mIsJ43pIhE5N/EXElyhzFRkJC7BEc4EV3QBpcjkHimBAG3Vwm9TQ3RRfpHkQ
hYiWdxn+loOyrPCdiP8xngX56ELmLxJQp3KUoSCwBXnuJdnCY3Mz2kLMilCkDfo40GvNbfTXXzKR
EYygktzOGSJDeOompoo8wxeDWXSGIG1ZQecW4z28iR0sYaBHApRzKvP2ARR5KJ/TWzpSkHNonIvo
Zb2LjBIp+ZRm8lClclhK1uucLsglMUjLG3+4ivMCYaINPNYp5e/3QG4YsANgOLaBoinji20m2xj3
pHNFejEi8gb34qrwtiPxWxoE+wpdOemQa/hVm9OixOcBg0Q6YHA3MNiP4JfxjLoJpZFeG19C79Nx
nXiCsp4HxP75js5UF6eON4xwQEEkX15fLOXykWtB+N4NMwBx+SrXQpU/CM1StG2mWVuyr9SEt0H/
4abUQWQMk9aWlOiJF34l0dowVUP1AuYQjmtwx+oOdNnIZ7J7sCCxrHVS07MvE3QoYu9JzXW5UZos
QFJ89mx773DAjFteHQKMrFQ9qO6OspOGqwVmdXtQztxs2DzCmiObCDQtYPV8EiIi7lYJYllsgluJ
pmGJnR3Oiox6dKqeF/YyeBPQs4gaokldqlUIzr5t0n2i1wjjmm62kJN0Uf25OfQ50wOtywQxLSLA
CNse/s18lDjHDJZHG17dYf8J6P2gUiRboRjwLnlEiMeCz6h8YoSwLzXrX/Ix9LH9spY3cbmnTQBD
jy8MV+hM5CaPis5xVSb4Kesjpk90V5s1NMh2OT+YV9yUaCFsKG+4RaTtLonvE5eu4fKVpxvkGYcp
SOGC/J0YEf0F3NRW0j/7exc/VTAxEXHbvys7wHN+57YZBWaLcIaikVovhNDepzZhaLtOn6xuM+V4
sjShH7tT3GGmPI1i7BTjXSgYHHdGfA3Uoihi17Qq8Q1PhiBw2dH2n1DRjhS/+gntnf5M1YFsLWGm
xi2azuW+uQ+uDjXQ4qjCsYDeciLfImm8aYuavGwYNuxAs9LmUT67S+gfXC/O5ypSBQH0icu3mqex
jJGnb2l46AU8K3xbmOPQ8VVQF23E0xfbqOKBC7tjWaCy4mElckGIgSe2wcmEQxpc2qSGjKGGjS6o
ymlMOlAyoMg6IrubxsIArcVO4kv0UqJSR8Bsxs87mOeiboNQ9oqhf0X2nRTqmuP1kM4f3JL0C0nI
8FWkyGQhyEeJ3yVRb2INgWUpcs2JN5d5keSe2goanOuJ8kO0hmMb/q5kMITAqaVF5XqcXaIvOvLp
QAVy6Tb1yAtVDoGV9UevY5N+mew1EelL42PEcG/CvzaykBKUFBzkiJ98fO3VO21n/JpRY6Gm5fgd
QaEc5CnZ55zbobLlmVpLwqzOWaUIs+bISH2kEPZxZAt1+BdUSNKhBjExW4KJ+usn5GK8Rbj25DvZ
vVU6IY4Y/2kOlc76rf5wIs1PYc7/wLX3qrRPAXYpB+JeDxWiT+LtnWKKR8sNJ7Q8cDNMJoHxo2cu
lpf334s6ljzv++SMpdv8mOLm5bcT9CRskbKkvkTC8Cl+VhuOyvTpmy7/fIqzvkRALrZEhcL/WW5t
gLV3aGAncYh7hrj8XBp9C2y6ESuMrvDDiGVP16YURiwF5LNKLjsrrXKmxgCClcDtftnfnnqrOPvH
/1czhnmxZ+PXhMHLwDOCinVaY5Ked07iRwQKhnuZcF3kLL+kIsAiyYujgEGYF20wheQKbnQwDwnd
+qS8jj4OJgl6EGt6cAPd+tR6wpE3Sh7GbjjLpm5F8F+uKu+Fv8N+0rLnanGADaqSXMzpbl7jBclh
jzYgzgt+c7U+mbl3QywTWWNYL6FNIxy9A7Z2oVA9igeHRBHoJBq4/2tvC+jp648gfDE2Qd0Mtpnr
p8oaayQrUy+qH4mlSbfwFjGfqerYfwv8bjU8tFR85Rx219Ps7k4DifOEi/mOUmaaRR8KBDPemgUF
YHV8EE45uGQLEdQDy1kbg/JCSIulk1DRfCctXBXCuN1K9Vsj4+jIHUJy17ibYuA8oIo9g/Ny22cg
HZaQh7nEI+VOCQhnKGw0bK3dFf+KBrLXPZAE3hC+BQH2y4b+JctwE5R0IcFCnP++uyz6pV6EPrxv
5I+ZLCThSCrmvHnazF90zwPRNWmmI5JDgWH77RUXPjOaRecBFzYl4u+nxC+sgAzNpjJgjybtsRPM
eA1muWo0WvmI/ggE6jLYyr6glJ3wI3a6kthuWO3BWDr/VgPT7erO1VB5rr5GEI7LpFxk3ZsZTo8O
ar2s9Qo+J88fKaQ1BhzI9aHmilV0CyvySXQN2KKC3cpUEnASDLj1ll4qyydkaiNG2eUicrlDDIjV
yODxIj0JYCDjmre/jUJFKjMd3SXtxqf8+Z7vdQTUXl+EfibZN+SFnA6WvwCX6CijHKFjqmNqGLrb
GppwGSI+pHXOOqJyviZuYx2vkgrOytSTC7zpcrZaiAimvlIsOa3ewIFdSOIyqTHrh+UFxuAmhnBx
mC+GSCWGO/YiAbR87GrEQ18Ah+qyGeYLwtcdgZD8n74N3q+FEy8WcFEohDIkdxxmGXafrc0Sa1xk
OYRTwweF/3kjOlb0iU2CeJudKJWAneCPhzun3KrUM3EllaRdwZXSnrDL28HCxmfipbpOgKE56OAj
vGsnAs/+YpifLb0+nrt6zRTmiP8Jz+5mC4Ai8nel77t+9184issgFSJ5Tw4Qi9jJq0jOv9qRoe/3
hCY4NfX8OorGBSiCD3wUdw4n8dkd/vV4G7gHk7NsrnjRlw+cwIe2cWimncvkx2tdu3NyzfmfiFwS
UuPi/2hrkoxIfoPMD2fsAu1ONTbVzfCcqPQJBy4PFGcyY36tHcacyNmt/Cfn8s4O/XHt5qMB5erU
cmJP7FuaJspxiVLJXHZw6MNsOfZXufD0DGVyFpToTr02GewYrJ0jJnkl1u7wUTx5PafjLM7lGxR9
fF9Y0537vZ48vwqpR/C2f6tbVydh2yyr1su6FsxDpssLCc7wjSjBmEO2hFZYXJJnUzG3YXHZuakR
CrxXoJvPvaznRLzohOVZyeiidP76G5/AxyATA6vU2uYj0gSjLHsUMy2qiuryek7yXaJ0BNmHWTmA
lrYErX5TttKuI5sjCnS9OwdSUHbaodZ3p7vxMZUNHPP0MkAjryd6puKDIBYeeYpxEq3qkjuf5KFM
jIoVndeuXG/c+50hoYS3SKc5zXYdX8Nj+92QhFxVOf2LiGUUKiwnGa0N6IDwKwuJSwzXf8rrT9x7
0xvxKxAI+bgTVSJfPdfjxHjdEo2Q5F/kFhfeCTm3YXMB3NYk5tbi9f0jzWQkf7pYYyAJDvx0e0oi
t0S2PrXNYJUj4Adgwl0nhajhr7WWqd1cYjCIl0MVEap5aST2NVNwbc0HyexunvkPSmquR4qIwmsN
ACnQmtCkhSpq6KCaqdFtIQwugBDNn/96Lhxd3hkygD2OMWn8LnCGFSFeI+EFccKjUmiC8Atj2S8f
WO8JmKdLFyT/qAepTajEk6Ct3PoMt8sNYWuxkmJXUTZbwM/TKIK2SwcbCyEjyFbZ8/ngT/nZ2/FX
k0OmCgVNj2SOrvsfIavE3Bzt1b34/5cVmGLXWYimnmxjzNDMpVxemmhih4rxDuDBaF1MIW38OxH8
qP5CxutzaZ51gnyw1SFF6jvi7gEkHaMgymxj8Lis3Fi2di+vksCRWO7fXYjvP4qu2NjQ73JDBA8c
sPgL3U+sgWl/Fu4UNiNU/oERX2m7Pzt+cFt1y4WzwmGQTWiSloaApZSkBaFzYv11AunaeLB20LBs
1/aGhNCYAaVk8dPvUkDz2L4MFWz+HvelRfYXQO+5Ux2N7jux30Pc52BNVGVCN/Dr/jq80fd+zO1Z
j9xtCFhz++mRwiri0Va8s2Cbpc/rfkgs1EDrv8Big3yRiMpMxol0cp3EJeSrMBLvoKVTXf9Imbov
DTzbLSZBxfdlbLhZmXc9zm/42OZ7asThM6WbWD3+OpqFP1sZVoDPz6RPEDQvZfkZUjdiWKINPtiA
zx5aNspk5f8sxoShMcprABCOLUvYA9U1wpnbeadrtRP382CVt2NJ4X07XPtAKXOiHBjW/G8KkEb7
+1qa2XlrpltzmmcWbl68yoUZeRfiC6CHfFKpjuaXLxWE37j09AvcVp4IZzy9tJ1TQTSxU8nc9wsy
PNI6EcehjPPx/h1V8yOwLTwgZ65eQ0eR4PCDLNhbWdeZW3JABFJA1F0Pb1l5wsmtcK2R5+nbC762
Q47iwLLHJF4TMFoGymPNXa84bOMSmP8YM/MA4x0kvN+TCrtZIoOlNwzS2c2osWuBgL7i4s0BijxV
r+SaDlfIscAQiGr+18xG20bNG1O4BbVDFTKJLgRdhdcLMUeKvb/YkOP6WWmXpLodfWcTZo7+0Swj
VIXdeh3gzV8iDJLbnYD53D4fGp723xOw1ZS568cxhE0aFh6xBPVPzzEXp9fl4XBww3BsrvTr76Jw
ImBPgECsuGZIp0/DfI1YJ1IylSb07S6/uHk/ePzObRCyH0bI4uWRIrL9m0vXxndBm9Inq1u9lq2/
Y1/4pXqpZ0MUpHsD9etPSXrUCdRU0TLfOcmyYQowuxydsET94wZLirMmHWAG1ijjS1MLbHtwKIij
j2KFTeqOgqxObFW2Dk8WyJGP405DOYgYQ9Jyu7DfIbeTHJ/d+hIF8cqutvD4tvKYrqMsHq+Jgqx6
+0VVXkGBZUGbPPDJUaDgMAtHQWte2Komsvzip5dmBrEWrkIiKDR7tLzCRH3FgAVLn9tKaGMRSH6l
wchijtMtPhz/afZuUlJAVoeroD5BhkNhmqhrZlRFD9OcRIyqJZyhGA0RFsgEdC4Zqxpf5K3zBtbp
vVH2T1CEgUL/Ie0gJDwJ+xtid2HQ12o1VojAaOzsxVjV4WDT6+wR7AjVgfYNEso/9jgNecIzd2mq
9qp6eR5a/UhrBnZfPhCKh7k2r5/zx+1HnVO9i9DM3L1ePh5dROeX3vThF+o/gKjb4KYAxoBMYHWA
Mmx0vUFQ7F9M88q7lLIMhsY/3hCnFt9Dcsn9Ip0W3kr2CAdfKufkYsWzbPHCGTnpuRntXWmgyI/Y
45Wiq+6k6HgAlh/u8t1Aqu17RLObHgrmR2j9N736u3EeJNDBbB+M9BhWhVOQMJUp8JwnIfH0gHx4
KO3eT4C/JmP5Yy24ERdQz1IovRAGkaeQ1xdrj5I59fsb2zkmvAytyF1Z5R2gF1qwnq3rQaOkz2va
4VhIdHKnbHKlTooOhbefD1PfKysHFBnGP5zOWds2FuO1Mx8vKwINc4YkC7jpfcoQMTwVFBYnmvdq
6O7TTWoBY8493c7/QkCZWef3jUCzkrahQOzSdx4rJ5hW6kHyN2lVKGHmieFgXh6RqHmAbcY2Gefv
LxgP4PyKT5ay6ClXfcHsSGY+axXZiUczoqDEV3vzq2fIuvQ3yq9enztTyJxVw9r2ReCgFMtdis6g
RvtjqTsOC7djf+H4eN9qazERf0wNRixabp95ooTc0kCqbdWVR4eWiilYWHFbOd5Ns3n6Zsyux09A
skuMrJ6aCA2v1gZXkCy3cfObWsABtLnIlWr9OQQ4d39MKerHbR/H1Ro7Lm/UPZPDYw2IXOny54qS
ioAyUmMzkyMk2fMS8gKvwzx2UI5yBgKu3s4yM78l1HOJ9eFc0/dopayH1FXtMimlpSoKrcf/RJEd
TD4rnCHleeTct+Z/8X0+ix47HlG7adW+dCaMVWt+F2czS2msH6AWz9VTIjv3ZomaHL0FChp4cI6r
loMhDpkURVIcZFfbvHXOpNXSWGmSLz9hvVCKil8OrUB8oAhAC75ABh+oNMMeszdtXet4tHZ6burf
XR3nTg3jXq9fnetxfbU+BEgZTVu5iDuGqkRWE9wAm4uIiqNPscO7NhsIU/Zbifh3AJphu7qwCuZw
5ybvE0s583w5lA4cNHbrOYOcHZ4GyR4tJgNujN0lNfEUj2OnGwrmErZQH58NJypycvWO6PsyWRN8
AkiGPZyJtO5Bwk+K48kIl3q3ZQ/E9j3Ugu5SyUKDvnoxfgWPbNAN/Epwj1of9QEICSpjfkuP/zCV
dGvcvBFys17qapcAKewrcfbj9mXzoapTU3ESxiZvXGiPXfy0Al1E3lHX3jsL8v8u9BLsllGOGxos
SGXzgI2G8crbUL9s9avq5LcxxuiqWmxjfpyE8OhUJlx3JIEu7zD6er9id8Rv3t6nDVH3HBWS/TMH
QcNeG/xzj3qv15DIeBoR62wGG7ECeB7ofXXXKw6Ss7x2nIK/zk9k2PVt74xGa5of/FJXK3FsM0PM
cwpJWzWnurxd5uezO6zGRVgjZeSzyJ/DLisPoRz9v/zpSQ84FBK/gKMmUoGcQ2F1JtXYO24RdPNG
qgAH5IuOmtrj6+N+3+6+tb9AMRW5rX3CDNMFlrFuVCJj/azOHrwK21XXFdkjBYvSZJtHDyBF1VnC
coBDEcHYopI3pcduztrcB+rT0IC0lhw1TQ/TYHlzkHCTOkIKVPMbOqHJqQKVoTZwZqoa9bgvHBsa
mNV6BR7uDG+/eyLc7PSqxNBdEH7Qj9Mfrq4YaFmIGqmvtCEYFaLhByMBOxeTW6iD20E05jsZc2to
chX/XpDDsvStUr7Jt5OzKbQ5a7GsjA/CWltjpBM9Y/RcdEUErATYY42fpT+imuWmpp+QqGXNAWjS
aGvCumKz0zy5hUhi3UQlzsrVYPDslwnX8zrcyBT1OYwosSYkLRJXANc9Erm7q8B3zOmmhPTkV3wm
KgqeGlFbdhcBC6rfuN/fVuoJ0R5DDTyajlEAeVB/RzQS8wGiVQhVIzHQXQjFU0TBwQfKRbwsbY9m
t/48HMW3kRo75yUkrbmJpjeQJH56kO+/SeIt+5Cw5eYP38+AumFSJbpCzAQtu83+w5h6SMNKm1Ed
yKSN1q1xjXaiFRtAIwP/DLFSjtqKFwdJJRN8VclMu1CiDizVVYlYzPkxMLq36EstUH0XiHKfQa3U
NOY/4hCdg8uvot4Jth5dolzML+suEQGych3D1b7g+a5yQm7kTS9mBSAA7+uG3G9uVHj/d+Mrho8Y
YwhbBDCfzyC3s+2u1eUcakdwwWPpvzLLchY0SeU8y/EcU5LYICOeX6SB43gTFvHqHNRtsdJdskMX
UQioMHYekQVDBYgs54zuQD3u116NQlAiJfatVsgf40IH8VNf+RDl9vN2aemRW0jv7tFecuFdyzI8
3O0KgtduOvUvZ+NCBwwooAhNa/+K5s6ItKtzCeN64jjAyIrmimLKs3keGx1kYkdvUmuwiyS+snYt
HCDHjlZWVrywVLPhuGq17mziUGR1a0BWPyW22iywEvZXGjGXOveiA0PcfsbD+9qSxfU7Pjw8JPrn
k5fv9Gkeavhr0X4XQj2ixD787bDrxFsRkVpQMe1mZo1wXGs1uZ/ZzaX2tBrEq4w4nUkhKftbabY0
hDpPQi1lFyJiZ4C6QgbGPUjZpiM72eFnC9qVYdCCt4qpOASJ4eV/if8BnUpJJy6vt3WekjADZl4T
Y/HICJIx43UVd/Kk5rbZmx6uKO92kTGA/2Mouuira6FCsred1eYLoQQymVT2neq65xQWbcBfbFzX
7uMdaoF8DZ79cvC2s2rFaHElr5IH81htG5BDASbcJdASS4S+DKdzmUGyTqSFL18aJU8ZC8bVjmjk
DPQkgXO0jPF1WWVAKvPoiLsLBd5mRdxGYiZVT8SvgSweCySWtwuqj5kRhsPXtYUHN5qtATu8U74/
hmjJw8PJt3YhXWLLLlNekNSQir25DswpnDsy2Gg4RFk5SPCIa7vn3SxIG/Nu/ig3eLfdUllSrZ/A
cDrlVyW4ss4NBT/BlROqthRrenA4RftZ32fJCuaVunHc/M37Tpq5hf8KsUyX5UytEj0mCd6PsQVP
LpzyLc9n+cLU+s4w8lJUGSWr4eY3iuUEU8q7BTqysAFy5myh3hfokVtRkdORTlvxExNZH0ZxPJ2q
x3acMn0+CmrVOIu8MyKOreD+PjUwTFxkMZjVatFTE0fdbJDd9oSu4l/zpzYIgFvWtbM7xknLphvI
33C4bV/fr2w2fHkP7k506LvNQBzI6CJH8RopIvWzJivTJQubGP/ylos+1RkLOAEzHqxO0AjpK5Um
9XIzC5W0LzruzZ0F315yPsXqTvRzQluWaSWo0fEajpWv9Qoo8DajGAEAOUBPies4RnruJASWyxAC
tA+Rp2X0k/5iXew5oIqxeG7q0xX3Gs8O0aJyFQDZq15hwdG7lIDsUJtNthRIUwKpHXEV9gagGKte
y8zMbjRGJ1zKwZel+4OHQmqzAVj9+benmJRM0b0/tL5ePEGlslP0bAVt3hTTf/UvLWvgBTAgdmgS
YOMZ4iVdxVIqmT5rppL93SND9f/BpZDYiaqIpeZB/MZ49uYg09fpouhK473oYNyyQN4ySHdgWSCH
JL5uy9K5tJWZQBmlByyaFE5AJT3LXHp4nr43vMdn4UQZ3nOub0wJgBcZ6lBQPzyJtcOHRo9QoxwT
St3RlvGCdU6s2AeqXZ8er3Axe6CkvLr4J8jTbeIwrsSDzvvIPHHXqUSgXO8FZ9x2/77zDz4/GwrJ
WnRf4oFJnL5A7tMJvAottXMVZNlWWc5FhkHqecj5geehJ416YXAhB/FFQI2tGq277crfAz7xIyxm
vbVieYfHZSZfHQqBgqbHtoqL9lfsoFzuTqdu9snYrdifP4aNWGr401q2OMiaGc2DLx4EMwW/CUKK
q1zCl4whNRPeUVKt+QHtGHqBFGbcGW7MsFaYmsIeATmoxYZusedmQyl68rnn50mujtK/8+2Ug9Qw
1nk2T/Wj0YQcO02ZFZDzzNa/EndyVUH6KjKhyCIrq23DtTs37o9Oz9cDWLLa818RwAR1PUVAjeCd
b1w+bdU093XtqbLng9hXt/BWmQiq7/RBdwyzjGDm1/2VOXO/dy0oGIRivkagJEOCSkM+SUcw512Q
sQVRNTqhd0D2DjVnpkajCbD2uAYJCLYgt1DZnoiCBjJMs711J2zDoO7mgraVkoX9J2SmqHJi0T6t
lNCEZedzG+Ot4/JRz5iuVbi+sHFO0yPYLpbnZ8PV+6s7/4INfIFslj2VBi8h+2KHJipGDS8GlP78
/rHlai5rzgcXi/sSjhwxMvSCnUNd9XQoTvL2duprs+DmG7Q4NUka0ElfCkq6te6BL/UB79xrGIJP
3VebE8trjGbtDQyGrURi5qKFxhsufzhVOwYllVu897BQZ9MK+N9QO7Ggsgw1uhA8dOmY1lf461eY
23WKImZlyZmaqUDWlnBb5KM7l0+F0VGsZSfKcjNtnPLS6Xv4OPoT7m8XzhzIszmE8iUCQz9GFeHd
uDx09pS3uEIlamsRoyOfiBWjyIZ7faE2GoEUYTCAapApaATjkD6xVR99qlIBJUbdsoRkwpZ/M4/t
CfEZ/ro0fPRQCp8NOA5t5wV06vC893IMwGCblGD95oMBldcDP3cg2gMgOPxk/NbGr8bbizKH+hhc
3pVnhfl+Cuo5F1+DFX57fDXaJJKNhU+ZNemMKAhZJFKW7c3gjtmJYkI3uVgClDnENns78l84c/Vq
WrjtJgC66WdifPRaAyNsm6uylEQ9fVdG3TY4RXuxDU3HpInD+LSXq9+RyPePWJWc/HN/ldzbHf8g
0AYM83hU20+yDbssbENINcVUgSCpyEYPD8M/he32P1YexRQ3nVAxW2XvdMEq6KRbF6LUJlzINA/n
+sN5g++tMUYJiEXlN6FodbC+vfpD+tUqw+J2DpQVKXRvyFsiyZWiXENiUa85moVp0/oQP5GTwkzQ
Y3mOC3cOj6ue9mZsekcEUNm+0Xs9kNXl90BhxHcD9l80N7d+rCZS7LzdiPwUS9xUTvYUePqZncC+
NYn4o83kcDSjH4wwgKb142m+GQfwXF16GayGXVMR+D17aWSTJ0sa7XGjncMZksnWEF3oK9d7OLyJ
G5LWF4xGnKoFmOnYREMC4GPZvYqXe72gLZbQ7G8zc2UbHlKRs7QvHfFOX4wJn4gtnYJEect3KQRx
JLX1F1FQKsNYx/jAwqkElRztqV+Zlx2erFo/hKcfvCvRRzq6XOHEzIdFNlcS69ff/r7TA0GSe61t
hGAKvjIHYkprShppgUCIos3hY0PhK/CXQSiQB9HGibHbQ7IBPLS2lLkW9hk8EkHWj527WEDyeZ2z
7bVPeNvUiGGtMqVUlO64ndZAvbhuIJH7BwIlXKb/6XveTM3fBY1cWjJDHkPezf1RiW5dwAUbfUXa
BVeki0AjQzRKXenjCJVwZ3+8u63WXk2C5XXts7YCX7uV1cLCpswNPS3SjT7QavUpDwpsAFAUdmuG
lwNpvfqHuWuZiSBfHPMCkx5CAqGwyP14xF8sSh/bi4KSMIMDEIb2Bmk9TmKFXdDVSDEjmv5IdinB
Qc0exOolyelOOIjwsH7natKw2CtQjoEJkqmR3iiFXXmbPV5u1tsvff4j+h7H59C+Z+yKzTUlXR3f
r0uy1b1wfyvnXxfWUWL1Jyd1IgbWJsJ6uSha9kKUsXjvSYxjf0G1QH4aMU5XWvMPTWb8U7LpU2Vn
PJCav8lGB4/T0Cmb9l1u6JBwRfdEKCEanCo81FwOAfD55PWiBGPNySZ10NK01qgC7XWoyibLnp6e
hFjEI3RrBID0CzpJ9uaRbmk4O1O8aKfAU/JrhGgB1IXMqwvEgvKuFNyHFo6hTR5jO6stFXRMuvjJ
zGXW2pg1Aac76fAE23tQ8A32BIxy9wqk+8W3BndHlEOoGrYYfieFpyj5rZhu4ZZuv0mGeSDYlwHz
T31l/7URd/sWxnwaxPOE5/g15cqh4LeMwGwCxtI16glLQpTuSY2l0nz6kqf74VaPWcOvqSffpoBC
fEJzMWPAD3mxAwM49H/LwtHN6Y2osbpRd/VLRapRd+A1n2ZSrj3HzDS22uA8stgNYiulDvK0w0xB
PkqTq3FkWkN2q6FD8IgcWxcVF0mepIWShXmAz9EhZfOMMY8l8fNqdr2rhdR8tL+X74E4vVrinQ1x
gfHT47DyUYxIXbvaTzvKUS4vtTx+wQzJfJp77LonaP2Wvw0iABOSyZRUpNoCu/H/aoBswohvGvDa
nSuC+hshi3uGPIxR7A5lLNVJDhcOZ8vbGPBJ3q6hVAI4A9QoHMyIWjqEJFFdE8eY71HQXxYdgk87
I5s3G23U7vHHpCTH3J+uxVNpygZVVFSyB63xRwI9o1nu/tkVNX5MzSk84kg7xlTeFygKiNN3iHJD
u3IfzA8yLGBusIAztwXuQUZrmfOvkEXruQkoEpXPV6PjX+SsZ+vCMVhWdRg/XGDcNPKQn5IS4ZZZ
WSprF1vgJEnA/YKe0g1Ls56/Y3EYXvk5smWFwvpeosCHovsUmXOlxHAfMXtyEVtai/Ua5MhmDSNY
ItZfKjkoeVMclalKZnW5cvBQXJMlB1JiyR5Cgps5mU5comU4MVQoShBesmbBfQrBVmPtjrFGy/mA
uhgBMJ7CQmhZ6+/noMhF0lG7K7oBkMKJ5DwHJJvZEZsESmrrZduyzvZmbrhkbaxmZyLVQxQaukqH
oY7fG+FIVudAnWX08WfUYodBNrP12o7TuHkj0sQfGPxM/9abUOFD6NLnZlS6TAuLtmj1KeY/c8fw
tmto5758vwVIeYXeC8Sfc+DPWKNMNP7eYr0NuxvCTbRDuteygTq1/tZUQBYPcr1OTFAswFFRJo4c
Z6sDYkw5g96O4M4lqE1Bf6Qcuog03pNikx43HY2Ha73iBz8mTRyEf4JApsTM8nBUpIOpxCtKCD3q
+984FRW9NZBIv3UVTno77Q/CdoFpZRLIF1/b/2MutCFg76nlC1L81PgDeXh0B1Euj3Xyfq626sZe
jW0MMJFHHSW61sSfLrgsW8/W5QPqomwZP7NregqLC1ES9Pi25uz1Tvfsz0I5JFXQ3bWon0T9qUCl
8srd6gTrxaCR/U+el2tdj07WkFBPQdWiF2RAZ1vsnqw5A1udkYywpEmb6rS+mi6DaobXDMHfvWtT
scpnR3ihd53RTAaBMtGcIxdUGHYyyOKYLaYwQp3zGCFXWBp3m4Y+Qot1/aGJIudMgvSfAm1Y2qbN
Wvm7oIWLLMcBvlceFoB/bJS65HTiXO/B5q89ybpxZ0rc0ICjDIumk8uhMV1ebeqn0MI2Iaqd5eUb
6Q7rR+fxyS74V4zegKPqxmsS+nPlOm3IhdEoMhzlzKSWd2xS6knsZ/UlsbIm8IU1cz0OoCW8D7gM
+ZKGGC6d+qfAO89dQphxhym0uRjCiYIU4vc3ZEOIfIs79ZyJ80pjOa2SvX8PKlKM2gtYqx9tv0iH
iCDQCdj2Iw3n6w8ldE+VZGDZiUH+MpvPs/YFzcUaryzzFZedSlAOWtI2N6At3ApW4JrznQn+MXik
hXxl2IMWXBBo8yZSjA6l3vVyaE3t+XlNT/Gf9VsnMCL9MaEFLIAWkeOrEQhlo/eQjqPmBudWRwul
2KNIbcA/jsyBKBttuz0ZL0ZxLKaXAIVC2ueXTZrzyWfsv5j16of7ul3QqNlO34AEiXz7uRfFRElA
pwqnterdN7qLIkV783U2l8XqF6G0sHLq0vLvcC/ohs2UAXRuvib3qYbsXLOk7jeUvSzuu1eJ5CSH
FryUeSWKHNNpzPSEneOLHClVvi9JyZd/YuZES/fCQ79+nVO6Dp/GOp70hACr2MMU6B6F/oWHFEt/
0OBGnUivcECbXkhojTtC8kOJ+kE6FLAOZD1z4PkfHofHZsYhi/x1PTxu+AEbLbNN3GWaDyaGoT9U
1Z1Z+IdvUzWuucsXdZ9+8hPDzX+hFccr0z3lxu6Go/pgbyG497Aakd8vQo5LhcYkglDabAeTvJW5
nB8wMmL7+x9rXGzF2V1TRoumPRcJfBBgj+WCjOAtKMupVcC8xzFhN9taK6H1D8SVCjcuJmeB2otr
Ckjt65iD51c6kRia5aBVSffY4/8c0910Fx16fmnk6vmj5LMxbO60fblBY35LgLCuBQEXsO7oKdEh
XVwe7+OtbbcsylTRZfwIVxdtEDDjSdFvcufVtaWgpNq/oJafhd5qOhdmF3av1FlHykkYZKwa8Rof
keFxN85ceHZeJobzO6nfL6Ta0JFY7hbqAsnPYazMT/uwIcRRrsqmdCXYodXyYj445Ma+aebGTUGD
B5ZrwNcPqKWZLnE8ITih7hH6h3ulmYIU3VozmG8HoEVAhiJg/WJCZJdbZCI7V+Ewhdcq+I3XhEEC
XJ0zWsuAiSulDAvtzxhvZWKJ9kedMPXfTFH/V0S4NwhJyULOEsi4gDB9rGYUcJegJwCPBPA0VI9E
SfbIjkEO9/QdRNDWGBwW9XtrxaWz1w4z2dN4ZXOgjoJX6XeZMhHj3Hooj0YKg1ByH6x0A6s9IZVK
L0Ou277arJlcAXi18opBGVL0CdsDXgex4BFR0rdQEpjjT9P5+uuq0SyV/2RQAa7+DDn8gs6LuM+L
kuUFbgxf8qn9XksX1P+TUGPZX9XxvXvIISqPyBnqsaa6+4XyPzqLIq+xkrgIsdTHmIhaipINZL24
svsBiRkN8nkU6yweO8Dm70VzIsZYw/m8tT+TItCd8+bWBZbtE7stGjIO+mk+uWbuyQdTiPsGZ0R4
01cxrIoomp1ckJp8v990wmmCyh8LYbOTYvmwpwROlFVvz8f2gQItLB74n2ws994TnFZruCgiZ911
GVsutlaEkaJpTrboyu0UaLh7+kNLGjBLCsMBiY8+2/Fo9OBVHT2YzkWj+ZXoliKKF3Wb3m50qf+z
M5LH9W0TOZY2q9BhhDlPQuljruCF8Nm5W4lFuELBo3wsG0By3rrnZ4KU4KwnZDsOgpN2nVRT2ITX
K4NLicFoizV3xQs6U2s5at8E7TS+n9IPMksAmUyfwMPD4/1yIzm1g4RPX1Paz3gdabg4aogmd6Qp
/nPTcuHPHNQtEQ6bGq0mTA7oD2c610u7+lR4SrFXgFXBsxVyMlx2eoRrjQMq5/R8+hvx+q0RUpTm
xzqRJna7S8PAxI0+uZmBldjUybqQLEk/5n86rc88P0PuqdPedsoY8sWldqqcUVdoW5/yuNTWDc3A
5PCBktHNPICiCa6mIURKZZyQSE7AiSKRu3Bu/rDNQvIVNmkXeIutxZie+bm/CUeCgfF63l47A7x6
iRbKTRzCtGS0m4Ol8AI7/Ahccq+r12lR/Z6Ji3+RrJ2zUptlrWP3hRcPs5/Rfuf4fzUC1PDD4ETt
etzuMugXVTVzBbIUh/GhdpDMpuLHQ+f7FDJftUYDMqAEt/pnfu1Muz0jl2yOPjjmWvrdMUbdzCzk
oLYicSVYLgEEFnMc0AfxmSUogl1qdM7HyYNfMfwBPjVtFt6HzyrVP1enhjdcqE2uMS+RXlfiFQk/
oPCis1cbALvTJQ+HWZwCzZdo1Cn3Y9Z1i1z1Ajc8UAjezS8hdInVh8BeBh+YA0I/ZTsUnA6SEYbR
VejRmVXHqqLfW0hTbd1dYFSsWnpZSaCSDKhTKRbw/0JHz/mfjzN9ouOAzivDYxVeoiyijxo03/h8
UNMuBNr4o0UQyygoobTGjsCZg9aE9dM8sBIzlQIrucrAhWUw9/erBcCyKcNlnKhs3kGaCKlr5Ca/
vgQMDovdUIoJRkLM7/+uI/btSWbIzoTLbyWUsa/jyStC7MfPMA8yuKp7uJLJrvuvFwRnFg1EGFSD
SVxW7Sim3w4OxI5BYivEqFeZIBbtXuQmBC0Sf33xUqkXNPbaxC/CDjpVBatK0hL/Up6oz3xdMur1
a0mD72znj0w+uKRu92tQU8W6lpAcn6j1KraqMtcYN9KTWc8nmfoFC5QGzASSZTARUumlX3aCwKLO
iX2t7L35XvZgH577R0RWjI8wi5HOSfz0f7q7LhAxhvIxZ2sEXHSU/7WuBFgjZk6HhBl8X3rT6goV
o4PfywPmNtuE3qx4X7cWA+EVckjpt8v47a0dYZHdXO/znL1RlJTJQv9j2n8vuou/q/klnC3GmC/T
42JZz74ug3rcIGNfAe+KKDcO79vZs9yVlIQNcLhsyXORCIr65aq5fD2TP3jjOX8I4CJCFTP8cOOv
KNCwc5pn5c3Uh1l1nU+Jlm/Jse6FMSHrzaUHMmjgDUH+VewJtmzZxF73Ge9xcVzYJ+iWU/wG4cWz
emN/WKQgRqgbWl1zly8qOT8g+B8/KpD5vPApz9sGsDmsAYyIembVPMSvqRA290G4Zc3DBfaJ1nrm
K8YVEtiJ3XJRsgFvYUGXN7akTAulvCQ5QxYwWDe8MG8sA6bzi3tFBG8vxAmF7vXaTvQDlJJvP1qC
xts3Lj2sKjOpWdHNi5bwSDvhOEbcwCOw2J7Wa5dzFi34oCPSwN+RaMEEyywgM+Qm6Dzk5TQzhlm/
CEYy8dQzJM7jMjX1immxQvpse70VC1hXWIrh5PfECaV96KS/+WZ3oUTleoIjWatebnCtbOo49Z/v
nVopxTrKvqfeqwGUUO36JFphC6ZVxjMDc/yKlY+iejW6ZjQCDinkwYdTGVBW2g8IH4p332/HnnZ5
VRuvlBhvhyYtDS1uoF/LRkMpvfJEGg6ZaKQT3YM1EGaZ06SbJ7yTiiuj7O/LLljM4ydliWUcPOzK
//o03yeuydhNgTQb3viKb+1CEszvedHFvNmhsih8XHDvD9FAh+OsvaWfAf6Xk/lxwmds/5s+RhIB
bysCkVj905PMpsopoAjoFvFVxe2uavfs9nZemBkQtaiFgFgzhUSMRHxIsMIJfxe2utuoTbpzLed9
dy5iHQCtAscaxQqgpZaFhA2/zbk4wDdoYT8CgpAJxL6EOXWLKuU9z480Zqu5OYkIDWnYmGSm2C2s
NG2EvKDxcKOGAHRdMWAUzR/cUlVmMlMj3oEv78k+y9gd11akPHjKQ2UAtm7pbaRBRblvSmaUkcI8
3F7hP6a62XlOUN4KxpnbBE46mpcdwFvtjI+cfsdRLR72ifAycihytiLIleHMduaeAa038qj/Yzt+
Wbw38GZdW3kah1FABq2ga5Egqd3CDGaIYuKt9F7193t/iCUTV06sEbWUzUXHnFyGX5FrKp2+p0Jd
R1JOqt4iRdRtvIyHDtEHWhvcr2kdeUsBUJnX99k8pvwkfQz/Qlg0Q7fqsH/s4434nS++vxn2W0lq
bvSZZiiKZo9WaqZznzommQM22kfRBpl2XZCqV7VlWdXh1XIsHevldUZY9rX3wNVS6BUDJNKjIW/o
ft/nSY0FS5ajkOngZXHKcgj8V0One97kwdPsC54AGe7dLVQ/FcjHXCJ74/QrOLLBX4TJ0PeJ47yr
Zxh8K7Oobu9Dv6AaPdQ2lBd1kjbnXo81vFhnA1j6xw1k82VQaY0fGhc7xihbaWKKO8HDIhp5l9ZV
VZc3SYg2M6dRs/6i3ToOP1JFmqf5XWcv7LgibC5fmFicVSFKuShZEFXzlnFCoMgUwH3RadIBIiA/
6OgKd2mxmKXqse9rE39KIfH1I4dWWL4l6sXXd0VCFCnCfUHYIXkwOjDUH1WDN5zP9srNVEpfA3hX
XPyadcyZtlLJDOY/TeqBmdgjjp3wajWcwwh/Ro9eWZIRKqL35XealSx606/jnWSX0lpmG/9qBwcW
s+q9SfGZyNh5/ZP4dGbucUGo1q0VUzjYcMPl3+loKtSTC2NjD0C2JRirmcRKdqRJTcIzmTcViA9e
ZXWERNvVQOKIB5qW2oX0vHt9puhgYi97oFa9RQxKq0mYiWksYu14MneNmzavKTg8/k6SgrEQ5wWe
Czgde3XdXLznzXqtLriw3H1jFBFzcifG8QZXAC3GFzPudJAg6uLCM/t2YhNypkUZRSaibcHznXjH
kAOA7cBo5mE5vwOskF5dGi7bdoJG3pjtRVR3NkbLLoEvqlfvyJcfrGguShT4BKl/mL1FEoGww7MK
2xsLRA6bMukazDmnmk6SvbMgtiPgOqe9G43oxYsJJ7IUuXXG2R5Qv/UmgmILVsPVSBAv45LrmBx8
eWvHbIUNiRhIT/75b3z165bSpxZcMb11DLzOfp4H+L/wyKPIW0vsCZROk74/kA5qlwP2yTCGj4Td
Yu79t9eKnAkFZfp7FB4troXalv1OytO4OxN4f+ujqH6xXg6bWChEv5g5l9KQ9Yq/RideQKd9np30
7oUaxKx+oWQ5JIjzOrmY8uBR24Ou8aDvaaftYk+ykJwtvAA5Y+vD/Im3Q8s63ry8WHaLa1Z5DYp8
YBeWldcBbOC5wM1NLfSX7gnJKa5RGcMIVphwYc1YIihnuxBLOMKMa66nWvDCsCx2gC+CdphnYT85
DDSfz1msmozf57yHHDmGKOb7FO9qfIKFtEh7efr36kkiVZ1wsaSbui5/NOYHdN49lNi2JMvoyKrV
VMRINQBihPR/yDMd+TqLliE2e1wXWBjx+F2pXMpXH0pdnriRLQYb/gd7+KKl4BNyiychqZasrFK2
JDcM0x2j2mdBhj1UZ6r2XcJ/mF+a03gbWj4/gyDQSaIISkVOfDQ5UABWHh2AuIkAT8cjd4HxZAF7
dRKqAPbVHONo+kdV3G3K8tuosqYt/9HCuuRrk+5JwUIeB6TqIAnVm5pEH3wihBC7MtNXwPMjrnxG
kq1RcofdefQoZSNAHsdub9rNIIZaNS0FQK/dMIS0F2kSEvTt0Hq79obQfDLxlEk0JjqiQt1NjGpi
wOsYAOddBY8Z01qW4HVM3NmRuIgVndzZrao8VZ9BSsVOtcwcpqZ5pTB2BITRFbPXz/loxLVq+fxT
yxJrbGYbPPO4pUn2phJx/68xllqqjrRJ9jsq/QTuQYFX4QCVbOsber3j/ll+IcBh0GRd7R9YQnD8
gRSusebllHZrGjsPBVhp1BPwNx8EKR+xhBxJTBJaY8t84rUHG/235dwhM8VS4GqqzGoUzeLEHBtK
t2cCw00icmHfUFSlLKboE4lU2So9RsngNywD2+Tc9ldlVVJGYFmo4USE5kj1p8GqzZmikHo8sun6
8TRqOKTa8pVoNue38vjrNWREcJHF4YTDacvAAccICQsmGs2Z8G8GCdR1qQp8AFt7RVUeLxiUsAtd
ub5QXPyoMt71PL3O2Gj5kWMUdCFoCXa3qA7I6LG9ytfbcW9RCbetv3gPmEAd6ozbWSGT097ERCOc
VCKK+WP4u5GyPtBOF16NLqo9UfgYSHBuM6BM+URHYLog2EO+IGsjhhDYXuNgUPUnBaq5oSDRZwTI
6hCUVoietijDJgncd/kG4M5vEQs8YTW8K+DJ1I+LVa1WdJb21uWXiakfQ6ZgKvdikanIARpUE5SM
CPL3i2Sw//RyptRZPxjl4aI26rhNm0jPq3iKvR8OVjkn93S/7ZsOyzLidOzqM3PIzmZDN/7tQ1ko
IZ96loVq//HqcKQZZaSr8J5qVsXcPtPqxKft4n+FbecjzMMoVEMErwf0KV9QqPyfXyLqCFTjAkLF
UaV/XGrMyUo/242V+1pEzrqNqKc2z7os3KFtQb38jWagmxzqNiJ0RNY4XvhI1+D5HSHpn0pxdsy0
GU82LCp9Owwm8WcCxAcmURGT8TLcXWWYPKE+HCWFTWY+umZ5bD82ysFeWLvamIfyXtKhS0rJ0ukK
m/YhEVu5Paa2zryAD6K3Z9WJ5BWP6X4LrPHNJh6WCkpJP0qopyhvxv1EU77mpHBrfoJbh1GBOmOu
dzIspr1XYJvsJ9ZGOAfF6lsBIzFGnf8Y82AaFK/azunMiymMhmYnMxrwGz7HkcDsK7T3mUrSYqYy
LxRSwyxST55tPoPwloDqY63HHTsz55F6O6QkHzuzF1NBw/t+/ONeSzcmsLDiqx891u3+SSvSqkhG
poOs3GAd6ZL8Lv3pqhlJuwGLpF9XkS86dVIJIopxrDe42M2edo4jKC8buiXeWaYVRffgN24vuPr6
mfK3QMN+JRxO+MHGeU0qqliqNpNTvk5dZh/VSbqud9jm4L3ThtrSCRoip+F9JvuJKdeIIbMz0x4l
Y4bH3Iy/VYQOHvKcT5NxBZKCNJjjTBnfeSlii79gWy8btWpzEZvaiTh69sCIk2RL+gmDcmbobUhL
Imy27B1aTc2ltdqNHuMh1BuNwi+XDy0YPERWZWf52/QDgyG1WcYjbmNh6uxiHT6P1cGf2hMhUArv
PJwUVVwOfuqYVnYj0FZHIrVdUT4pTODd3tob2lcZFwY/IBy4dkVrPsvKQiqbc6IsZR+snfPovxuz
avQqCtt/FSful/NWHtWa0g8q7N4Xf/k5C52oCmcSCfh83F4acFUXTYHH1R5v+WLE0J2lD4NrS8Z0
ApSRuw/FUoCAEgEMXusryUZmqbVR4LUkW9nbNppZoDbxta41gKpuBntp0MJXtdbvTbYeFz0p2S3p
5QE/tdn8grj5Fr0TqF4IkrgoGYHXneI5pJ43hiJw44+HF7O/9xm9SuUwyLMVZnb73lIamX5Xg8kr
ygtFDGxhhqH653gRiIntiCOnCfIYmgw1aD8+FuSneUKON/Cv+TyvVm/MQq3OGL5sGcmvNHJARr2L
I3V/U3UBou3gWBEpekjZJCNkd6JLGemlzY7Bh8PeXdgDhw9Ry9/cQtfXRG5AggHwG7vfR+JeObhi
fKn53k9N59OI/oaNdMnyfD2ctDntz4kX8lLuPSgj0MOGYxjgNiYRNTZk08DGy5YSqYluUjFzaxt4
cId+8jZfVtokOs4ZPtldKxAM0jI5VtwG/4LHwATjyajKFOI9GGfSB/5GLmlpJjQ2BiNQq1X9Pdou
vrw/cwA9CZE5xEn4WkSMf3lhEEcge5p04OofhoXTs+Gx9bVf+HAg3jh+mlacAZN1cFDdfuWm6sai
E8cHsJ0R9YVrGtocblRd95a9D4nxpssB7SUEjU99uEama1X3fZwLK1Gr79j4SeKqCwAJJRmHJ5FC
UJVe5RQY9Ibst8WA8LlAIT33yPSPY/xBYWjNW6yALpNKPdktqackLZZ/bIShOGhWJY2NoyRJ7OLd
RMlt5s6moAuMYIGH6c2GqM/JwvjiJduecH/hJ+aL2QxP6ZzL+I8whjGJ5ikoIUR7Ifm93uQwsGKW
0DD9xNq39TPIJvRS6CbAzTgE8i6OlK2fmQeIO7sKHhMJqUmO2yz9Q53ev7gp8gBL9fJQy4Hz/K/I
mzvnpZRa09qFqahaNYvT+zoQGaHr5Rqgzz0soChmio8xvpOs4rJ/esg3IxsaM5whT5WGSAze0rhg
B9k381PCRAXKvCOG3dk2TIgKPAS/m99olmE7FpOCsmeQ5pYUHGR0nyKWvV6WSAy2jdv9wuVLHlAv
3XrhZ8N03MyxGpLjw901vluvI0wTkuvMJObKmnb4RsJSSFdcQunTSvDhqzKWuAs3ikYghmlEzll3
8NiZFN0veEig831J9d9hSbRPhi9AYggTr1/4PaL+nwoPFUYCGURGDvmnruTwoFlt6P9R90bD3m3Y
/TP2uVlQPq+RisA5AApencIcAkvF8FIKltoXC8hkGUAkoQZn/jEXK2TlF/qDw+mmC7S3I9i3AdmS
PuAWkwFFvsXjyIbchGgGpeWrRl1uPgt6K44USVBeZMQWkpEvTyh7dFgxJ/X78Sf0qZHCehYg858a
wXXdXWCXWB+iu0lnDaSs2bWZqr2I0KKJMbwSAw/Bb8t/+1GGwoPdWDAWJSpMvwoUG0QKvwzULCx6
2ztnyxzq7NQHBWGtxUs13c2u4frmZjN667yhrMjOYKyGcGRcWonqwS1ht2ETz3gDfV2tshUUuDdr
FRv1UQXigWrodvDuXJUAywTBrfXN1yksiX7Nnzn4Nu6a1MT+qSfLIOqkAdyO93cO+C9KA1g/5V40
2rH6j3VpJp6cEn9W41OVZoN4ak4W58CwDf5H28RCVsi3qk+gYrW26LT7LCpU/4409+onZZiRJ5LA
n6PO2SMtLVZBvSxe9wgm2WiZcyDybtkUzmjHg0T3D8u9Ku1RNgqKkYihJVLq8SboOnnDyUarx73l
p5igUTTfl0I3HNPElmuO3Bt6ETM+Lqt/7EVXRLRfTZ6xrGTiM2/ffuWMF7Njb8112NGlhj1aOfSo
OCJfhMbvS3uOJ3E8u+A/LAf0Gv1QOOU9ON48O9coddfVsZlzvfvpddepykx2zUwBdovh2/G88a4k
M4/jfDxoOgDpRjR8Y2MGytwO6bZnliTzi8x4bY3ZhEmuYXl2B3xuIZ8xduC8ExB41T38LnTbjkGE
cBCrHH3HDGyoptAJ04uyn+P/qjenmt88mgXlxqvjIU4y/87t3YcBFapu4/Od5R1f5KpSth4WE2NU
zVP+1fUC1FMRTcjk04yeXmwgn0qm6WShHoRXvqkCRySHYvcG6ij2E2xBKTXTlc8BFrwwEsyxjYRp
g4atS9dkJk8jt7Vf246YIFTcvwx4CC6TG1qwJVzSJfmNpRVSECRWDiBBKNG4NfBWrnigdXN92skb
jdKRizz9D2fx9HvzgsT+bcYMtqtuEFNkq+egpjwNtQpuhKz+jHa5TnPM8fLVJ7Ri4kJDGvbidwIz
IKm8O9kprhWujbbGjywqHPao+00Y0LTLcRpoGbrelstFrYckbnOOEtSvvLu3pAxXGBl/nZqAVn2l
QdrkhIJQmiEO8Yp35szCWEtW+EPH7nxezLmuiCzo5WQfX6lEPT8pw40W1RUiHmh6YuKmRLIubuKq
ZNb2bbwqnwdrKL8ayyncd21OnzLxJUg5DOIyCDZlMkcoo9nN7T+pdxMsFwW5iR/ezvEstHxPuuzS
vYztrXc1qpvAH6kyZPTLCNoF3ZUqxGpHeZT/BDjVJiwKTSG/u7Z+pg4pcgybRH2jw+GRPBfwCywq
Y+u48pIKfIo/CTsSiUwO8XCQYtVM4Qi+AeSd6m7Jx+VqqKEdiMdRDzOcezkHeOKNLfpSR8ve3EAD
+ml1kEZQhXMrQt2gbHNPZlgZNE2e++969FMIW1mzc/JCVlfsW7Xx7DcmuWla3JExKittxJ3C/VGN
W3CMnRDHY7lmZ90YGxFeDQpyoUswBadpl/SHE5QBJfOVksLwR31D41ZhGWDusX5+NtJw3m438DIb
OM23iawJ6ftWU/8EEk3Aun58VykjsI+jhU6Mqx4n3DdB2sLEtfxpGQAbFHKh9hvtpfpH8fTVNiq2
PENMC3UgKXKZFDc4BZQUOG0UdidYyWtGSaezg084osec4q86+l+5RLdJhTU6E+hogQMQ+FgGG/XP
wHP7gpvKzwEy+lAcwOj3OdZmL5bHYDT/L4DTYo05+ZxTTSz4l4Jj0FME6V1Zu6qWEHn1g5bSUP/H
C5dMElc3usfvf25doVMQwg5XsX9hHuhChIgkesn8P8yL2RbbSVknG3CIFWqD0GDhh89ZnIv32dwH
oKWZi+aVbeNlsCKKkRnYhtT/1aXbxm7koS+iiB4pP0UTkzPfUtynoArvsLzDLu3fX8X6ClVaPwt3
qMpnzdNFFwA+MyCPZaGdpy24y0AkDV0UwAqe+VEB7tnPek7bCqoVF9W0Urf9kLvJRcsSLCWJzjWk
bUqoLBiySdtb51hsZT3CJN9BW5cgLRNhcBL1rfu2VeM1LnvHa9HPkctJGBONBKU+XIlua7jdYZ6p
bRk2ZtbgkJZ8W4ENRrVco4Nlk/Vnu8YB7WLvrVHm+RJ+fL2ak3UXhxJ4hzJYWjm2wDdB2nLkQbsW
KXrscGkNcMRUzxfcgpWr0z3ByjLTUET7+1TnWJtEUYt4JRmWHM23mx1kZSQfGijFGfGoe30QFYq8
rp4/mFW55nDvK4CTSKdu4Z3oSAbOcYe6vR68WCJtvBbLkQ//r8h/hi4Luf6PWka+7tOQ9pBJMDfi
9NwydNrV7x/3oU35HUHqDoFIwnniBLwh+QrWG+tkvyQy1TbcSAvjiQHQYQpJxZ6CoB0hFIOqhuh1
PetjkBFUuO8HnQbbhzMvrR2zF0Ki7bl3MyK6gJLyv49Di7DQmS9iOh44OgHb9FxJIeQwbOEf5hSJ
1KlQN2EWIfBe+UXgK6k18EBy+kn+1SU2EKacntCgRRDKzKZHb29qhrIF09EwH9sRkI5UYiwmsFPe
9MFQnTQFqcG+tUiGRrewC6Msugw8L9Q/DEWbRtzjZu8D2LdoE060jB0UaNw7ueJBz6SER02MDopm
b2lYQ4AP1YdF/SYlh18MChlEp/EH1R9K3p4XoCSw8VFNYHuP4HyBq4a3w9jeyWnJzmOZMPWVacfG
9YyXiyxsjevBnwjEwMe8ivQaJyJK6T8ixMDZ10KESu9ZKgsGw0yxnYMQuZFqCdGl+vYJAQEMYehR
2BFN5/+Me9kW8pffu3ynkbLKiPwfcm3W48ZNboQ4vGLDfLttEui1g2r7Xvif7FmKK0852DF06rXd
LS8BjSNOf6nJevtogB2RNbarW5jpD2/hUX855qpzLZLcPxSMOng0Lm06L7HlObw5UzCm2ngvjqhJ
VaDinp65AQgIlrW5C5tTFMEleHq1GUNacD1KLn62ZPIl827EJ73DFrwwseWiWuiLhphP6hj3uEU2
RKEatLIV+PCsZR7RoLUWRSy9os4SJS4YfEdiRNneA4+8DJWTbG9135inspdRzdZn5XQ9fDwAPrwK
fQY+BGkL8r1ldBmVkh//yIDneJ1jvdj56Hege6ZgghlLozuwUm56Tg3lmNdOyyN6C8j444V8Unkm
UPhmuj1ZOjYTKw0YfQRGUh8E2ygPlx4LO3enL+fBaphYfBjL3saLadVaOqS0Ub8CRtpZW8eEl597
eI/vd7WBJlLztShmhK4l2Clj+mKXK7SZ4cVZF1ZvKLFKJsuoYCTy/pRsnG/NPhOmy0vRMx8WPvEp
kZ4BydjELA+TCnbKjQMyISA9XnYMZY+MXwN6bm/m/Lpfoybf4iUZI9N7x6ATZFIS4UhOGfIafATx
WlCGSA3b8U52sR64nkANy4MoRNKb6NFa4qPHNv7xttwTtw8T7xU9/Vum1828Ryb5Kmo3F20qa45H
YLdEbFFkZL8aRXtFNiNBy6YDOsuzbgXZTU4CR59m4jlq3shSUz1AWs5advYfsU7aom9kt27tpjJE
NKXsdqyTeH3EXIDNlzfmS3OZn4Lv/uEnQKRjXugfpUxeis4pwUc+SZBpIdhZhhZMO+3Kt0ouFmVY
p6pxgi5o5vKF6kxUjobAiK51koa3GgJ0IWMgde01Ike715O4zjA5dtBdmTWHE7CgVD40+XjkymuX
GHRCZCHLKSdzoAdWLxt/vtci9kaPOTJYu3UHbfLrabuP3qGVykkUFHIEqc8OdxaV7KpUl1+XUNm9
JHoucZvCoG4U+hrKblwtXlE/cTpg11is0IAmdG7MZLMTkFLHNuCGlx8GCVU5D3ORcYT1srF8sFYe
/hy1Rb3cBGXOCmARQwTYpS3alhg1ght6qGOm7dlgEO3NDYTfB1K7VY2sQz41rIbREW5gb0sPQ8pz
cy1jaNVSDVMkAAgUuY5HlIXYmXy7oHbMOypsj0dt8zj48dtt84EM4/f7/vIMGTvsGI78xD5rVBbv
YumNDmWEVRogLvs1BnAt0xEikCbjpihiwU5Tbe2UT2NEZEbqKuhwcOTjCdnjY41LxpUmd/pM1vq7
Q0wcHfBYDxJGRwy1j4zzW9E2yfd2AtWBLvnPjv2RFmdKyGeiq2rQK2suE3S/WbOion3H/+UL6jPN
6pEsA4hez5bIVPmmuzqHIiLeH7rSvfTh+zMH752RQOpFCWluhzLyOPNjtnZXJiQbOrkmV6pQm7mx
9YB6g0AbUQk8Dhf1KROR9hcWXjtjn5kJJnPLG1jFDGVT4tbkaWnYp9ryAssiqk5yy77pbO1QmoPH
gBVpHZmL/oQ72HcoJselPwSmO45XIZcXKDGEQrjiQ1Fw3m/m+pxBC1UZS7HxKE0+yHyUQ+JeDTMl
T982kf07t08mMdkTiNDk1Ca6IhkmFx7LygH1298f+bRWTXoL4CjzdFLVgiD8dMZ32ptwAV4aHwP9
k9y3Hb4dHo/u0W8RTM/WMWHr2T8zA+kB9my4xwuhmaghz8+EMOyQp7peX8vx4zubEgQ/zRm2snzx
tCDR9qAcNeorePJr5x839GQxsVGqM3wnurDvlhOH6wvvH2SLiigdrLDDj2l6kvq8NizUlpTWCcuL
df7Ki+jqPbBsKsjSH5QZVAfGj4NBcya5NmebpPw4bjQtDmjN3ZclQAdejtE6c+ZoR3ifM1V91L7z
PWKZZUy2dsUri/k45YW8P5iyY//uw6S64n5XrhKIhVLY+i845UzRoM3iBbfV6r0yxTZ0AXnQBc7N
M5SjOFhg0HWLpggCkt8KPuzLMWUA8MnQEktvo+g8VrT0bhapAgIUT4VO1Hid2jtcWR0GhTawWCnV
kNdSmg+gTB63UMtmV1j+pYQcRssuz40ajrPyGK5dp47G6wBsT/XVDEgR1g98OMJ0JXlOlXVnwfij
q9/jiD4uIaweaKvzb2QOzSNRZMn84oQf/hKu6BgfHwaL1DPRKkdbpbelZc4A/ymUt+oaGmndBvxI
Cxzx63Wt+a2ersGso31eFpUoP686BhDx0SpNU+tVnIKoxq2GhDfbF/3MdKQvrY1ge0lCdJdl2qoM
CN1um2EWJR0g6ssHZbvdLXzbgu5Bto5nQb5ErVuh+sH6ySz/bz7z2O16NWZlV+/2g4ZItCwtrUCG
VkxkPTCFRyrok/a8FghFdQmhhuE0hUJ5f3wmpflL5YIbgTDq99yPZMMpSnHACG2dQpGhyLF/8QCp
KKisxPmrntq/CZEs8+LGD4yV0wWxf0ZA5XwsuBq+FbvgdDPG+ap3fr++OpTpUvG7+KxyVifoISC2
k9x4XNLp6a+ps00LoOAofZAmOFG+WNujhCs85Mz58SdW+HFe/4ZXbqKxWSE4U+ePBVmIMN4FNKJr
RTNDUnp/Idm0MX2ZtbkZnlUlIUpqbLVHUhlPX1VWC2wHqU7Zi/QDGaukocXM+y3kuvpdIs6befU/
7OcaMlgoup5VS0q3vAXbqnjCreRCwdgq77OBy4sbSgh0jPYMnUPynJplmR00LKL4xpp6Un6/Z7px
FwsUJYxRoxgsU5EsJ+aoRaqW9zpylbKg58rwWdCQLEOREN8VNKrbKPb7Xe1yEArqSltB+N3kr29j
wh6ttdIkRHfjGT9Mh3QwTY9w80YhJUYmdq/d4GXqzQo9Jj4Hb00DVEpLtIW4bQ92utoxwRSkRNzO
/2aeYbl3DI/aWXqcagFd59pVPEeNMxwNMPx1VyJspbRCdRvTPGHwTWHTdl23txd6NYL4LOV1PXYo
fusxO5y1Mpm10gGLG+Wd/1DLlx+Ay1zk42lDTnAI5mmnn3xtzloQSs/CWAWlnuG2klKnvkoQ+f+p
e4KRViiUYuRMd9RZc6LUaBwxJ8YUUy+5DpQnIjYXhxE5MeD/v/2qua7Wxp4QeCH2Jz9kJa4kHMPN
F+ExdBS+hseagnEfgLRU/LPlTetkiYRQ/Pw+bMT9r5VPLQE5jnhGxjt91SdSomFRJ3oc4JIyrHRK
VwCHTsynOOOah6V70rohsMEcYm7Z1D5l1XnK2FftSxYc0ka9eBKVKPc8wtn/hgzC6G0Ho/7uDizN
kwUgiwUFGU3D3QgcDU6RX+n1KEo0UfWU6qFfu6F+v5n/JKMLu+xW2eOaEcx4pTvCB9Ox/8jfROhe
TelYuCireQQLHfCiKNXqxv/EvbMTnfO1kD1A3e9lDY26eOqYcmtO3RUgQWnHtTfpQgW6pPhlOYBR
u70rhZDXQMvUD79fgwcgXQ1K6Etz6P11Obrk4h3yTBhYSP5+x7eNHidg3Hq8Grq5rp7v7TVElm3o
TC424eMHk0Ng8Grzh5+EO/uh3PztzuVtcWXkn1zAZDw7KkS7ICelwURQGPPBCNZc+AQMYw9O6HOP
tBPM63BhOSp6S9cY18qu2OTx8LFvna7HdqkOgNHv9sW4NSIRh8WLdaccrjM7mz8AlWPrYkEYaEvH
xuzwj1FFqe91wsI7YGb0IMShQFs9elEznRG+S87Qm/+j5CcFldi4v9lBvVKrYpHl7cTs+pik1pb4
GN7r1aMtwbJa9cyXBQN0x1pAz0BBFM8Gcj35y9Z3GaP30Q2BXDDLaS8NFMHqb1ouXwU3M51bSX9Q
QC+1UjczHdnyxqJKw9911OzP6dI3lxAcC89u0jJtlk4bffcy+lr/t2UUI2nxae33sAG5jamc9mv7
xPd2t575kTblt2ZgfuULkWjv76d1FGHTHb1Phq/Dv+23OmGtw5sAHYKQYZIbioDI5gCt4RFTCJHR
fTfhb84X5DmW9qHPgbllCIY4rCaEd9bY5Ei9NR+C4TUjqiSQoDCe6/0EOJoKEoic+ycF59rahbZF
BcLuUvbmwUrACOlHv8dScWByqJsC2zheMkzYtjbg7Xu4amEtdXbseoSSJR5OzZ+fxmxsEm6jztXu
NjultTxIv3lVgry9fW2u4G75XKXb4e8L8/123xqD2tMHNBSXfvHwyxainNtQWppNH/UpitjSq1Di
gLoKWuY3Mfu1fC/73sII3ScZtsNp4Fiw7CbMRS4LwdU8qSG3XnJjupjG6EY5y7WMUOFdnNJPQqd9
re15ySB5ZguUjEB+9DEW2aRz8rlp1HuJNfm8M8m2ol7A8+q5fg36EpvWzQsn8lD4gbmnIgfdlzEx
uT5zMU++41VPyhlI8aa3BDIsX1aQuI/jSW1yg2heJka79ElDuEtnFMmtpnsuhIkyTFXaFPFVvn1U
hEq0fF60H0FXcnpImohOyS5jp9UvuZtlMBAxTzfQ3jQK7hWeDlV3GgTjQWCmxtvKm/taxGVxXjxW
hQGJKk6rG9GKqPRlRP0CrtI8r4R1eck4LlFJd4XPkAzn+Bq8gpXLXuEffQ7yvwMXgboOHK4XcVPr
+2w78lDscf7ZW6ZpbrVJcbSD8Kl3H1AQ+8dIQKJ4bbf+HZEnK5KE6hFvis98GcI+jQnkmZVZFkBn
8r762+fUSpQmB/ZMTD4xuKJJe7Gl8IY4DjuWvk6WWXmNQwJVmo6i88UiTw2YVIkJNFEoUqAU7zUi
QSaSRWNyQSQmcFIxsdfuDvFEkRwjJaXQpgrE6O0O9kD+1QRxkCT9P7DaSkC+p5MR8y3eNq43o1IZ
sox+cI39mdKjA71P+SJtAyja3fCggQnb/IE6PvGXDDg45zv81lHSxu/vPdZ9AZGq3gGuhOw77weA
Lui7ZPqoOeRDNRVnwzH8xOxme0YFVEr5WCtexjv/skgVDq3fHNCP3ZrId/+TS18Epa99ZLwbGttl
YhmFNdcKoymLO7aoakOhMTGZzGe8JlGeUu/UBAtGOuckEfc/0ZkXdHW9dUpzm2VCWeC9+ghE86Dl
/4wyowL0t1szErZf5nEhkP0f+tS0zqV3TaZ1VrFZhaoHL8JO33JyUWMT5/MDlIP6r2bAhNO7RcIt
oPeQIhKkd7o8ctBavfDqbW8tZCW8bln8c1n8cll7t2LKp+bo/zgwqmVJZPtNAHlL1wmI14YUhxLL
95mTkFccn59oiVQt1RNSMut/P/A5D7AZU67UmL5HMLVpseremIpQiVs51KeagsO1n5uVoFb43izV
6vZN+s5kafLQ5y6sUZqx1fnF8iIULx94M5k57sjsI+A1MxGhOOEMmZIbeDilhCpxEI+sqcQ3mMCU
z7++ygpbRn57ziGCyeyeXmMbSlNDucY6bW8mYqPZSiWnjtJkQ99ptZlO3uKT4Vf/xO3ZSxyCy8PS
dSDq7W845AHupMUEK6ks8o0eFO9yeMaN8GvNCtJhma5FH1Y5WZAlzK56Tn1yDa9wjILLKdG4wae/
niKbgsReWI0gkH1kkyB8rLgBme5EKRpZgyR8hH6aEDdMR4luZRxF3i5sUpSQ5BNV8KCl4jKE/UIe
ctzRu1nc1j4uPQJQAvS6a/AVxs4ZT4SMFymr+m3+ASJgrWNnFuZoue2ykAxZ3o8nuUoIUqHVlkTA
zTOoKcf3LPZMNPGT4R/qUjqFUEXqtG4fsiniFib5QfyHLL9xkO85mbT+ge3mU++FNOhuxX0oyhMv
YJNPR88qG9W3hqjS5iitFgzt5Yp64zlkP+moutgtP/XsZTGwBR1O4Jtdgo71sr6swt3op2rDkKX3
EMiZqsK4kifhrsqQVNtY8DrgRK03XYK6WpJjzOs5ldi82f3dXv/pmOVLXj8+5DKKt13yxFIuJfsz
5U0IKK9TwGx7VK6JxPuHqe7E0IX2qNIuciyPq29zLkBtitsauMk0H39uadbfbP4TiOnfkhy55Onp
B9IEr5RZOyCE/Q+4KlHPy45fjYEVWg89v+htIS4g7+bOv4jCRPNlSF42FXkFgM9y+eQF/rNjjRyD
xuPlQIjwFXw4YmwG2PPKkMc6rYC1kHJvYWN26Q84KUlaXnD/sLyjWhXJoaqSbn/6kXfnQpJ6p0Zo
BiasOu5vw3zHSkafM1D3cRUFymJO+Oz6EmRwScFCh0fgAO9yWM0V4/wc7pWusobKzBJ7ueDkQUsO
NXVKx+LYQEkrR0zdvUOdBgpi5d0/oFgIGOCr/I82twBcvxjibytesINgT4eaytny2Wqt+3PPOn3U
QSciwYhu92TZZMRVyN8NiBtNHLX1hQ5odEutMcOdRjPHH5dPkgslNZc0IBma6Ch88VWp9XzFLwm2
U6kOj2gxhxav92VRs167HAMT/yTqWa+9lo/e+4xjm/UAqpr2xftgLjTgDi/fa3EhEu51s3OM05Wc
G3CSQfqvzSTadNLTIwIKQdQZ2Z3WSGENLy8o2tQWeXnQDj5x36USTYZHdUO8+1yfj0rpV9GhwWKD
pJDoU4Q+BVfMhu1DTrGdSzyifvZYnPX25VsHJNSrJasXQd3CvFSevMtGMt/7SxLjCHy0ztNCJA9n
hAdHJQIftpzDtnjkmfzcrCC51PYA0m17vVB89Fw35LE4qpnFDtpEPUiW7pEXlC/Pru0R/CpvUxiE
ttAeUhIorEnE0V+85lgshWXNbPcrYUq2bQ3MHr412VLMfh+OiHTJJ4v/g1nj5CiJCz/3qsZw9HrV
fQi/oOFeEeVICqP3JHHP06vhCqEW4NK86+YxjDflJS0rNqFFHhXQNzF96BbA7bgy3zT5BlgJrbJM
wJ5idTmpz1wZ/mKux2eqpxkl54ajUSiSwnu4J3n4JRpGIEQ1mBqMuGD+fnCNYZzhihcBMSxWOMe9
uSksU1WBz6YSSNH9sZDuX8HUcyReuhTR3G9cTjUWl2dNWeTygpp9XVe592fB4wKXijZivXKDQ6q1
SZsFrxIqVwF0ZVxEev0ArXMU4zZdXL1NoaZBK90YVes7NzVHhF3h8bgDB5+QGmkBW3pvW9iNle3q
lIH3TE/XRR1ArqyenuO1xefIau3s/m8sBvBkP989SSlHs0HpYFlfqciLPN1s8QgHK0bQ6nHylCNQ
BhnGxclu1tbArCy8Tdr3pyZlRrv6nnjFiT9c2WckgCxRHgYzl3+vXW4TZ87o1234D7Oe+x7kpcqt
mSseaomiSrq9sK9RGvFe/Re7KDfKRuKo3dwLWal4H3XXQ4eqMz+4hE/DRf1m+hCuzudKT9Ujwskk
MAyU1cqr6/4DBIs5QfhSuQIAd+m9afCsiYwS3Dvat41HIoH71pO/3jm1JU324MIKsn48qehyWJv/
mjNpGbNmVSPwsphvv0Tj/mjkxhD8+QZTL1OtwniPBl9oKQagKT8fb/BEzUmj4gsBlJBxcn67SACI
UYegs2bw1aQYiUvw4nRxugJk+sZRBcIwPmA2V9YtT5qdI0CgF9JApw4HoE2Gi6IKgTpzKGemmE5b
KKP1/bxnbfJJW6mIBsszd33ldcew9U3zx9BG1cqRD24TsE4bJtr9pdGJ8UF8yMvOjHTuwP8MD9uC
QzTX+/saar/gG0ySkPs1EDej4Aw41kKjURq+m1zWSwPhqi9kmEPv+DAfOdftTXGAeZFQqQK9kKvp
hXkyQYt61X8DwlcO7FreUGmQtD6cK4uzT2Vlu/4oKrCQjXCUm9hbQl144Opt6feNFMOXdnuodpOQ
Q7aJK3x2DS0FUq07oP6csqxe8uKopI8kgH62w5QeH2wyPi8wi6aLPRcLrfUAwr7jWFiYYVytx5Z7
pbCuIg8q/fcN6IjZrQPnx/v+NUxWAadkbKqoWZRLP4eUJEX6oEGywHTQ9TYjaGKmSHst8yFA9UDZ
duAhxYSrbf8qWSZ96C0xckPTh6cW9LQhPSdQrT1wOJ+JLTrTCZQSHlCbAKcqm7XMuUscMEqBdSBV
D2KeO2EXd+1Uvm1jbU54Sp1u3GF0U0XD2F670O0sTTe0nDS/tV9AKFSH+gCn0bwXS+573zUHxAja
edYIrKHX2lWs7vnfEvL9W5Y9j6RO6y6SJvpCP19tnnu/vxs1/QUGu9QuoZMu8242mDo8HOOOJEiT
AQ5993rfRd5NJRfB6vi3NOjF++vQVhxy++2FKZi+/MULnWH1ZcvCUi/9drUTjqJ8GHTDoEvVwYlN
k6fb4UPhjqTwolwssxf8FDkCXdoFslVD+Z8VA68cypNaqQQNOWAAYUTDkoW73pyHGyLr60dHYwm8
3rrVgKGpXNNmkQcw2A7464C58Nn4KXCBqOHQ/17KRmj0WLyGm6v2vPtX4+B7qNqBaGR+4LxBZKBm
IvCeBGpIFavN+PvEoyY0OLO5/lpetcWscGt5SmUqF/C9Yg4LaRl/PDWRa9Xt2VtuJM+VdDEZV/Fw
M3Vg+pEkCkheCHfTthANBhaKrHiM61Gn62ujNyXOONaiX0K2fcqL7kTXkGWlO/ERbKbvWF4Qtpaz
G/4gZ+KE+yO9YyAM+vwvzeskrXkD2InC879UTl0iUeccFTgQQhfUNN8S/FxhRDRfwg4g3B8Jg+J5
9f1gnw1nuuWBVwP2AJI8CP4uLRYQFpBcT7Yk5k3BepKSV8eTrGXR10yeTTjU7Myesq2JiIEkcfiG
BqKdlkQ0LTP1x5P8kimjoOj4/ghQAW16Iq4djRu0ly37hMtyFWQ7a5yZSJYMknbSfQP0+VbPHrAC
0ToMFMT23S1ItHZDKk7XwKM6vkNalbjmetXR8i6rTZOyx/l0xP8PnH3E0IuP8fpAb5YJiJpE6SFI
xegA8iEsTbn8yc0VFr6nJij9hxkODnwYlBE+wtkd1R5CcNDUFN5ladgAV/TAshmQWzJkNXwDx4JL
WQ/VkQF3EX8TZOiyazrP2SNDNNeMw1BdxLdhD3cRrq+UdhTtSzkSzZxhSOu2E6cIUDNoFdCWbiGp
nCzZK4ld4MOIOsUkbOltKsmC5HxI8WvESBg2JWHGW4KJVMqd5V/JSGV9NwiIMW37hBy1hrV4N0UZ
LEf4wWnwIZMy/ho/i6466P4vlor6bh5q+Z/vnwjS6Jj2RlTmfGRoD8uNopGPdNEGg3dzfrergiJg
Kwi2tiW1JkG4DR7UqR3I4yD6mrqxeVgxI2cM2hLvfv1xalR0FwzfIIW6ixyb832qai+CanwAYYs2
kLXdK6bs9l/8LV5bHFetaTxQBNqYeQm9+pKAViHUpRedRSCuZMzviQYLLvj+2/QhA7IG/7Ntwv4l
GnJuBzPKC57qysLDpM99PIC5nlG3PYuzrpY+5p3hZlqRSZu381aJgSveGEwjxWk7W2pgSh1bS9Ok
s3sJ86qG2nyvkhrcX8sduq1Gq22NRDCNC7qnLl0ussFXy6NQ6RLdqsrtfisSj0ekHjxMxKx5Byja
8lKC174uJk3cdfU32w4ykMT8+VB05MsMGCrDtFtJRUojM1esCuhl7z4yYYkcrY9Km8MjFpFjqIaq
y4M4d94+twToDfjO/ipnhVet8+fwyCHgfTEUlz3U+okTN8foPm8UmtomnYj305ghmvvDU8PmAqsa
yCre5jjJRlazSMG/YdyH9c7FwktvazZDqIy74+k2AvlN0+vfMgovRHwrTOegG0NMB3UVrqWYoPQ9
bL5z7R+Of6BJrztOWi/Q6v8t9lGAIIOP9iZrLipvnxhbNwVyutHYQf66muV6NI5O4w0Q9ayasA5o
YONTiTL8aC+l58o9GyjLQgfpcAV2/3zA5CUdEcVHn7sDs8yJRuGYzgDc/vKtB7Q/yvchkQiLWuS1
SpDbaSgHlNqeg8Ir5Kht3cny/ppNQSeq8P6S3RJl0tryR4lW8aqkU7m9rD+mtWV7GGmSPQr2cyrW
sim9VouzXsAI1T2aVA8uwNZtQn1l30nei/+8j4fNhsEcIkpFqC61/dVUiH4zSiRxmSZGbVvX3Y2M
nHGvK5kQ9hv75KmlZ+TRSi1W6Yif0AZtPFaJzpGfu0DT4LyrMR/XdNR98ZYNgvygctAV1obOIHsj
tIUorv/4XIjt3FdNw1dNu5gk4UwQkqsszMLAB3LzBd2UoelA26uu7lAnltmMuBOgaE4jkjIrFuHW
V2r61qdsm5HsZOXw8snOPGDShIJaL8uK1rVFLya7w3dCD1b994+4xcW8Apu5ILI4jsXE495SAo4m
laz8GVJF3ZBwEb8rwMZXqQHBUyFm7wpcsmhGKAN2XdVKXBZ4t2kfIthECL17Qj5+BKk9rW4608Kk
jkoPbF3HWTRMP31fy0sxYPZaMP4ZLPmDwY0GcezzF1dZfjbkgF3Es0chTT0BIZNpPb2iVevi7ao/
p/ll7s4yZ2WfDEIIygajlEYuS3hjFyv9/2smOa3JaWcz3KeZYtl1E+2mZ/3zP1xzLUTKQAKym/+J
OIvirTCdjWxTDmc96sHVN9VO2pE+IZGtWywoAmzXUaKLRG0Q5lBI5ToHHUr5PNnC9w8b6YOumqO6
f3G9VBYN6+blXAW45dM5yKQ/+spWnggBpboGsXXSX8WiwO8rvEuz/k1jZFkj8I0doC7w0hqrJNvD
f7tp6KlZ9KCW1o2ZECUQG/6Qwdv2LyGkSHWGOW1SbtWK03aX2V9nc68J7WFVpUJdRolBEwvCD+kh
3H1q6LRSeiCUwsoHVoAMNCCq0On8fsGDmNgBRx+KqlOicbJxTMI2zMOtEXRsiiFSL1ICp7U9TVmd
ui8cx1yRi/8Ym53sD6Z04T6jM83padRRtVXQbEwUujLGZduU903NHac2k4PRUeXPckDD5C88co4M
/MBDKaGy+MpiuQArobecB4o1mNcgz+lKOf5MEtUkVPMAQf78BK6mQjsNBB58fs7P8F64aeU2t+5x
KtnI05dCBV3R5ZbwTPiwURE16HbOqoikWnJYieJaiBHJtSVpP43TfMUyz3TcJQkeCg98Nz6ZbhYF
prJZ5CE8lkrHcKL4NnPmltzKb0EmOnWDtRMr9zuzTOCEXzntwHKOc2x4sjc1Y2LHXBnqYUjsc4q8
/oG9p6GVV3lGcD1SVu2UvALIw+i6Wl2kPw9QNXvZqsxqPxYPUdT3aiBmievNxbeM6GjenyYq6ZH/
oGrqRnSNW4Ch8ZnRmNmmZJXBuIwsrWX+8eC+iSXbLDa+oZbpwIU4N6UP96ES6edYxVCN3qqKZv19
lW5FwN711bCaX3N8zmZ+eBjW7EWmP39traRC/r4gdW1eDYQS1zHbeElYahOtAzNltrR9DlBwBxYH
5q+RlHia1jc97Epbyth1U1ee2z2KzeNCCvKzovqDONpVy1daF34yTkKJXWH+8iEQsfhTMR/58oPS
kn/jrVe3y1RhZy6y7Nrg9iHTvx423YhgJ0tAaBarWhlLolIRu1/kTbRmmOZr8QaWDBHtb5aTEoA0
m5G2FKRXke582memOWEWbWyLLbE24pwM/U3yPkXUpN2SqPTUFukfm7cOYjGhlhsJhz5lAj65NzRX
f1L11AQkJGNMD5QwlMIrbbZHTGMbNBJIozf+N5J8Y1cDk/2ZhuSXsZPFEzwuVsGstJNC35KUOk/1
NR26cB24oVYsE0qUm0eo/dcFrJ0Bg/uCD2bNJXQDLdnqLBrCvbCtN4JahAsI4r8SRFsv+Y8/Z0GS
AdT/2IJJxCV5WmPtF9RvOfmYz7xnMSiiokDUssDxHQpuvkez7lAKmmHck1B84g9zFtmkeYxufUbk
y/q/LbESkCZTVaHAhasGZVBfgw7VfTGX8LExIyeDbjXfZNLIQRl22BCUTA+KK510FXX29cZtMB5N
3MlfuAK1EDuW22kW63zyhAWkBUbN2Z5YBm8fS1oMLUm6NOzh6bTxKLjzbfsRAdKzOYFyiFJzPorI
lRBvh7QBohoGy7AixNyJ+3S7+xmK1C/64yRK2+ycqrARY6t/v4HXzEFFyurK/lRDaz+DpzmPAYUM
QWnH6IhTa3RsLYh1qnnrFU5fzlqq7YlkAFoz4NA8OR+PimvG0z5NzFYv+K+m3UlNAGbFSo1+ufhT
HJFAYX7X8JR1qAv69d0wwrq3QJNUSsBYt09SEn1g7cFeWXA6oidfvrM7eyGh1R62bqDnzrclOV0W
QyBr9CCExO0P/yJaunAz5slZMMqFhyWOE0Hw1FGQoVf2hKhJgzEglnpbbxh4BIeoZdYZAn2U05AA
b1FeybAkJZOpAdm1sebJVKHmC/w61yytGbrip1nKs/4c0Ig/xoqLi071jEVxp/u9z5yGzV+T8hiJ
LF/RJ65rmT8C6RyFSZALk4JgJZycUBRUncemDKK+6m40KBF0JHloI1Scr1I8fZ5IEZQ/G+5YVjQw
+q8r8c56Ra8TywHA+/sK5j/eNjClPn79xUZ0GsA6/nb7/t2Ursblip1bk2YehEW/xD0rz3t3aSZe
YCIM5bxYZaJsIibvK55+pOSP4wdKl8PAKsCcl8UU4Hs5VpCYGLXSZ7P5VeUGlIdaNoVDxRgvLTR4
6BsQfbIu+uStqqZRHzPbMhn0kiUFa4Xg40ESZgWN6cQTFYBLs9UNGTzhnVrhFsyoIaHcK/MTvC9S
ktVAz+RgmJwOgzKSgsBo0RVFaHvrz9+s49XXT+t6+hdrz9OT0/Hzcskg9QBg491k4OvzxwAmNt0n
4rKTQ61dR4/oeFLbzYMGDeJ8gTemv6mmOQcVIeKCksNn4gVnhUY4mFMIGbarpW7ewrIzqkjkXJ9A
0VgfwjcZzNsoj3fHBS6XbkKd9c9856CnIndADon27i1r/ou/ns2dYzFlZZSaNtHLF4pm+U7EJCnh
IQK+8i3mnYM5DToyrdjT/QnIAm7AXuwYgGRq+NMNU0sToEk9DJVQrhA11c+Xq0IfyRY0cNfEbrcS
3v57Y+MENg3g2csl9obH5MbYtvOepuLD6uFqF03BuvxitQ2/h8kyXC3ESduqFyPBmNzNiIN/VJMM
RrzaC3mi228gTjLjyzXGm6DcGTW0lsPoz8Ms2Vvzm//TuGvmdWrO0+EbajdZaJ+KE60gLOHB5lJc
m7eSiudIXkhE2xU6h4ENclvuV+/T1sp9g5xcPvv0uvGsxfF8U/ednMv4s9USqMV/yfbJjtzEcmVE
uCWquxIw2A/faJBRNE0d/RhhY4A50dDRyCXIvnHiJrC4yUdpxAXX6l33WzV1bv15n/zP/8qXwNqb
PY8GaM0dGbOStwG9W7eUSzkG6p7ixI9AE41XY7qd6MUGMQiycTqKEjN8Gmkhvdv399Ew8rRyNHxt
kQfx/7vNTQ/goE4qdoBGJUh8NdgjixLSaE8y371L3BoCLcdJmVrj63x9YIO9BNCOfg0auuJG4LBm
uE8uzaBBQtQ01zUQc0Z6B4MrR0jrzZ5QR0owY21/A13D0x27kw9iUPlDY0z7xBR5nZOQwNt6FR91
fIo5XbrrQVtrKQ88sjBY8wKNZ5Kk2woqfgRppWXyswnjO7LpHdeOv0/c+qvBIQgiv3iz3eisg1Tl
J2W2gpaGPAWSRTbXQrhzSuYofF1u11y2blALEcc53jA7Awn2FIkh0MGU+xix3TtBBuvYL1+2JCvI
1NzvG9sObuszXDzwKcTk8k8/pu/C5zymtrZsvyRVOlHBN+2daG+t+vfvdNjc71xnD+Vny8swt/iz
wXptRiinif048plUTM0xTQsKHhWleNSLj51i8zTBp+YauQG3nMU7ow4JaSLOrfTaMgT17a+phyjl
8WN6OvVIqKXvcRJt5gCWFpyB/FwcQorDw4RvVVNewFg7rzxC3OTZifLC5z+fsTCCHgxp/7fovTAf
k+B9fd/nQd6NHX2MkVQvZ/YEh1mSRTWCEpbZArG3kwVFBRfufN9v54YZEh6fTPFlktkImLHr/Vh1
hcgmGMeNgUEuRpju4l2Wlh2sx0ytKz3o4pAzvvOiZAndEsbTOFQDXKM4OC7trnMzh4HvAkyria5o
IzyZA6rvn2wq4hNHIlCI9cG6fPAlioR2Y99EULAZs+lwhCJ47Zqgw/YWXqhEUXzgwjrv+WgbSR2a
wUkHZPMVWW9F2cBtmgkEZAGLNOg06z9h+dNBcQTONywprxEnJ0FyQQGPp4ttTJqMCHV4SM7PAz1F
NLEOhwBQU22l86MYniZfDzMGcFGbCfCe1znmkRj/NhrWD+DRgEg9GyOmRlk8gEe3DNOLtcqCdD05
nDPRJx7fLtW1zDLWDNzhj6pA8NYVcDLkIXy9El203SU+2xAqLXPV4QN9xE6eZEtKUrZ7pD8v17Vk
RNqph49/dit495g8SDD8NN/Lo8bETvgyAGciuDMEoFdlwMJCGqjcsbKeI5LzhyBoJcE9oLTO99A+
iigvPogG6x1Ufq+M3vrMSTGWReCFdetogogFd/vdL8MSCJLhvQjjYieEdxPiOHJK/9aBgB41ucyP
J12v03MPdzTJ9A5XwvPwSEktCTED8E99zmtPcsF6eM8xiHZjV1lOAGmb1n/jznjic+D/chCy1v2R
mNbaYFqT+i0dBD/Sih7t7MVqxwRvbsQOrm5b8coDuOnz2zaMdH1INT75xvxEWhssdqg4PJ047T4r
zvRaYdyPiwvr32Y5AifpjTXUY9niLi6mpA0ZimBGIJ8D07wnHkAi5sMTMAzd6FNSJk+c9gxIShgX
7eRHEYPci2+D+I894+wH/w/M4a3ZO8j5Msn2f/O5G7LrdTguC1n47f7KLTxeUhla8Tc+Pu8MYoN4
TZFXshhHWNb7CXnpuTDQ+zmdK/QZuRGBCUItCmTWhfxKBN+TOD6TW2ZH4DcGJ4+uS9HMVSVAQyKu
mPoG6ukvQ7FN7tmKBP6DA9ZB4OYwNCRivWV1L2A6IOOP4dp0+x3pQp07EViFqtN2CqcaXlpjrsOH
GLoXIy7Juyw+YsvldVxA5qURvjDDFj7XQPr0CJqZuBXzVvmlPwFlo+XUJA+dTWWNCG5yp+jNwZvq
uO26piu2rlYp2LkXXbDIVRlw38AJnORnrjbkQIitmwdY491ydunuyvaEcZEkrgJC27awf34BafEb
9B3l728l+6Db6UUxtclg/YiWWYl+Ygg9Zq8EBgvg+Ur8nUvgERABaTOIby2pH93sm4QeSNjBb37B
pfazqIw7xJG4DdLxrPECMeAQaNSrv9cEX/SJDLDWG5zINdJSY794XaveWAiyivLrUVkXXY2vMH6x
lm7qxGE1WovyXO2lFwFCP3IQzt8Fs6wQ2NREtpgxzgNJNEd3Ytq/hs55amhvhB/YT2l8bnLky/NL
HwALRDR3wmG/RU+AcTbTDbJ5Fr81eVd7wxDnid+OlN5+w95C66XetfAGhp+sobOTpxxie3g5pJUj
LHQnN+ojCYJqDwxQTO9qBy5pSdUCI6pQs5zyEgxlCuCjeQFw7nyx9W1gJ0f7zzu5TS6nAO/oS03O
YVYjEebSbt83ikkOdDivmPl0+VMe7R7t66pH3Fq+hcDyn8zasqs1JSKRD7hVDyWKzhauf9o7m5jq
O9jltvpYMKlk/viQNmJQ9TTgflvV+7m0UkFc26dCJkuqvFdq2QnGMkbCtol/GZsFX37VoZmW4gKR
7ezehwDG/xMu0ZY1UM00b9BtfJjvchY++cakCR+K/5ZIS4J/30jbbVROH7fvYOi1jt54BgNCUc8m
dYkD+j5Gbl/cVCU9qxtQpMwl+d2fgc/eQnBsCYvRt3J3VHAABPT05DdZEtN4Pb97Odata07NrK7S
GmYaGfEYBBQDYE69dw/nhxYRJBmG80okvMcw/D2nOMalohYJ+0Mtl6PfYCvjH95lkVe2r+u7Rzbn
Ehz25cFO+Me3JUSvuq6tF5TQmaY9F808gl3pSLfBTEsjpDtPSP93msQQKMvMpw/8v5+54DtiCU3s
+QPlpI5ALCBDP7xx6DyyvRjSv9TrYw5n4j6yCUtc+JKTDcAAXm8Itoc+D90twJxQpV+Cx4lOxyqp
vDxBWxfJ96OGfVYeWjSKIChWBtdBrz52yAq0J6cNsJ6QRFG8/ObXDctdE6q8QkSEfGITSqRsb5T9
PjF57a9nSmxMTi6teb9wt2SMCtV7DPaEKz2rhbDGNQXv9HQ750v7AnlDYmX4ptlin5N3kP7q3Oan
wgc741jC18dm79ZkNqC10NMjK0D8XwimNRKlf/zu0Zz8CqBZh7QYWglD0sZ4SlWhc3WdR7k1RLGf
LmtXdws9nQc4IG5ZzdDnitL8XLgfhzW/FqN+EjnJloLgHgKLSZWwKNPg9ZsdsDZZ3ce76eh5eHvS
rEANPBnmWPtYTDVObh8pdJAvtmvw8aJrvYV2X1FnfqKJl2+Hw5nYXaoslERU0XcidJr5CbQvBy9y
SVBtB7t7KNo/r4FOPBkF32OI4XDGXPPc9yJDdHryKLUVxfd2vbOT6V+ts6OsRMy6CnN9pisYl/EM
sAbXYMyWYb1bJsD1flqP5EmkTSEgQBka7fEBhFg+3lxcmAr2x1nma3YTU2wZe9cozKW4qrZ/L2bg
+509VhTmdLBJgi0QRd8Na/u+GRmMDthHTVf5sAY9d+EA1XNx5HD9+7OXYe5xFenDGYeShdhYG2Ot
t2gdSh4FAI1HWzI04ypEBj7zakZdVhrFtCb92WptMTjSQ5KxqoqgznpcbXtFrUfjoiruwwAePxAs
pwo0NiB858AYae0RuuLMQVOTDuNRER4eUHSsqGhlg+1EL7UzIGnv4ohzmn5pq+si0aLr2X/U4z0n
JXhGodZGox7z5aELXC+239n2aIqq3CaYWkXp3xz/a7GzPYdsV83Ib+NAV2ljJS5NTF4Hn8BWfNdi
Ga7rkV9gV6MX7LMxn9/IAo0AQd0aCaiFVzjAQwRTwmMRJUHr8LoHiWSTYwqb6tjjjUp+M/QWkEvv
IwBDaYoKfJg6F4nBNuscOeiJyvrqwe6ZTnH5zdTiLbOkh7Jjcc2GWOFn6PrHtgm4deSX/jh++n3H
JB0NpCqE0jMPxPza3wkF80nFma4EQ0zBtH4sRHL/rhAdjqT4qcF2TRN+K/riAw7LQJr/FntwlbPl
gN9t6n0eD9ui/cvt8CZMnF0xf6OYdxNT52pzG+9zAfAJr5yaKwickHmYpU/+GVAF45gaXGHhWUmN
fnLq7kvNHXKLrVqjJsh1MINf9yAdzLQg+avQHmyKYOybJ5ZMFjrouK5ys099TKa4Qli7cCw9RFT3
8YPMCf5ESKoSRL5VF7sIZI6NpjNRPE/+wRzxwvf663qeFoFM4Ljpxngqih0tQwpxZbZSyTGCQpZX
LkLh2LZwHqradLzXRJw3SsF9lm8vPVAdqioA1B2bawSjkwG73XScn0qjU/1GAXxYbBKIQQP6drL3
0wvHnnakRk6jRLV0iT0csdNqVlnNbDwxxR7fbrdJM4xj4nm1KnqGXwkSz1QToVSQCrobFKTJpzHC
GaHLRgmCp710f6zf0i125+VLHcRPd7utG4KPAOcTNi24C5cePMGLdem3kPZnMswu3dx5Fr3iF90D
W+VBMSE2qhuQGD1nQwU4UaL4URauf/7d1dEuhFIdrp6njEkpTdXpO7+1M/9/8eO8Witg4iwnfjEj
lb4IQIdBGqd9UnsVGZKrWUa4ozNUafAmyGpvHRxgsv8vf0nCp6/OheZMvaRIO+oX4M49bur34dOm
BQdP6KYY3ttD3y6bWOAAbuEf1KlDJa/glqdcqPJ14RBTJMVu2CXnNFdkoadSr2dfw08lYfkYMLLK
Pzfhskt5/pDmWnNoW8MHbOyfTIhUEafd0424Xry6do+Wlu41wB6UAyWUTwK4xgSLLu/V5/i/8Sph
o/y1w2ATwHz8LU+L9+g4mfhcemIF5rX+B4XydSP8tyhfE59vD3sls/Q4r0oKRORsPlE1NYv3KYos
FYx9gTNE1MeEvhID/rtjdcYCI6VxXbglGS6csO2h5w/O5bJfuqklp7LBsgp+Wp7nuaoifVUGg1hE
e+4v9xa+jMsPV9mlR0cC9RAxJG8IqX7sK5Sxywyd8JaEnDqBe/5Y0zYP6uImBiMmQE1e/QqZ0FOM
BK6DapxSdsqcR9cL9hTJEE7qQSUJ+D71WJHtgK6juOiJB+aQ5oh7TcsuX4GAQ2xktZqtsMiaQn9H
BJDbwa7lv5BlawLZKSJcvMzxZnYv6zBj4rs+26R2imZg0ugbCdC9kaTAx2QcyxX0sdEQP3JR87Xr
7vjsyp3iedoZmvqJr90A3hmtaEdXaiKnlnGfgENigt7wn7E1T7QgvzCwg2w1DYTcJ8tOMe/Q+Y4x
CHRPDoBHKEcco0TJ5glC1D2evBOZW7/RTzFZG6sxKbWRBetv39sa9MqLF2p8+w/GHRT9WMf0OwkX
Cen665hTbayv3AMlZ+FSJ/JwGF+ErD1MTquqR3sSWVjsvFTz3XszKk+Z7TCJXIiycC4zx4f/15Tv
m1EMvcLZwF871SDwgUFsA7vt78BbVcPPYVniHNJwynevD8+HKxYhmbGVHUM/YNI2WkNrrAHDu0o0
Q8yHDbyuTIFapQlgaURQNOtdyO9E4xkQN/NxSeDDKr4vVcNZOtWIrwEJfwMImb0As1mPw6dw3d3i
ICG42OIwuI7Yuh9plk9nQYP7m8ruank1GEx/91aXQYFsUjrVW+iNvSJdPq/X5YTqjdu7uo4IjtWt
jJ3Qzk6V/ALcjA5KLUQ7q0roE3d9o1twgcpLp/r5DHAjzuPwpLopuXfCiAhZm6qlxpFsqRYiZ6qI
TevQa0QMVyqgjWum+V4R7hFWFzuRhzwm+tvgjZsreI34ZcfXhuxbvOvvZVroWie8csXZ3D9z38t1
MFRSh1AI+KK7jN8LBMd6coNyUoCjCzkjgJdzpMZ+neT1G3L22cKUr+1KObwQaU56nlGF22fnrSBh
L5buRxJCaQaPlf1z2VuBPhSZDMprfBrncBsuOWKI7zW2HXvKITv3Qgjg4+Y8uSYVK/hZ3c3/XjkJ
BLg9jtik4Q/E0W0NQBflqIGlwJuGce2+UQd9DSlII7nZz1aJF1KghjAwC9EBvYibhZmXTKoEaVSl
fNRsvV5BXqJq9lVElkJsvs6LFcK598PQOpN/cksHzF6woew5zPdJGyx8SIoVjbmEMzQiKaIqttDQ
HzfLZxie59Ry7lOTlvP/LKNkBPfOtuxRmNt8XVY/FKTljPEHWNyEzDYwH8P4poQkACb0NoLV6ZAR
rTi5ME+cWdl6YNFdDUl/68S0Opt0Q3Hfod690c9v6zHwF6lxaaQ0wJCNLb0MzfKmdtWz6AUTrnBd
qp5n7/XtMTV301asLfMWVhkEvN1p2hlu87BFGUykMGhM0+y7inqCMua9RDXEIwelSOFnZ7tLq0vY
6XoBU3lMYqTSkGQLDVR07zmSaOr0HeNuEt0k7B0/erneAsBjfKVgYxereU+FRH6aUP4PcOr9tdGr
27rhxtqyxFK5BoiHetgVeqF1E0lTYmU/SxNE++h7FBFER+WbXyBzqnOb4cAzzmASepWt8cIVXXvP
nejhR7ho6snON59DLuUxG0nzXTvuv5fUVLzCv2sNvCWB8r1q3ngjTTFb3v+WBr2rzHYWl3w+y83z
2+rFixeu9vyOVHlIe/QPqibhJKG+5SHYyP/fa/xrtzoeBs+ryAnA1KVzU9cU46h5U70spU/jKOls
Y0sZxchw51oEkPjUrqe2uAxkM+XAdSO8gSsYSmuTvUsnAQMDaeJlUc4rg/VDir5f8mLXUE2E6YUa
6p9tykl6eLkKOEDL7gvh6SEsa0xiGd4WkjluokG59Eprz2hTpN4bM9izkk6iVEH6xLsadRQahkGd
UaqoXiVOjChOSbiea2UzAVcKKWMtZ/vJ6Ne/4GCV0QB6ArzHyAF1krrwzuYAThPrTRBbhZvRk6Nk
cP+c9p3yYts/ETa4izfCyGj8kOly/77zwX2rUfmfuldW5ibVl1bbFF66R3esPVxH22kADaVzlW2H
WXrWUdsbDHxji+rX4+oAdn+EqMrMVMXfCUiRf17vtCyqCi0UCHXISyxn3uXpEt+V1LKX6/b8iskZ
nrs0D9mUGjAfRrMKsZEMpUXwhyOsBwqGRj6NeRIuUi9yHKQa4nMHWrosAxxPlNdT/qiVlwS0jaOs
8uk/nrE2WK9OL6W9zNGfMgL7UkO2Imnf/Ze0BnjspG7Us4v/pyXIpw7yHrFEAdUv+WzWf1lPp/ES
uwGNldOs2Z57Zef32qH+dWST02g6ztIKiFOkiR9XTMCMwaz1CdemYrZVEq0YtwjItxAelgFHvgOz
B1mJ/3viHRlX37rddQXzwRudit/6thAKzP2Pa/oug4uS6zuil2fxEXwbjZj4fmKEdMzTAbeM9wZ1
t5lTERiF/tLfCLXlwAgH3NukLi8f/VD1V13HGQYdPAUpalDwL//WbYyvu6XbY3Qj8ABIPT3XdOJW
rISz+kTw4p7T6WKIYwKbQVTJ/vx86STWL8F/jMma0rvmbTkSPAu5ulDQh4kW2/6xQkQpAI1HJ5n2
efuH9huBo+dlLasIDHIfN+trBBFfxmgO9Y+vC0nhiIB+tbthKwdgi6x2asMmN3m39B1ruxTua7+k
Z7s0jQNlf9UEsbnnxbR45so/07YagjH/OJIgovxiT2i77wiSfPzT8nyqpVR/YfIxBGJQufLNubYM
F840c1rvotuHOIBMoXpwWzbafGyB1UwnWE5AWwVwZMU73P+IbS2CHniRyRDLudmOaewsLtnoSvIC
NuG77AiVqnWAJ0lKXlF4obD7dK8ERtTtrDPm58sOwFd4KVUKf0wKjDB+lGqp2Z/mJmN9ZX86lrMU
pBtZpbIcL0/ppzl7ryLZEraGPx3oC9a4o/VtjF0FOQ8zydd6WF8r12nAzb7bamuipWztwIHzaP/f
gWbzPR2cr4wmFNr4zy2Zt103YOZsbMIrW8UUzs9AcflCi3Twf2L0/zlTm63cA6+yVp2XeriYkwVA
8SHt+JLFWBBGjgOJlpAw2Q6sBj4TlbJn7i8kKGnFVTOZhniYewO0niWKyZGF4pNxPamEOoxZr/Cd
5KKW2QMBwpygpj3gIrWipz8OoHi70Kh8mnKoBxeanFsTu6QtzII07695JLb4OGW4rTNkvIGTc4bw
lgcWASJBdzE4dD9cMNQLJwAZagpK2UeqKaY2Wycc9J8mZGe4bLLRcYF7ziqPRc4r36nP+AxN/eBw
KGGcFUE6Ztt/5JBBfwOYR33QTIyiewxJI22+WfwTnE+EaMqZVxZklC7iJv71WBydk+cYo1n5DodS
JCU3EwbqDGJ6iI2Pr3qJu5jDgbkdzhERdGl6BorjTU5DKgD0Rvd09p6Rr4mZSSpEM/+ZWgvIZka1
RyqIyEYU2EHACG14vCae1kxz1+k6rGqUr2bSlasKACfp25Ba/b3Gl/E3iqviioBH6FuKnfCFJbTP
l5wNW1v/CY/0aHX+IZJdjJ3HG2QzdSJLio5HHyNxhSqtZHhcPVPxf5lZH3F6m5e5aHONBCN5qqH6
jSu25ECq86LxE4DXC9bSKn+aRNF9E8Hgu2rBzpFf6QlSRdTnIKXa2R8ZYzhquSfinc9Aypmdqz2T
Pap4JpdUNsnWgyMUge6XE0YRHH69YGgcIq1xC9OwaenYVnhjcrHQ/+8Sd3JXzWo0/GcHyuSx8u+G
taYfPV8RtM3YKwduqWrvvHSCd4SLd+zIsQ7c0p68Rz+DL75C3mpYELhzPNMb2FLlXCHezk14XAsf
Dx4b5gThx3SRBib4a6G0btoGMUvRnXTwauE+mQT3CCZGKqhOdL1Nf1d5oJm8dvUV9OmvLuXUZUwg
RnkoH+ufb2kaiUNAgfBylHklwtYOzmANa5kynO15zTJYu0e/Pjh/5E4Q4pWjvNCfO2h86pcIxD83
OX0kR5AyXrZYLvCr94hTWF/uCgQj6Rv5XaV/+HLZOp4n3ws9s1rBwrjMoMO7/n2ZkiqO8samAE3J
TnG19W7tFm0WEcMpojNvboPmNF3to6Q+RERt6nmws35eEAnZPy33L0QDmNiWUDmXePvkkFatYZjP
27HgSQ6U8lBjxIfrPxiS74/E0xiMIaWZ09Dd/XC0AxUuXH9W0B51B8dKidFSoQWSE5HmkrIAoMYH
AjEyEELN4ky4nfqHou4Ma+3WXxh3cjRqxMFo2aackvKwKezJqpv/qNG71koomPoZB1tuqGFxx078
lUMWOLSsX1CF6CJUHqWUrARm4TI1Qs1VIt9ffRDI5YTe6kKRwgODr5LXzT1WwcrGe3eh7nQHSiLs
3AIKaBazmxyBj72InjGoh43H/HQoOa1B/iPSCI7hg/jgnbXLgXH6w/SvHNPPhBgF77jBA13b547B
0MYPCXe/3bhSSXtLfUFe+CryV9AdaSfTRCsJApBVV3ucUKkasv3PauWQ82QXYX/geGA/5vgsTVhp
PtWyTlWEq9pneen5H0gLCpkIRU2xiwDILVviW1seWz8sDoGjvvx+qGuPThA4dUKitoVYS7Dd6n4I
GG6pR5xqgPx/psRx167ZtH9KmgqfLcyXvCtEKOig5p176O0wHnJyDtPb/m/6AxqspveI99dy/27O
67k+LRaUVfspjtLnzaYThBa1YPBU/p8+vM4BU9KzkX9MDrXeIfYqWGDOhV15CzA8AkaBJBbcutJ4
LVzbXt7w0fphR9mWJxanyg6WvW6wsdKans9BMv+5xsY+Yw23qQTs6uSVtycXq4lU51V+RoEM9F2A
YxN7wdi606kK5p+FGcRCEUJhpCE2DeEaggyWjrLAhl15KOoHmsTc+ner8tQsdEw5TuJWmpGp0sWq
6tHvuWvc3cFHtIzb02VXZoa7YWm/Se4msRtUvvxlf7F9XhdWI+F1QEoQKTIBdi8hZZVx16YKVnI4
09Pa4+xtF7YVPPOMPBQh8x2X87sqCNt5komHy5BW5QTJiUoCmP0gI9qXvx1BN6KUZzZvjzIkPc+i
SQqUYK0ppfW1EzC5M/AU4dkVxrSr6MORooZk2P0OlCxg0liYZKA9QFtVNYShQRYYY17o8qaHpF2Z
gim76UiZD7Mn8YCZIv0/rRxrF0l4hmrkVDV1fgfNPJVlpxxzW27jYzoIjy2bW+G0NAsivY8cCT7m
xxoBhEI17hnV8e9a6Wq5ILwLCy/qFaqCC67qhMs0lLIwxbpt+un2tA5LFHF2g5H/OsAcuU5U5taZ
mPqJN1vXTTDmpCnIj5ZHWL7AF4mWtaVkjrTwGiYxcJP5NaOgq4BEetdymWOlAZYj0Ax+t4Z8Y77J
EZ1O03Ks8XJOkxSymwMEh49Ngh4t9tB90YWko0Z+Cjo9uJDBrvjtLedUoLOiVHeDCzjtBbDQmr+E
PXuWIH51ZvA322R4dprcfJSa1bRersImJLcjUYUhj9/vH8bbMx+oXqLNGF/YWXfMjH6baJdSsIRe
QC9gaj3eYtxmCFKhEAVnFEil+7NpgQUldNITnXdB5aN2tJWR/f70tcYe0wfZWrgc9XG2VKiy7NxY
sZHv/tLtgESN+5yBxQo0jVowvGLn6sQQN3qqhNhgm3xv6src/temhqB0q8r1J0uNtq5X9fK0ehBQ
OgSQIaNVCSH78h6geLr6+9bhG2ytJ0IHLldQ2AhPs5ls8tpNoUZIxrAT2kt7M4PHkAkMa3KP7Aow
WkHE3s35erSCfnKJlXSEO1sM7CLm+pGXsTu2VNNN6rd8w65pmoGT8YGNoYdFoOfxHY0ixVI8jbQ+
PIA2HA4q3BL0pYpCEJTIih4HMutwqTQs6sngfMyoVLd7lPTZ3BXenmt5OO3vr0FGhlnY2KWVkd7F
a22lWSt8LABJulyvX3cGEIZzzuNBEorp8HizqTJeItlXABNlS9nfEVwQVBPz7w8QoudWdWJigFUj
WJfoHQ4Ee1WvavtDZyFwRMBu5Wtq+G44qXwYQG8fe593QqtmC+ctXLkip9+HUILX+/3RqvsWTk1P
VVhqILcaQygLATrTSqP8j8NvukfncFeqoFH9H99LzbyHkVs0yu2ZGHAc0bxomKG7Xyxit/QjVrPl
moo6q+oZd01Mg2vhYI2jE/enuTfBT79HjIclaWRz60y7c0sNEY1qMjnJAF0Z9o1/ANw/oQosCQyC
+HORCM6tC7ABpDqH5seNZIIHAe5D2A3jRBLEBZzuC8VIEPXt7oaRW+GyGoPhCMz/LLW5Ajd5FeeO
0hmu8B5E635E7rlc7skgAUg8uCoRgy+c+ImSS0khVCprAWPIK8XNRXnA/QmSQP4Uov1i0F8q+k14
9vrLq1td0E1BhRAlt/iy2vmNos5qzjbYNizYnbKjQV9hPYNrVd+k7qN6QuJVRx0/k+nbJin2FHmd
nxCL6t4/WJxcGi8VkTUDpc0nPjfKAk18Exen36PhPKP0/v0Xt+fKvvGn3XiWR6Jsz1BbQvVuiN4P
RUWqY5Y2MZJXBcTSx+JDkj+bMMdcjj4tJCX1xMPSfhkImB2cnTmhQ2F3jzw2u2xBSf1QNHiJI3NT
ZCfNVqhdkOvkq0xaYey1NOXXIhp1g46tgPRl/LI4QJhpNhw5lkahpta6biXwDPiPD7n7EuakSoXg
9UH5HSiaWEsj6g8lL92yEmMNLymn0h+cyPlKhJLook7q4aGCMwr1XjVQyGv0E9EJoxRHVC4hcQrh
JVQbIeIIE5ahcfBykvuwMvOWfjB4Gyy234umo/LQ5p76QbX/R2arlgT33CE6SWT+tGo+ys7Vw7gH
qnfPOg8IOIrQyIR8dk/oPJLlLc8ywVVjTWP2NUlHnQu3KTCDXBMS/5hNIj7xFl/Tt5h3Y5DOlTCX
Lzn4Ww+WIshTRHXwNCHFXMymeVrpUWQMXEUPUuL6tUsnd2mj3ZnZqWN/J7cNat1jQOmjK9ThKec0
H3V5kmJoTNwyDlWgTMhhIWgS960lcVOcQTbBZ+xxeEarU6ImegLKZ7Xet/KxL4ndHOCsD9/MKDhv
fkvRV7p9tDmgdmlZeRyS/DqEXJ1gbFx+Tz/XWODgwPN0REHnLGm+5NpPdJYugH4DaODchMXNhV7M
3C0e0dAv8NiRDCNcJ7Rq7XKmZOHuzK/a1gdc1L/ASC4a/Aw+a8qsA5r5ofo6sJRWstRYAeFM77Ah
bzc9812sSKm7gmX4RrDFeLb+NPIQABXK3hjbKFeH2kDgK9bRJHKSPFwyOi5bNIR2Fs8JXPoSAyvx
n+MraEvpDoigH7xAkXb69UDKpFpEW62KdpNTAi16whwm0yg9guYFT8DDgjtQ2geD8WGnER2is4BZ
UDYX+vKgSOvMirpiAi6pm6T31StKF+xqX7EsMq7Bc9aV3KLOhZgG99i1yIqtGH/Yps4V/uAi8X0d
z1au55qyAfV87HVJXejH8THMV/C1jx3hRoIhKokkqwyYBceFnT133Db8eSZkpb1qquG0tQC0EkiR
b7pn39d54TAsEvoYraJqPTsu4meR+JBUC4OKm5np7eCw6T93gAmsvj3PNiBmbx6roRKTfiDl8ERB
Y5ND2hk5P0GoD5jm2/U5iOkzdInyPH6j7JBGFTnmw+GVkMpRK/KLMaAKlOcvMBJ425BStR7HO1xN
x7N9BPqxlROenbR5OLNlelq8X+c3AyTN0bGrSHGF+EKGxSyLTkOIvma6oU9/SsoSIGz3aLR69d8K
/4FRiNnOxdSFqQ/IZxP1XDknvB6/07TlTyWYZJhX8c+FGK2JLFgVzBInoBj/bzkDQLX1grqevOsx
DRqraLgnXjG4tu8JLL+81nOHKLyOXxyHZWZ4ONb97RuHWyRPg3FSwSkAHKWgbSUqWcq+RuGhTCmV
n1wg6ygkXTAL0j2fkCltuSdZN40LUp0dB+vEjcx6i+pW+m7PZ8BsXx+co6Zd0OYT68WcW2WnR447
AhhGNvqaiS1nNhH3oo5J+VPxvr5fBocjEXUm7hk1SUJybpD3+q/zM/lL0qhvhPkCeMkxrnFIlwNd
YfPxFYgNi8jpoYwDacDjrk8RsfOXbOs8DxGZcWUP+EGVuGitHQ5FKAp2gK/5pSiQyBvMU3022Gp+
tAmzVU2z9y0p/oTbcXzWetgD0mPkMVWjoQSHcFA+wKFOuuguPIeJErXjjcLAJlYuA9JD0R/VbHNg
E3baUdu4WrxMNle8SPjUTBPiuyu16sm7bGPT2HKZiR2ON/Jb8nFyf+doTMZ+K/GXUin0Kixm3Lbl
Hpi/8tYvIKDPFQ96dxQBXZ02aeSQjWCyRLiTQi65znrHWQzSefS2ujpGa5CXFUrFcb57AZEEU18U
WygUc1/zoSwZ+CzvZLqewMhF+gXqeflnuSdStKWyu+A7SWx7e9c7WES2pfOYDnfrHV7bOXQIozro
sfdzrOpEqVllt3LYmE0Xzb/z+r3urh0LTHm+QGh6OgzuqM79XoNDNiI8bJJf0VJkV5zlXTfpY7ns
o10G5eYp0evWHLbx0nVVwiXEmwpCRP1knTwlV01MAOua8AXlrMpZHL85YSP/yME9SNgrYvnm8EZD
Sg+eTsVIUvHCFG0qy81fao5Wc6CEA42xtwLPqe0R2zFs7oOMBtP+2jZxZ4kytT/lPXDzYnsI0lBE
U02Fe71CJGe+SDRpD/ll4yGlgXuDmrJkxdNxomLBxqIbY8/ScZa6QNa2MxmGjsw3eqBHRvbLB52N
0WX3VTOSPQu4WoB+k+VsFdopkbUC8iwuBpZouq5WQhaontZvueidKgafhEiMJG8c3+Igzg0J2zk5
gB9FfiA2uMQEe+77HFPMxVA09zImt2bkF/sF2Cbt6kXonT152rVCpC1CZ9765QBcE9CTa23VsPPf
B00Vpsx6zysk77u4bRT2y3g3GWnN/+ld9oKGYgdE9m640NegkVeL4UukLiEq2/egYDXYfbZP/BZb
uzAEwTz89EBQVG6K4NIneJLOqv0DJQLsZgF6rVRPWUm5voGuS6Ud55KzE/g7EwO5JgMOcII6IH2f
1cII0G0kyVRS80j22+t6wSr26mj6N9WliHNrXUAAt5Sa30e5gE82yF38D5fKePmlt6nhTVz7FY93
JNwlFRcCRZ2xJhYHVyRF035sF1i3TzKVGlsDuDfz8eiKiR3gSdn3yikwKQAklTc6POV9dna65E1v
RuBLPwyAyeGcUSuRfLVHSYAziw2XzhdR/uQxghlrzdYUdrlfEMctQH353Sajjqg1hp9EAoEuovRS
Brkg5xX6/t+yuvaNyTZjcNMPEYLCx6le/WNE0MBFUQynpvn0XqfRmc/HYAIHL49CITrh5yVbNUzP
bTsBvlHO+HlM1YhxVavaFEv66xftrTAxhVGWjbnXT7Z7Js2V5RHGEV6tag3qLpgXxoeWz2J5osNf
ydbeGOUg00UGCn66HKU3tHWMp5z4VEy1oavOYm+ETTsJoHBtOh8ltpLB3GusljOdoi4ehvPfktij
HDu0SByQY6mYnjN/3hQ34But3nlBfkMK6k1HEVt4ExgOpvu08AzN3hE6N8abcXq/kwUAK7WcZxCi
rn91B0SYV3saGuTLoMHBgrlhxgdGqZR3PgX2La97YV7ejuULzUCdHKOZJSNabTCJD0e0eIhhhW6k
MrFFJ5SQt3mQ5pdOiuiQYdktS81Pqu8l6QqCDDyGl53WzGPECk48UXu124YUWzUL/jCgpZT+xXFu
+WG0WrwG12rg+skJc1jojAC6QAtNNpuPFDrCWBP43be635WJSADEIoWZh3SWulr3iScP3/VHLSQU
XxnVTAovWPeycKZMf8NAS9AGvmj1Fe8wZInt9cQRoXKnAunIVin/5cTuHJu/4OHLhPms1nMMsEo/
qGfj1ok/BmX72F5P/Ep+oTqNW/VqV3fITjJElpw6DrN+SHDZq9r0q3OwLMf0PNALtTvbJHCSXQBC
WJEPJ2DxZDyRTtXVQUd5LHpHN7b28twbL2JaxQNlWJxy2xVnqI0pHF/KNMyYGgB1gfjOhv9Ok3ba
dGt8t393JDY0pmF8nwV89HGayXe+TUBSfymgRrDs3nGQJgq5ERP1/qzWID8h87Z5CC85l0IEN4k6
i9sQ25V6CN7EhFkBV82RXL87UK6HATLfPZXnUp5jCKBNiMnMPDn70HX55Bm5MuUUBPr+7hbKJHwa
QPimRM04g3lZ5SOqMezp7s8cwlcQl0MZBDZpezff8AlJnIXTRD8wANHwhC7wPJrI/KVm5Z/Mm1AT
ddErum7jvsUs5A4FOkbH9jiGMX3RrTomCjrQcyF3sV9359sM5OKBDuQEDc5TnvKkiOaNVxWhyATQ
0/+l9XweDBi2YTq0lPIGc18WE0d4DrCZxPKhOtCFlTLuk07Vv2AiE99jNZEEUctPRd8FYHulZWjs
2lKjMCCTq3exQsEzqeVeg/p+yIrvX/7XxFSbwUResjJcG+xeFPgNv6lbHphg3yY0oQHWUL9zICPa
08BCfnecEPJ+Hww9A4ktdcXYTxZorkfIptatM/OutmLqvQRwrslLfSTUKJ98BMq/LwEi7D7PkWTz
ul+ZtO8KQremeNkSrViovuP4zboIWKr7+NBVI5s1wbe9VPH1LnMlLzh0cjFt5u28KTEY1TeFZBOV
TABFbQ9BF/U5EY4yPMRwWFnwylKNwomS8N7vMscfEu5ichoSJzl0xbs17KYUnKjqITN31dZ9UyHs
MWI+78DqjGfJF8U0k9ITsV1tM9lGjEB6GQTUUwvOfrGG/xjb5gFq3ozzzUzMIvh0eXsyk20t1nhQ
LpeIIxfE/qAbgBlx8DSUzwRoDeMGsM+zFgdoYSa2lZnJp7sH1SytI4bPasgSSfQz/ukE986qAPG9
Nw2aDJx4ev3UBV2v0n810dwHUXsOaXMSQPnIozs6nMU2GORnX2h4XtwncBMXWHO9toKdBxt30xXi
JUq5+eh+zhpzjXIFPbJL5juJ1X1dGESJxcjwkRepSJxKqZjtgjdXNL+ceyygSCI2K7jFH+PCnfDT
FJw4ffuJ/xxvnE+KZ2h7BLTJJ9JoXOmD185rLne/KFeCiFKlO1dgpYGsT6+c4sJubA1PtVJEmxec
y0wqdFMDsCe0AbxJVN/OMr+4CJd2MD7pvHr7ftE3g3i5EgX+pq5A9JPUCHYPUaarAuCyDUmA9szp
9xTkhcZvgpxrsUWwjHb1ezI9BSCdl9zfLIAfz1/Hm8yVw93XPsdu79QUhtSOOqQ9ryHb5U1KaTOl
3YjPJcRCTQLAfrn/IDhRNavyzFRWKFpGTWNT+JkgWMYYPDfKCe5rK7OKPDN4QyHgNupKzJi4vCJf
yHkQ9h5Jjkoeroldczr+gAxLwYjqY6p1aFlKJ+gvSgAYeqk3vIVB0uNNvrXg0HF2iD0cqUzDCd0U
s92DkAf93ZGwpMNH1UZC6TJP2ZeGzka9ap5IvnR8JSng9eA2kutJcM4wBJHF0gFEJ9d7y11JbfNw
PRoYZeS7J2u0UoiFg5E8N+Zbcf3xtQYWJdGXVPEVcXIaQhzra/Edo+KQthwaqfCU9ZLygi1Rv3tz
dF5zA32+S1Xu6RFgE0PEIrqliQtV0BLkXg4KcfAqWsOtEnCV50vYXIurtZE3tgso8HbrLlz/Bpkr
AM5fV8Wk2Vmpa74QD1E6yJeRn2RLnA8QfO8ZvcqEIjfUSIJ/fZKwICModsZwbkug9RysjU/HJQye
UyBMSPy+Vg+je+Yf3ExDvtfnU8Lrc6YO1ooXMVsTvM0X9k2UmdLw7tO80jc24jTmLeFpqfi3hVw1
mTX3gxaPS1xI5efKXUC1WB9Iow3g+1wcTF0XBaMQD1UBsaZ1Saxuz7arg1LqL/asxbsUd5MhtucY
Qy41FnIGGlDTVBey5tVoOtGhPSVw5nRXQV+LpDrNmcWOjn9JLyuJs72RKF7xxT6Y1F2g5kiwM4o/
Cs716ZbQ2QC8UMWOr0iIjZmSPjkESpvzaXR8e8tsfy/Y3j5gPIp+jIdQcqbxcjh2XsasnxMBaR60
tHulrEBGadJTzOyuBaBe84dz5wvyYvsQa4cZ20CK1XXymdTJD9JXsQpyf8++Rw+PMdEn1qdEfw4L
wQXm7wGmVhD8kdgC7pCXSb7Q0YrWM8d2D+35MqCbiOz85MqEMiblq4/iY2mpxshm+pazROM6QZiL
o6xOOLoileGr9f5MUgTGtd4UMN99idS1SnVs7tT9OWpXUA7VUZb6siLQUevDNm9dVHmdwog308Dz
xDgogLGVUwUYyownRzBYLCgz4DcdM6QIMKzrdKdGKxDaLDhlzgxanw+Hy0TsYmUHlklOwFn4OHhD
4PP5WzPRVS4LweXdTukEDtzA5zmujHqC0v8CtB0lwwtFDP6vl0uIfkrTyAmiGp7ZD3ufYYyaoaFR
DVkRxDZbm0nuEg8j0FJ+1w0acC+EtfOoevbfyVIbwyeXN+Bw7sxbgxC3nZnl3qPh//+qU+bIdhPd
pAykkZMZYahfknbHUL7lF7IIlZOEwhI2pBoKN3r5sGbgDgDtsk6uvu1cOorC1Esv3KyNso0tvdwo
Ego1sSbsvRbFvWqOb5fdT22AvN16Jh2RAPXRh46ImEdEouTG1WGqyQSm4ut1/zr9loDKUYtr20ll
aHX4AO9FpUi4Uuq1X4r+X0RZB6GOJIorxt6wLghtGwmr88jVSbXYV4vJLkwkhxPNC86eGwq/Mn7N
oyDqtyXigylpuK+/Slz5EaTDZxbJiPXapYhAUTJyIFRHdoIyr2neG0x53qfa9OGe9yt+Q8dA1iUB
8ZOthsPglQW0ZqOTNP9BKyq0a0EyaAGLRozwvBns38h17CsVoEs/J5K7rxkwu9Z8mK6M1JWBj8mn
P0OhKG0zlRugPzzOAMuW+XitXuDr7IsCM+UnC24iiTRgNtMR4uJ5+i9JGNc3Bw72aSrmZzwCXEDZ
OgBu+d39iZkXnTlj/69/JE7Lde8pWXa6e1J9qjGTdWgBmbvNW3Kl9bRYSbivL/IwAWgezx9n31KR
vKY59K6g19xKs+Mtzl/QrSarm2JbxPPDGTBG/H9Gi5TvgKQmOoJjqQ3U49/xRPdcayboKQLAUVQO
2Bjud+OvGb+jfHAayTiOkIqTIymXFISdKBM4lMvCCr9Tyym8M+i9aVyzxRXb0xDpHo9el7nlogd6
AnQIMCN2fOK9xPg4IqJY5C0wwEKeRVN2gy94D3Bf6ntq9t3IGpYlc3BiCgdkJdcLuZLgTYRA1Lcb
2I/j/EevndaZi69B5IJR1EGB94B/S68PmACH665osD+gbaVmMmyXFU6PyIT++AJjRJS/zWHS3/WC
mXW2cPUtfmtkBjxRU8glNAPUdPruzb6QieJUu2on1+LLBjwWkfEklAugiIDlgL0qCqd3A8GDiB7H
X++1Y3H6hVU/gRu96fVU6elbaSxjEY31kvOoyJ/WmYp+OVwNlymA88BWTBqL71RLUf0ug1PHqGej
euTvVwt9xesEx6w0AzgAISFK9pWAjE7s7Avp8TBxKTlEnAUqokyHXor0+siNeyRkNmUEDTJyB6Zz
+HNa9Rysqzbjx2dVLfgLuY/NWMkzzqBPWhSvmYZUDtBuTVwnhH8DbP4mXbsOBCbGYXXIYFQ4O/hG
6TWibfij+Lv/6b/hCf4jdbzpB+rPCKNM6VeyJUZ/qbSNYLE9lJgNZGduQjjeWBW5A7GThTe4cGOF
0qDjwSJwmCMvfp7K5TrZVOeTRMj7CVQgTA1HyKlaLULh7wIGxFcwqz3P9YE3ACjGT43wX4rwuN0c
o+ym93RgvTglY/4ILJUr1sYjvEefL9tZ/UnPNF/qznhm6cFojg3CROZ6FnHArmUVvBOokQHZ6Xjo
q8O9I8oc6W3H0bbfDMCWWgApTxUN2ienXDlzCOersmx0p6+L3MTkij/wEsYrv8/sxQ96Zhhjj6zB
RzhKonBqwK47liURDAphD+9lNLsnwJqF7GJxg326JDwSYU++3kTVKpkWDRNuF+oNJ1gXd03gk/IK
ryw7647cNLaEnUat5oEWEvWrPm9SuWokeFKT/gw7alz/QhrSpBqsmHRvghmXy8f8mbNyGLxhuGlc
vq7sfbw7xGIhDzCYaDtaBs228Ypj/TXOOipXPx7d3gRZPBV9uDuZtDXDgIfE1Gp0hQzrTmNma5fP
MDHxnUFhFb12PKXXK6V5m+PIeSyHjuCHQJhdqRyllTJMtFFVZEam6z3qRf9CmEmpFLHotHy49Tpl
6OM84R/u8324Tayo84rwFp6Dx09eEH7cLX3sM8t7lEV/+0tZ1cwZ0JKjgq1jNjfZDBeY9e0qfURd
vI9cHzj5CuAwYX8MEFtYlgPB9LqaMlQTxu7uJG4D9LOyRlZ+Q6RdT1mSnNfI3KIqcspEhOTMfwE3
eiPrnIMfxwJFgOl5D3hBBgFzBYdY7LJ9jD+O95hImPVeoXnmsRcCYBvzBc56p5o6QHayvggv7bn4
6vDQfrj1bfsnPMFENec/2/yP/RhiVh6sdV/3aTYfrLfUeiC19i9LKqqEM11A14b0O0j7RVPCOYLr
N88/tzZMPnbOJ4CYuKthQHx5KBObRgSO/8JwWviGRsULULGAGoVnFgSpJ1MMp99iATT6Lv65C1f2
ifFmoIAlI0AePhRcqPUJXyvbYQsU9rwyFnLl7uDCD41qe6IxZtuWHWra1mm0oXWoKniD8H470oBF
MeN2S/Y3mHUcjHgQWYkIAgwk0e+HWqe9tRynH+zG6gZSb3XER+7FlBw8D6+Ve1T84K+yH8fmkoic
GJ3UV0b5AcoP2tVLkGXE4ntaXMmj+3rHLFTR8D2+nbChCRbbOcjKW4S+pznhH6LAzv2UOYFUs9fa
j+5YkhUbcvLZYcxsA5njHnTbE8jsubI9OpktynNQ9w742Gw4A9Ut9jQqVyns46micL04sIIKHBdw
WmHk3Rz/ixLcSqMEo5X1Q25Jt7TN1ilHZWEzqinoekSZZhohcQusdrUoUda6LKAXZAOfPqv6Tygl
mIUSx6wizX7Mr222R/7PRSSseBeU9lsoN02PqIT0oA6KFtaZQDZjprVJ26dospl+5LqRivV2cW/g
6L1VsZYU3ZepXzhlxM9rZ65cQCikolOkmBxVedtK15hqkaabL5p2yHm2xk4hae2BXegLZsCn3N/9
7bUNVAKcIX5J9mZLncprUxbdimCgqp5EmMBQAFFy2zSxiX/RZ+JXfaZ771kQ2pPTi/GmdC/BO/OP
rEyX7LJQdg2U2iqnk9LyHUZnWiic1bCcqYlVVzgf8zJnq1TBcx3HO8GPKTfooTe3t0zDHo9sFTNZ
uJcn4ITRli2e3MlJE3BpudULgaXHdR2sJeyJ4UDClTcZ4UsjZlBHgYahdksh9+jzGFH2GBawr7i9
7jsDuAxrjLF/x+1J/GN+kMczHDsy1c/a9tQGPRVf9l0MXDO6f7hD/GRYeM5Rs7dUaopyptfSL8T7
bMzT60x+hw/Zh4ifyYpz1c3Suwez1lr3LWv8I742br1AqJ61h/nMmpEiGDDefez3hTPjLY3r7Nwv
ejlPVCHWTpcA3JCQfKXQA/4G4BPnIYRhEIUJDDmqhC6j8TlZ8iJBz4QmQKM1Z8YER5euMvccLf7J
UFL+rtUfJlebTbUV8warr9kd2uE8H+rfNIzUwV/w4ksF5jyjGw12fR2zjxS9Vp7BCMc7amNjvb9E
JffBM1px0u9hQx/NSW3iKSC8465/KVTtMPLuen+hK9sOisM6hpiqNlsG7221TlJSg7pWJ8OjeG52
rsPzNARqfk7aKCWYdxZKkyC+1/4vR3I23Uz+49DFlfXZYCR/zHpoPiIkjXqAnZzeD25UnqfSO7fO
jBF/TWKNCsTc5WQWhdK7zXy7sY9jB7PlOLMVyZ4OvFlvQK34XYlOOUT41arU+qmLAf8wwh5IeaY4
r+bd0BAqr66lkX8TsxzUbjqyD9V612fugJYUQd2yA2SgBJH+mjCqbbSKz4p1r7ymoj4kFEkG440W
ALePrAfGqyEpVbMUMiZns7o3eCYBDWQco2DeTW4kH5kvPDEorlKoqDvj/WV5SGO3Rs+c5KiQJUJB
vnm7zY2gU4XSOlM0NLSl7YvFMu3Hh5grWT0K+Of24VBYqdIVKsaSbgojIjL6F536nmtgh+NV2AQm
b7JLYC0cmxeQn20KCUylhSgf26YsyZwMHI8oFLh32bqLSr7AYnhPFhLO8kb0CcTao2mlEGGLllEx
3OEQYQ81wOH4ik5h/qFIObT3/Q5s7zv/ikzgUW27zFZS3tPhHGN4EqgnH2q2Ei6J9XNUdpjhs5So
4imwDGpspMvBX9TZ1M4g28q1R8Te5LsmlHdoZGySAlyrcmyRsmbP3euf+gI+Kq5l3itAXQ4rsWL3
YgiZUj9PiH+VZYHgmuH0bDvZH60IkS8VxC/5JBVgUhWSvxC1vGKT1pwuimJJuJrp9r+QeHNf9R/A
XM5mgBAEHW3Dr3QiWtokIpAOyLTVGlh/mpwLHMAJvJ9HmXTbjr6uOSJrmhArUv07RVhZAPYuNkm9
t5R/05MLK3W/MDJCIHNPjNnkkDX3o8KQfCdQhEEayxASy1h/4lUsTHV+VBHrZ0A4VNZt4M9cmQpp
+Fe9D+rGN6VpJSleZ9BKOCBsk7e/OlqnJZgMj1am/E7SZ2A51zwVz6HG0b4NCAVzIWygiQEynDtg
ebeTfrCls0ZuP+f+vvMkTyEzDVufiqL8JdduJEyLzhqOV8iDxmaZ/qivcHUoprXbzEVzx5QRV3h8
0gmhL9x+72rGTBV9fwSehV3gSEPMeapESwYe3tm3L4DbLAKuUVvhauNXt94RqvOs6ooJmE/zWITC
z4srV4JexIccCnFUaCzrS9w8gadb+iDLmvt3d1fytEYo+X6NF0Sb8gyZ8iaslQA+fhf/n77f4Fak
ZUHimygTvyZKVScvT2sazvw+TL0V+8a+7D415un3uIfGpo+w3cm7t6mS2iE1VNuZdGd+kqghhiwA
u0yHeM8AbdQ3ZBevFRa+Sezs5XdbvjuXNughYcLmVJRiI3QAxOpbV7c6P6l/saVR2saJpPDquf9j
0NXrdaLaTZQLh3rL7oS0zPTZrXwzkAfwYaBsAVnmDe7dzAca0fHZHOnF97BH6gN87fT7DYdoOxkf
gTCXenhfYCAHJxp6GimDQMp394T9nsfYlhc+C/HlZCO8kSvpHQV4IspFhiQfO0HClHniQ4pU8CaI
FPYEY9Eam2y4wTEyOjHBTxrA58i8zoJnLWnOyoV5SnIDC2nPpsSlKt4HgYLkYlkxOzeKq6ctuqiH
nCbJYvcBau9Cn5e350OEgnocSOoE6UDUc/81cAmc3V044k8gU4DoqeqG7Zfj7ar7XQX+IV4M54mT
aIFKP8DM0hLymCD/MnUgpxLHd94FPEH+ZJIvtdaDVvqz+/Ja9BXKwqidy3e+HBW3JNkEYkASalGA
jNFcuKhf/ew7d+EKg/ZIEEcBqmh4tqLk98hL1QFNyAnmYhn9HKhmU5NfQfQOqvKnfWuauUol+Wur
k7Kb7un5z6gwcOYUXRxUrtCI/Oohxg7BToqeHk+eMN6QnNBYC71pkh3sUdGWoX+IU+2x/1XuBG/f
/AIpVq3RXt2ezdYFi9+kmQ3NBhb7NkTjd3eUF+F7saLXkDQyqBsGcA9CXZ2XY+R3gtRsvra+DEaY
6SZ9/ybOMlkl7IB+FcwKaZjq/v/sqXI9Kcx0puwIDCo5X/oCirVz/Vo6kwbo7YYV59d1x0BES2yH
uRXx2cU53ZRkTrSmm2JgN9Rcefd+NzVaCl/V8/4Eeq1/w93XUcdFubItSTYhizZWt4v00lCLXWz7
Mn+1lishMlEAyAj2eCVwcj/on2coBUVYx55Y5zR9fFpw/BanZPQEwNpZHD3Do+beU6ucOohdVB4G
STmJw8xtYcntziHSxV51AtuOHDoWSMWsFD3O5XfiI+PFOve1Ckmc6gBNTacoWKY0/SOdE9gstSG6
d6K7K3DIazXVwA39fmfMjGyr5UBvcfGT9zmlANFORiTe2icZz0ISBz9y+kNxbTkCI8z8Lbl95z4V
wjTbXtT1YG4UKSzUNs3a28XNckWBFd7IZT5sKz6rzokqLQkM00LcYxSSM7jHkcqxvliTyYdhGT7g
H8E8JAKda5i+yEtI+EV9pI/cpMTDZvuJLMUq+RUNTn8HHM2lXDCdHq57gW2N3YGMYsy8vf9qDBbE
Lj/FeVyKn6SurlzscaOvWLgPwsAXXVJbRy8ZXZgXDot2t45N4sYj5woNLGRSsSierTRN9ZRo0sUn
+bYJ92dXHey/WEH9bUwpo+gBuQzmwRReXA4UNi2wQWN3/CzjxssiKmHfam82EOC4zVmPKaYZ9mCH
T7zwBQaPtC821RLRnlxcdPkiHTrhwhe70Rwco+kV75NS/tVm1Gm+ZxKEihRUXHOze2N98HTIURWx
NBb8yPJb2HVEDcW7Wg8NEFJAtdyNBLBgFEu3YEcDiNyx5DmcelloPrvJFdp63UBw2vpngYAyiZM+
e4tkuiZIp9PfS1JSEgUMLNr4/q36McSL4jj1bJVx1Dou5pFJUj8XbXbruUGHZFzaNWuWOo2I8fb+
UJb2QLItbnGmEf9GBG2/D1vRZrQ/YoIxaNpYSesD1D9hHNf2849hATcqQFXSR8/hV8LCd09Y+C4v
mw3G9Ke+36huuHcJdwa3Kx+v45c7DJNb6WSiEtTKYLW4mwZAvxasL4uKsclZ2A4deC/OxueCWf1/
oxHu9lEmvKRo/AzUyuckz1BjQbO78i91sbNQD3nP4/mQLbJOopeDOgBxRvg/CrtcM43obLwpy2t9
CKoTQTyOAMDt0GRP39Eim69L5dgG7lFpjg3inxbaWafrDocuTYaWFHoQmvEb31b/V1YU/lLQBi/6
dKTU3S8U1mVMehS1PYvUtXjL0QW00fpLIqLbrh8U0LaLzGRTR1IaNsj5H6+PwdGzOw37M0d8ZIm9
YymbCOXSp4bcZLL0D/LSrZF+kc9Jiq4NbvHXLuTQazA1sRamn/x8nPdng+zUzivMF0Z5CWfb8BzT
CXpgxmqEiD64ktnD0x0+MlZCKXqxCbRJMEv7dwV0fxYciRNPPzeX3Wl06htIQk41mbQqFpIve4fT
bcHv2wEVbfPqwpWVe56ItF4QmDRHBWxwEgU3RYVLqClnMprpuJK5ilBa7y6oqWPRYBE/xsbOtaLK
9o+69xriuYVvzsWq4lSTFNc9cZivcmvQJoXxBRD1RwarYdt2hYPTwLHivBabxphBMlKLXhW7iA+T
eY/t3sJyD9iXDRgwNB8ZpvWtUJKk3IbeaUK6hP74F7t+0bVqucPNVNRrfr+0Erff2nNowtdmErw0
G6zb//M/ptNXcOfqeVHoNLZj+8LVM2U8VgZoBUFXmPz1D4nPhXLN8Oe9BQ3iI0Nis7W7oYw8uYz6
7/Fzc0kiskffv2AfAUBVTySp7LrZykW3dgrZ5lTaVdPg2lM2GWht8QeBtODjVhxLV8B/QJWWzBXV
/tvZsU9pGKbxF1zW+xELvqjbyoYOdopXqY2Aq7DZf3NRrcqVzyymvUM1vrsCzXIq7FWDb+g3yZqB
lQ34IRYrk9KzVVZ9sqih5X9I7fvlJCLtagBCLjz+90M3VMQvffOHLenlkMMBJKQ7fcLs5IkopNDA
B31+ZivXup/zefJXeBZLag8VVqg2TkizEFtO22Is/plLmzZSf1PegWjW+aqSLPuMFMvTtbV4x7Js
TOzTHGQvCS1ocJ8baOZ4MS+2/9xpkWSr4ofhD9n8Oo3/t/d45NCRke0rRkcDoEkwEtP6fIl9wA8B
893VgJliJ5I3QUgDxhaghMe6IuC7wjMVbwlF5Y27n/8sR/2KRaZx4h4ybIEmeLDl3PASqrzceNBM
Ey9HINYjMUUct2dFRTdLuiZ1nHYbeKRyGOM2eafX+pm8IM1O+osZrMW3AuRxVCoBydfga59d3K9A
glb5dU1V6glfn802CUoEPI5t7Khst9nSJZdhmKy51WImca1WYnlFg4O8ePWSbjSvpQK6bzp9LKL0
uDR5ERmGyZDVhUmyQ2S3k+pefIPrXOjxxPV9+S3Y5AGLLoKVEg5QNVZRtuBHKsbOLSfwvrI2Pi1V
ZU9LTVyGKHEmQ7rS+lh7HhRxEOf8teVJv6Rj4gZ6FBAPRsxkaqMvAFYchLsfZHzqvmAYhG1l4czW
fU9nCZH9PePrDAB2Y1j/vZ7jkOySCLMTy/vQaN29b7wp84Kzlowho0Eiey6mb0F49TJGBc9fwf1C
FyPd7qTeAkElCk+qafDK3vKfWEIN9NkRrmPTo4P9CIrx/KDcO0XTCJ6ESNtqXFZmUZBlze5Khl9F
UikqSw6kAxkbJnZzIqF6x+DemLL5W6WtxqAQUJv3ERKcHKfs420L6eqD+ruxFGBY7KDsHW1rh9PQ
petxsQ/35zllYvhQ3K6kZWwA9dD3A0pIaUXmELgBOO9hyesv1F2VqG4iHAZ6gsODQcHkwCpQIZrF
VJ5XOLmkKN4KnQ2sjPRj5QOZNe1SxvOj+OiCP89nWfDfRO+okRpQg67YpWxFRMszPfvP873nk5DL
T7UKgnLcdb2gQF5MZZvaNNvxx12Sv6TuKeNlOoc8HUZyPqPKjMGlvvxUMabHRWXWy1g/09z9xYvD
/p7t66oVRp5G7C2e7DsKDsSxUXuM43rSoMH5sOK9e52om+I6HyzPyXnkb5NX2sscYOYa7A+mdX1P
Fej0MwDF3/9OxJZvnPkEdBt+thB3Ld9sW3MzALMdkF4Rg9huRrjZBBWOeRnTpsUx239wEze1TmpR
D9fg0dYjSUjO8duJVkQXqg7p1IB/fGzf6VG8qxlVwLSYSeF0nD4vBaot20s0GcGHLjwRXCaoy+mv
ZgQ4kYpgZGvVDROQmiVPaCMyEXQ57Nh1xkvIpxG0z9vX0D9b1oSEuWSq1reYHV0Rr1Dxeh2ACdDr
gFXWoDHjn8mk3dZWpPmTRFmy4tE7L7GS96zvSnYRgkTSE+UiMFnECCwDXHgbDW2rait/t7fHE39u
MzaA9qnIX7Ov70rM1joQlSBUV7rm06sCPy58jXk4JAjH4ebL5FBxJ1JtAYxbadjNJKFGsCm/C7x7
8sk3qa79IwVLKlg007jIxI01xzJpxpodIxJKkBiNSHg6DtE+VGaffk9of+1iOgoT0p78sg0lP2Bq
qgi9O1xSjBbFKMe4BMUWKtTy5I4FmQw283Pz8Nq5Tp1y1rdMonGjscSZhs3yQ5D7vXHn/T6WnpLC
nRIP8HblXjDMPH/v49M/rhbvJ6lzx3oteUETRTPOmvZ65jmOLoU3vmVOrDn4KW3kjP8xxIYZJ7jA
OQAiP1bVE8pRX2JisBk72vCOmA0oqIqxnbE5Gzujl449TXnmg9omKvuENeUSV8wBvdENJ+PXbWsO
ydEsFEBHEjtokGDks5cSGxviplWVKHa6Sey061YFOzVRR7MVQb3LDRTy/7uB7GF4nkY+Qk3wMnHy
xAtBIL1Gou0dysIJ55tCLw81qCzRVvuTpmikM4z3GDrenxH3kmVa2L9bWwEMCIG6KRs3oOGpIia0
nFBcExTsVakgjfFiw/0+wUorVBGKnsD3XC9TSMnZWEVhfni70USrijY1ItA3zvZpnXVbXG57Q6CN
4jAT40bNVVVgZKWcZMfdXE18gtDCi9P96yoBauX754a1RV7MvCG5CgI84hQ0lhxIzHDX/Sq98DGH
Qg0OcKHMJuPMWjW1z38DO/C7fDQTqx6CYn1A1cThKt43JLUxMh+2RVeKEY3JBWsDc62ul6xgBbyp
qU6Voj8fAt/DWjpm88sllz9WdW0BXN9VNJ/zN4B40oHS1QFdAaRQKcX25v42rZTeX6pA/feepVKn
CYt8nKIuTyOtHlowTW4D3WUmXIBoydNxGNFx1iqMGCtbHPJxDG/TvkkattyAWLEmY1jpmUNOF/xJ
eVltpm9rVpSCfHMPvucYFPnE1OfpByl/lsMK6ka0Wi4JnzYaAWPHgqyEwSbzPXcNFHtdxyyrBBBm
QS43eaE5dUsI3GF+WTKcAUK1bUbxQkVkS57UFfVwXNpc0OS9/KVLAgbhN3KuBQ31f3A/LIEVBp6E
pDHv4ActmeSGEOxPwRaml6D9Xrnyi6sOGlU+J1Fm9WI/7B8dSeQ9kZj98+R26gHRH4C/nmeEw52s
enSZwhxnF9pPgB4VfSlsTpG00yWLxVl3GCRZuJVUomBOOksFDL8o2KdUsQXo2D5FWvZJpOFPrUeV
vz6c+ekmFka0lEpqlZ0nEHtr5i+7gnM0VuGmebCJDVDPWqXXBn7GS6945kXbPA+UYGvtmeDqdTaA
9b+0t4YC2YcfTD/iiPf2Xd86MzCy7EI9F/qm/r6rIdhD4fOjhEL6snrOTcQT/2LWIRTpVeLJXm+6
9f6pRpaNjFXmMW21lLy/ZpqsnSijmErkZn2OFMJNV47n5L2Lt0pS7eaKUnKwLByl4HdIA+7cXdIV
LqEbZAveO8TOIiRvYrfZQdqEvlzJGNjrZlaj50U6R7TrFXToipbQc/902kFFOyqMiLxlLPENJn2q
cGudm3PzWLkz1rNBHPaDdHhpeNjqgYR/iBej0r6zalM6mMLX0JeEe43U1Y6kjbbkU+mxX07efq0X
1ghkRKJLMU1AUm9JzS5yAZgG3kf3MqnscUVFA5tks1COG3Jxk+EoV8/32O/AhEdZRG/DmMPSNhZk
zK9EdFaF35ZvArG0AqnG4o78hxwc3tx7jkSuwLmsB94VPNcuESXK5+yUuHb+BWpaLmTaHQvf0w+3
L9I7I3kLR7JLkxtAZybh8gex7IUZiknIalHArFPzqFxxNgNoRHj3ZuIGG0bLNIkEh5DG6/LWU4Dc
fMrH4rXcnSVHishjUNBYE9tFc/JUezel1h8Olhd4It9bYzKTuBSC3+rc/oFDtPUZ0Sc9Y/Y5O6dO
lpIkDb4oKLdJaj6BI9pkU+K61SAPf9Mzr/PXOhfQqHE5A5CX6Djf0krXoPdmPDNL3rtcdhuEtsIs
4wOxJVplL8pKccMaEBZE5M8D47SPt1QnClDVwttJLjBS5VShT78H9wtxC6uPRjvcb5ihN2aPZE3i
9jN5mNG98Xk1PnDuFZoDdKU7dDwvTBQYJkfgAw+Xf039pmGmqbKAkRpNiNkbsCrPxcSh3zjcR6B3
enuLiy1wHwBWx2yNjHi1/rgVMX/ZmDgVRs2ZGUwcsm03AxhBlRCmdGl6crmy3G7XAbs1GzYn2fqs
aOthhfrfs5dwaiDnGoR9fDOaRbUHrvCjQxq4Uj2WBV2kRb7EW/tTBM1CHe5Qdn9UV8bPP80eLGu2
jhWhtxVYfg+HQLNmZVrVP8q1Xx47MJ8aoRjlkvXf+6E8m2sWQaIzUJ4MChOMOx+63oNChcPS6C38
qjByh4I/P68MDerwrl3PJKiZbp4qWPDQJffkK9X/bubdmczoso7pRNnOTc764och2WlVNy4fErHi
hJNVWI79K6yOy03dEK2nTV7xNB4kz/UWFk/S+WLqK4UGOmMChGFCojyIZqud2X//01pmzaaigt8V
et5viOBJYURaaAvM8aapH1myLPIcS5OVOqcLZ8ZcedC4ava1NlquUB0J7gnfZ6hY543gRyheRu4+
K7gvqn4Vf1wqvnfLAnNwVMpZdD6rqcaRx1c2zJL/mkpa2czPXGfEura6ouf0X9lMztGNPAD/nD/0
0Y6/Gje7GcdZoLvNFID5Pzgg8QaQkxBEzrD8e1lc9XdQPtokG9nR9HZaMnB3c2cVJQBZ8YQ4JAhR
r0bFYtj7l0JWHZqoMAd1EKj/cqF1v/hHdOiGrMU5PTkcfJaOaJQ6+xmWbMB+fsR7chRkYgnmJClz
8XSAoYHUSxLAasL4pSbwsd25dun30NtSQTRsjOBN/T4/12laPtll9W+tuD+2K5gn4+J0Db92QuyY
YYvywMLx/AjKQpFX8m/KzGzrX5mwHNxIvuRRfIbiwXD3tlsaneb/OVpYcVqjlAGoolmmEOXdI1IP
p6tTO/1s68ZUX/tDIKHjAELV2ZTZfixQKSoc9TJO+H6xKg0aXyNT+USZtp1R3PE/GTjZNBY93ho1
wCVSW3ic3+OAz7FK9bXuGbvSBKS2S+TpFXJr3WrlP3jpR9W4S5m3WjwkuhQrFcApJ2VlWpOJGWAf
bMOHBpX87SchbfAwzSWVuHt2esSTH8RYzIq2yb90zi1eWvW2MK1oetvhIT5pP9akdk0uw8wux0kz
C+czUGYNEm/iAMDVfDI5UalFBch7pON7U6owoGI1xycdRLjfcxzUE7IH0jSFt1NKKMqCRakDSUml
LUfOeuJ/PiBcyD2Ve8qGZQeaDmZEtQgZD0GnuNxEe8grruJtAgEXlHItZtLVSCQueepwOeuo6+CW
qTJvJ8wWlXb4we8uuBuaDbvj2FwELYOcS556ZBn8/MoPi7AfXrX0lsTK5rz5Se+eLzElLYPB0EHI
an5uk50rg8fa//ewk4IJSbPFIMX9s3DeYMftCofuffSw4nG7391F2GzNqqlMHgQds4OXxraJaV4z
QUp+rI/cmLfwGkqUp7afr+uLv7/Fg9KZXylt7pBZvKO6fMwh2ypSjZAvgvx6xZ5HJyqJLq45JO72
kJYGBl1pI3yJhR9ISGRt0I77dmJEt+KktfItKpG2tIyRg0L6F4ptW3S95kVAq2TpE1CS23cqaoJA
64o4MNPRCyzn2AVt5Mf79uT2cvYqeJWTNBk3JnZBIxLimpRQBEiJRoqWHJah5MesZEAypiEZ0LPW
2zgKTB4MWxzXeBppGiDbDffufmUr3imepy3LF+94bQ3XagpQA114J6Twgt6XSV1xTk06wZg1yf9/
N5tj8xzSyqkCEo/XEv/Xm89BSCJmM6g1B8bwRmcilwrWpaZM1HtZZ0pSJNpiRPikn94o/6PH7ZZW
UiW/FCdTRD1OXJP7SErWfwqY6WCUun3d0/wfFscpL4WgxFD1aDk+4lscFdKP6DWs1FH78TepZrul
/3qHGjlOwBfNVlP5308PvPjLC96rA+GBLaMLUIisNn2nO+X0rL/EWprnlCAUMBO/d45VcVppE8Sf
TIN2LNVqYgfTeLxO5cKAQjxtr8NflgRzZFxgCweAeeFyhSu9HO6WtjUGN1JCAPv/CjcCbpwaqjzh
C8fnJqtMHBcZPKVp8M4hF91XJKkEUR8jMhBVUPoCbn9xBO69sr5NCtSS9yBRcflo8yO7chiRUNJP
UIIO61gXMiqW8vT7tFwOBmUu/NLx3Crcga8zcbT187aeJ08EhVfqYEu0mc2BhJuLDFwWReq2EiDk
8WrEFX2bc56fz4ZKZf/5ovRhGky8qoaAz21fu0/SSEy1qvuIUryyGVyWvE5hHV8a2vpeKKQc1FPC
JcEQ0tjk9XojyQQqnK26DfQlsnQk8UJt1gsRz6PWxkDx8XxizgUS5EU5P16jMIOUj3Gp0Oo91mK/
NvfZqqttUCPJbOCLK636KIb7Ibd1ZpFajlHMTgF1I09fY+RYS5BOrFYpC2vlFZktIy58x47iC6he
UN5s8Zelzo1+WOB5Ggjgcku1E8I2PO9R/BSRyVdtTIBep0GfhT0baxi6CkGa0/uFdAMuKNgEOmNA
RtNKGaSEHmAsA7PzvtIpxgtCinPFe2jgKMn8N3TmppEx7z41vcGMoKm8qnln+Nfq57z/xS40Utsz
Cbn6a7wM+uzj7X//N1lD5yQbZ6C9yEjTPaVMr2v71yEwZ+DJVTbGsb5tYF/XM56HXuLrhbWPESH1
Et46C2NTYiPZsXZVZ5h/45Qa47Fu5jT0q9EDyRq2mKhUZJRNGK2AJxyMimq2luh1BhX9+A2T34G/
0ceA/usiFDiHjkn4yi1Lgv025wV4F1BV7f7BXkSffQ6mtFjdoiTpBQu1+/wCzQ3Ye9PyyjjNVCHM
XSOdmFseZH7s6MWbdvEf4OcfEuztgMS0PoCgAn9VEhsOAkMjUMLp36wBz/bmxzBd24gprytEasZX
v9Ncjl6gxo1GiA6GeUJJ+9EIO74cKYdGOXJl6k3GohF+ulP7kHG9Ijz3vyapDApdAgOqozTJ5EkK
ctZys7oeqVloAH3Z/n/1QyewEL7AADKIUNNmyrWxeCELNn2h76RqSnXruSy5HUMZKzxcX7jJgFUH
5fxSyRgeviwqhcCdM5cyznWNALUbHClR4AvcnVfEUmvsWHy8wPEpytg+PJ62McJPode8qulsn/o0
iJAvBmWVYwCnDb15CVGJKv84abWRCFZhf3Dl5om4lMb7aN5luCq23Y92gq35DBpFeeUt7C9HQyc8
SxSy9qATaZSaBCN+NuAYNsYr+fOFL7xC9TSZ4kbnmCM2JQTuvh+BzV6rRl57ux/GN/DJxGa+MoKx
gbRwcG88VgIKMBaHWCh1bRgRuFm5/CsZ+w09qyLviyO8yLfywJYHuJnaa5wAA9bEqA7sHL75aRYq
cTz0wVQU0yUlZzu9p4gfhsffY5mQdgb3lMtX55ZcxhBi2zXXJS1pmhNPEcGHTScponpMd4fpulXY
OAVsOWlecIZ0734OXnVFzY2Cyf+fqxfLG2Yw1mYZs2c7QwLtKpomv2fEpQzhelnh/XpQCVkuCEoJ
b9M5LO8jXU3LeQTmRUDZ1OO3CpKi6B4+hkzXgUj9Tjta4WyLgI+PVozJvYO9aBAljgYgicPhL9zg
GuVqnEiFPYwf0AArw8a+cuHd3fMU7H1AX8h0b+b5VR6Hb+3qSzTyXbOp1KSBF4JBHab7OCq3HWWE
30hSlIX9tig7APpzHRWL3IbL+NlcuxvD5Eo4/qk4ToiI1YW6KnU0an7U0RRek63afnxdeBPS2t+9
DY9zKamdI/y4rbAjeoKIjsVwDWNrsgcHj7FtgXpLKyonesMN/DshjLGtI8hRwqVMCQjYP5Qc/tYD
jD3I/JZkEoEn1tJ5iwNmptlORzxfrUBZKm/hmiiIAN6lL0/9sQFS/BwIfgIiDyvwM84+JO+JSes5
DdjCozpQGeUaNDIFho64X5elayNEvapAAFLWDbzrIBKxJfgD1HiBuhGf+6RR5IbocL+up9gDgJvU
hB6tZOA9ThJg1FxHk+evzEdkMykKyPj7164hUXZSg5h0TujSUDno0ujkkwqS9b1ycYXY3WZXHdFF
TtegbBkAp92poHtcjMerxSl1coLS/7JaK38TiDQdB+9Y00nd8BoY+WotJLOwXe6YJ9e8E58quSTu
oQWRtC479EU3kz+o3I2vD9DKd9zkQdrv/+Un/QeIF7A84UX2BDHIFYfMEK8zehyqP7TfZHGPCJg8
klIemxBDP7EP+u2CeP1xQcE1XwqXgHa7dKkTN2QHRFkWY5F0XlT+m6cBJ1BgY+UTD4buS5YzF3sA
hPx/yRqggIEHh//Ba2TkHHV+bN5dFguVuCvNWmFGiFmx0KqHwbaoyGAYbA7tj7go8WCfQHTcmRdF
X4gcLsth5vgN2nve1gzjv+VZM+WmWTqBKmcZ+iEqyCYd54tSmtdMDukVeHa+H37BvHZDspZ6J2nh
zgubKUm0Ja13q+Ohrpdk4RyZWFDSYxjMIgSixvKOxfV0ya+chcqPzEuklUaOAQ+dNzY33MTCUS6r
FyTU32PLVlamtgO4RBYRutjmdp7WptHxZDeoVCup06eMWIxLQdOQfp54IQoVteVeHfZXrBF+YEbX
/1zmlL0cp5Fp7ciaTHzxJk+wstinqOtVebNg2uUl1IrCD1UF91l0REqtdIduW1uFRmi9N9xHfLXS
7v23lrDDbKcZnd5/aw4uGkASEYxAUlg8EAfPTpRy8BdQ7pHidCOkJzUgt+gdtY4Dwkji2FwKtndN
CMGOSXEP4rdhjmmYT5RbpMOuM/26/oh/WwsGsIi56FMEjNeW2WeL19IU11vc6sZgLnAlnqvPYASc
zWHdcVG6D1GUS3rgsdupPx5b0CE3SSWbIibr5JY5bF7/y6xxpK1REDVuYB/ZKMpGuWyiT6IgxbW8
Tlo3ika0eBjv37F+p5mxlwj6IMcuaU06ECQT1O7llnOS+fgZvbSqmob2Nr0q2E6XsO2ZFERzK/bC
j3FG4iVdPwsM7CXvltLC/2eaSJmED+xIFz298EUvd31HaedwCTTdAVt13MZkV8mC849DPKzF4KdR
RUoPkhZvOPmwMOafXPLThK5hAp3cxsPaRmTt/Qdv4O7KZiIAruM78ORxtjXkCG1gF+VBd1RlBCs9
QDfmVmdpoIRUdUYQdw3iaQNy19u298T/DGy+QBzF8zbz2KARfXJsxFHBExuUP3/RKd2rdgR0dEoa
hFdreXOxAE9WgHmGhZFZPgtLFs/ylMntX4pTL6ZmgNtd+AXvM9quiWVOozVMTWNvw60qUd2gKTdS
l+65N/OcIebKb/UJmUjCwyF28hbnDRW/KPVj1O1Y0jbj3n5LbAH4rfFXPHKo7Cc4fFe/mkA+dxDF
TUGXFox7YsUCnQPxECfToO1r/DFdwUQEtliZ7il0lX/S/vcn6wzq8pX2u1H3Ny9eaQS2PG1ymUEQ
YINyHtIBSY0uebTqVD9yZ17ium8OWm21VxU9DwL95KSgnPJZU7fR738/McPV32ML9PPfoYImWtBV
IQcY1prbAB6Glv6s3Xap0G9ofm8F7qBHp/Pk1maA0o/ruQUmKsOtFHO3qFWhBzfehwfg16xdKwME
XXCrBRwgwFrCxmhOe0qEvPMpIy4YEOu3a6zdwmGo2rMPrL08qTSu6T/1i6Uh8fvup0FOq4az1zqH
0akJKtfmaX7YmznVxqY+SrgBNEGjvulZP1CB1Lf0mOySJeRACX11pJD81bFwLnTD5hfb/BNYzyCN
2pOmK7CCqyPftg88rYWl54ZwZzgotqyb5ZI8bViJ4UwjiDRmkxFYiP0nk+pLBTyzMZ7iVzaW9+fr
rVwHc1qwiWPpGK3v9qqAB0iqoVgw2ZZ5a+s5unOCXBqJbCyiSmeGny4/dgFAtYpNO/KvRUstqg0h
b/QbpmF9nZujbv1+LHg7Mizlp1PQsKNmHv1cVj3NXW511qBFlGGpVVIW56SKVvHV3kkfuf679GHC
iwNpEOfAt+uQd20XwtdjZdvHXJPK1LoD6KcqcaEjRI3X+P4tjrBl5p/482UJBjdW0bA+z3/NNqng
+WjTMN7Aomuo/Eq46+5jxm14G+2qwdCSyfJ9UjgnUlmQw9J5ySAeqXc5sizJeI2XzC07xGr8IORF
2QE1UygImawchbJqsSWea3xVKZpACwGTv9ko82QL4FbfhzApa8ebOkcPv82Y+EowjW4PwKQFbaz4
/ggMGFEiPAuAyMeBM6KyLMyGRn0zuagMyCoKP9dqw6HBFgutdd9QVpLvuQJUct7jIRGJA56mFP91
Qln3ASg4GanPhL8NbOslceSVIwr2Z9efsR2pa22kg7kjFhHIkOGMq2M37EL45djdtJq9Mf5h6qLG
Gk8nQI0o2xAiDFSNVB94bhZhTIrQahp4Bi/gTn/evVWttfH71BjO7WLGJupuM3RzKsQyqkaLHfP/
gnmh6VskwTIVICyOeA+LNGVVotpGo+Dzh6DyT+UdeOMlrhXgGsRMRRTM6Ffgnc/V9PhLawvKOzqj
xcYkL0xr6tjaEkBDObqZ3ph/O/OLuv8DOqDFlShiN3r6FdYSloQS09aewWJf5OkCo1xguO+lkEUf
R8gp5Vqpzji7KnfFz3ER/y8+pf3VVzWqjCIHm+57wglHgj+mGH7m6fgz4pzGscCyx/T5P5GyWQ28
LSixl051oDjJbipI8Vd5YAVxp2E0FrWqejllcK4oFzrD5sU48gzSBoZMRizXu9HtrL1sqgQ0q6sm
4FGi5G9aYXUkfKWuIYG4ueKEI0inKgwcnjVuA/ignGGqCxgCoji7cGS+sV8XVF5WhVSAAAvni2YW
tdkchQuz51QfnRouji/IEchqs0qPFoF1klW3aDZL8ODctixrrp/KcWL1McCP1n0Io6AdR7G4KcNb
H6H/HBcVCf5nzGs57dqZvW9qx2GbxiZ6Y40caoWokZSx5kYVlRMDrDs2bfnu3L4zy2n+fdr4M58l
tqjVw9iHQhJuT1HOjj7y2X2lQ+VkdKVAUfgQJ8+MEU2InT/qyyYrOPpRtdLZiMO8NFNzS5Vr0RcD
IZxXREwP9OxEtzzB+ayzY6fp/Eu/9w+sDrhmlTp8dw0q8JeO1STmuspf2fKuycuVsCla/iY7Hu9V
UaXIXUHBN3pUdBqyeexB/CXlbpA+u0sRc5Y0FapWUrkQ9wC8wEL+/jdll1WGM0KAZ6Dx636Fgt88
iWmhHbv3ahG+TwRK4X+v3AvsrfgvxK/BS8M9Hrvek+wH0obIeoHXbdAYUFqKiujzOQeXSFwFWLe/
2+8GWJzxSHsJSacXA7esPuda26NO2Vsx0nt1WpcaSU+Jc4hB/7hMd8tNum88SLH6BffqdkCL81A4
ScmAcubdlgpEPARZ60WiYxqyVzS3G4mhLB7vN1OssegW9WLCnHmUAZpa2ockA1ikja8c+ilSroyt
+eD9uQO9OJ/upONqaY++vpBVqcBRtxZu/Xn/q0t4yGIRJQtboUM8yqJtyqD2ApfHS8MgPSepm5O8
qoLBXefLvwD8jtu6DDEuS0gKkvcsf5b6nPdKYR4AHUzv5SkCi4ClPXfMHshL2FlK1mC3cFpPI75+
sfSTQznSkQqA6/0R7V4lT7D/Btyxp9C+y73XyBFzTSJub91KAHqJiIAUs+w5DOapKnGuFtLLtJtR
PQTxQ3MBx/4h2o0OFdBi+RsxubM7KfXyHsAe1WelyWTMM199neK5usbeYRofj694N1KgZBP5yL0z
DPj9ahvo4uQuHZYbWHF2JRfM1yImirw9sg4dXj1FtP/9Gk59XNUZ1d9+QIgxJ6+C1mfd81XXP4g7
EMG0T6utOWrnU+7uNXqZMlHkPKrX3SEAaFyAiYCDLOzpvmoCXTfd7do7a+h68DId1B47bOPXq2Ah
M0mFcjBvY0ImVifjGxDm0BUPnMd3uLm6sl4qcqVjrX9nOm6qOKEllsO+YWRDZNEdsduhFxLgH7sp
bcyGFYNdiQU7XTJNKNjaoYRQoJ98vXeSO2aVZ9CwB0zOjXXm48Xoup2H2CzF7Pa13sOAVHbrsFQ3
39Q/TAAvrMNDYPxl8q4AN1lK0cNH66ZO93arYUBIGgNbpjsO6B1+Jocdg9hqTGaueE0dITGF1Z3c
ZXNYKh2nEfDfbKmZy1nBtrF+5fpBtST2eaEgc5UhYddcyLkmSMEPQyqNlvboCncbrKqW2bfkhOzY
FBL0FUAOXxqBo7VRCiXuEiHKFWH3pO8zxs+RSGtXq7B0HsA36Yk45mcmDPDQqAV5spf4IkVGF786
bNuMlHu8yUNssWj+siZCgA9U8Niw95W6QHxUSjqsEqHnJRbLKY3Rr/bHcyNsc3bEWWB2ygKimp34
2qE8zv394jA/3oASzGDJNK4wWi7kWuW09MynQXatTBW65y+pV4Du40QxrbMZplLNONtvPvkWFJVc
yt45E07TvimbKzqAELbH7ByFWa3Z3h+fBCdoXAv6rhRE/BaoflRgNIlziThyBNGWxtkEh6o1/m/W
x1pZp8Dny5puTmKttKX25ELnZOwkxJKmnB/T7rwqN36ZafxI6n3Cx+L+gkXdKuS4vNa1NOY8qEQy
io9IFq8LIqwKnJA6NaUHuQC7/dtgTyqp0ZWqzLXVpZcbFbNIh2QfuXosYnPxfwkaez97HMJs3jWO
3BpN0CSGc20h+MTLcdv/qLE5QCnCHLEynxWAtrcdw5IvgAKej7KyRvclCND4aoufPkVeQc51yuz9
2x/yqQPOKDTXoIbF2pI+p5xf+OinhHzTtlXr4/ogEhUiOzsX2Ko3oWL/SfkNwdbif6udQz/m8sGa
OCtsOkWFiEypsjKbeefksLiqAgZgC/yq7uUEgFh+5nZy/9eptQhHM3lv0P9wdgNa3voOKjMfQL5G
E5fCJ1DMubcjOTqHEEdgTob6F2gwE578yMUkni9rIB77SQgXv7i6Emswl25THo0MHma5cG2phDTO
G+XCSu2U7faR86ykSlnXJjC/QTVWfAqhXzU7x7YTvKcAvTLKp9oAXR1OqOhF0U50XVn5TjlKzEg/
KKjNCZNeL5qV30ZEcZKU+MWXB+5R/Lz1Ck+43DF615QN7CTirA1oQwUr2xbwV7xoceeZDYK9ddaB
xo1F67uFf1uvEjlswtBxLDmwHKkXQrqjWhUPlHCehRb8wqmL1GQ8UlFEHRyACN7tH9EeZlDFVS3e
DbwvL/qsAzu95t/nwRnvsfm23UXhYf2vYyB+BJMukcgpmQz59ehqG7mtre9r3TjmowENznrP43Uo
FiJhQLNbDAxBLcB5JOl6H3DVts+hB4TQW/txgQXU7qSl7WMQtlV3b7nodBkTYKMqBqoHA0UZM3RZ
/hz5Nw31tOEFgluKP0QtF9af1ZJhSz+WKOUlMkGQ5xMavBteQdMCm5lEn+cJo2umICzX45+VmQEi
LdEC3m0tg1dJWldmwpLIHw81Jvt0u/iIBzd1Y8QUYsX32uF/Tk1mJGESQh0FrzX9Z+B7vXncfLub
mlO3VdqKXfK436t4EL5CgWV5XyDd17XEljCeohSUdqg24eKazE86JMrb8qOkC0tIeNOnusrRXhfY
tKfK1J7culzY/q98nztAxurauzQ4mA2iB1gHNejM0r1r7r29Auc/MafBmI9esEjpoPeKZaRxUkS3
dENKFZuXjEw+wcNDyZLsagO/IMI/lk90OrY3O4ZJ2YF+YPy6UWz0D0H8Sf5kziEYZ5y1EBJ1tWqM
TIElVzfsQgGtL9cGGjrko9htPpGsdLQI8zDe1BZuqaXdxRozAwS+x75zPva5UZVXerskZ+YrEPxo
1/yVaJPzyhjDHab0Cs8yyk13rnqCexGMJ3+QSuST039PiuH7WcG6chMWMgkw6mwVthrpnYBZX473
lqM0kuWfYPvg7HfNdDiK5tLmgwjk73u2yAEAmMhd1N2TB0zh6aQcoRXUC8Qj7QQk3A9YRSnmnltk
dZmS4axv5cVEJyac7YpM7bSj/eyQ/nqy8eVu874RMx4qluOKMNMHpFj/2uEp/I+Mv+PkcHOua2P9
9rICVUL8Lo+OoMEfo+7yOlTcuDPWgibwsBgORME0gZDJd9uYOAP96XvQEWRA3RjwIdcCXtwGRQ75
tN0hhnS85Whbxk2+25seqsbUFYcUBn6LWS5xzbp1NbuwGkGozb3F06ILp2hcPmeOVhGKcE4B9bWD
foLTBNAgpIibTAzArr02LYD20yQJPzRBpIIuh/bUXWTWwv0fh4+PQgfCR6P0yHMVs3/WZGUeY7O6
dvShdz+KhgrKbxSpy446Kq9k5wAsom2HR5n5npdYIqUZb04TzGj59UmM8iXnWKyJtAkSYVrpauCd
F4HXumZ0NtqgFwg/PUZTtg6118AxJF7toruRQgEHce6BiJzHLbR1bfweQ9rTsDCEhL3EP8gmJ/2w
SdQfeeyVejGnVXEgusFNxhvT80lGoqtR9Z/EYVszwnynzDUTrnneb5JKEtlgkO5FSb6y98ZTIXCG
9HHwgJL0ng5vQ1UxWAsumxEwZwFhC9PFtm0dfpG2fvrZRz0LnHZ7WRrp4X0clbk22Y+6FqiX0C1f
`protect end_protected

