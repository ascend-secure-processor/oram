

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N4pO7f/y5DQ/0OV89xtvgdHuyCLtXNOAURxfDelB6Bm0My0l9A3F2dDapjVn6qk6UIjRBInhpDns
6v8eZdGmog==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JaFVfX2+fy7c3yrZKJNKoQhXzMP5N0vz+MDP+AmqnrlpwAvsDGLYJs+Q4wHKCZ4nHNx59Hcfxlmi
eCrCAaRfpez++OOWIcxn7/8fJnz1ltE8JeAUg1yPwxB0xsDNH2SnWskcYgoGO0HRbim3dxkUe/YH
GkzhX6HzNkoANJhjFjo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v5cFJP9zqSpxZ+TKhkSH49RVF3aXsGIpoBiK0fmtl0WKq4YmRcab9LIk8WvCmuHvU+9VoJO9tOc1
nGkU2saSawdCwaKhsuG6NKJCqiIWmNpDCzvMX1edDysRggV1xGKlGRxccEJSkoFZL1i35RLZw1Kd
fBHTuSOYkPqlFyh+yrZwryo0bAAztIvVgPtvyEd/8Zaq58HOQPHMjkSgsM5dsQHZIfT8HMcWcq65
1zj8ioxXSIuS/+61XEYCJO6RbScc2yYz0SgdkrhBLACVhLKYFG7HZdJbpGE1NzdUaNNSkjo1r84B
EH38K/sqfrTiQ+oTqy4s0YTN/RthPv/COXrgPQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qc42FDfbSzbSWOsPC7eUpuAf2Fcfof5nY8ElOZpbBTxljsFUwFU8NYY9oHzNkQUA27O32P4l/9Kd
pniEn31prlu7/F0x68bZfHO7wdHY+fP/cLSodF0H2+ph9yuYf8cDYiyYEpCkXvKWbdYnnZe7Zxas
mALDAXAuxHn0gEIjqmo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YyhcDZ+TxLiwTbR60JcWOOHsaf38CpLCWqnuC9NQVZ3QsF2pB8dsYeksy7Ho760wBfHyaqUpHJX3
JG/B48KuHJbsy1vJMAAFMU4xTqMyaLYi0GI89v8MjugOjc8X7ViA7SbczaOeLXanXeexOi0Ehk1x
JdBSFHFwgd3YfK4mMvdE2tmhNgaxF2PRJBuG0yiZQgIaWxQSjItV5lYi+m3laAT3GFw8CRK3FT1c
TPFaSfg3ZklEgDEPVvuSFiPjFM7I4MZ9HW1NsS/ccG5xZcg5mwaor2SQkrZM6NdXk/SOPy3frrfc
tIoOI2HTdFcG1KjlVF0VW4zUZ1sMdE25tNAidQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54432)
`protect data_block
ALlT2O9GXmfYcMDsGYETbqhtAj+wjb0t5MmmrFZT5Q8Bg1wXgsAVAshb7D9HieFR2jJFtLstVeTd
gcyg54NX5gY5qmFPan3ErDrxF78QdxKxJq1puE+qlj6C8aenKWplwVueHB5SzOcGpjxiJBmB4F4Y
bvAtLCB2arRxd2itLSCWSYf+DIJpzJZPWC82HGjXTT1TtL0/XshZRXFLBRxJOkLYJKOvVX+MjNsu
3eZ4iF+65AHou7gGtBbhIw/Mkg6W1Y/O6S6+SobRaROC7AqtWk9ipiLwrRAi2o4Y3ZURJlUR/ezJ
nvlSn4CkTaQQPYUwl3ZF0Xl91OEMZLfsogEDjrtEMLfAUUA17OSR9eat2387c4aItum3jgiRRxa2
zJL0BSRfXo+mOhFek+z0jlQ3OBudoXQiCGIiOEW7pV7L/UZg3W/j+zRm3CkAzcC1l1u0Bg4VfF94
z/6BM0bs+VNdiJbTzIeFy7DtWyQBwrZuWFK8fgljFNY1tQwAMFVSL+WlsYQXxuJCkkL/VPhy7BC1
DFo0U5wUJqdR5MfWbF1VjKQyOhtKQVg+6HNwNoKkwlAT0lU9LNuKcgYxVgSOXWk2ygeyor6eoKKz
x5/FblZrFT7+gnpQmRrjW4j11t0UwDlhJnvzebm8dqJA+ZccSXNzKyCP9hGeZU/10CoXqmK8qj2W
FomEhG4/N2rMYMwQyun9wH5lW06duCirlF3eQebpV/onhDLBLn9w/3OPnpMrhTl5ElEV7UB9CVX5
imWKnVwuxFJm5z+/1KrvHl0eEqpMZIFFXvHKV62lm+LTAlyvpminIa8BPIpYDo/VsYTuzJlfOl+6
X3tfyKFhrCBVZ5dJ55D98QERJWi+ABGMNakVar+3xU8H0rAeHvh35h48kWKZt1hzMDpnJfBpUzwH
5RNqg5vXnrdItLJtUUMJfsxF01akBBKbJTgoHj2/oxx0qcM5fJhI06vK5zs2F8x0uyWM9lfdimGs
aBFqI7iMtaOflmxAU5Vc5GCHtluc5HdWy0G9nURDWeqLUYJUySRjFnWfvGHqP4VU8BN+0Gg/rCbl
zWOBcXIOm4fAJ3C2NNIQnbBX26vl5qakf/b6qgmXH+y+iTlnS+4r9Ke3++nBU/T3OipqEInr8Nqb
TK9BMiJx6NilkBRL1gRAMCIEMiR6bNeOOxOKvrYUi9E5nm9/BmBvOS4Rx7H/fy4E1UiYaEl0b0dl
ppRho8tCuDLxepmxaPrntfMXlroeiOWJDpuXfQTbRikFxCDNnxy1BMtFf212yCfL3O7ikVj/hYHi
BuzOYJmJYDZ6F8pda9yZQl7x4HLyn/2J2nzL3AOA+3itW4yEFMX+ftey9aTUyQ88PX5sQj9WwPI9
onq75hvznF+azjmq19TLsFDRy9lQuGPF0ALW54q+Y6UhDKlix0jWnKhTdMdCYp2VD2T/A4s9ur2x
vyWi5acb+yYTYfOM6OU0d6UZRJPZF1jbAzUyxn/Ai4prMB/OyMyRzIFHopt6qlYXCBqBmF09IFx8
cey9oUblATR2hGezGqHFeSR4CdKP1dpSTWTU6xjFK9+Qsy3mANrmJdt7u7cqTEeKwYe+jU7oX56g
PIB9EOx956h/3SZCJ3NfEbwabIBym2I+wea6TVTmOtF7MI6GrBeIggiUGa3clDvNbg7Dgkc2HJTm
R8l+p4b+UTg+NWehby/2ma+tY9ezK7DwSHRbA/cXx7v+tDnzJ41IvNgLGq9yu00uKM4xfMgV+grU
Csk1osZKFApqGVpUYIosJar98CkfYQ7YWiChGIHHaXH3LmCWe7S6dv9n7h6mm0CoMR9mHLz7sQlu
+sq9Zlgjat4TaK1VZSp3ZkXARzTDuqUV6uqqssrEYylnqor4X9ffU7+VEufKpJiuIpAhdkZ7Utku
46TnQ9sbCMTM8voZmnAIaJsG3OCgJGxypXqiAu83m/eSJSMuxD0apZ78GePhhiiyRO3qOxDrJDKm
OPUCu3cT4snjkgOs+/ECLJaj3shpbLs7vweG6GroPZ4pBHeupymGQW3IiUlEx7DeKm0bvnvoVa+z
y75weYuXy9jq8nDNJEK17MITQ4lWnJFaksJXjkrnhxd+2r12VlglqRfqP5hmYRHG00wHNh62yVRU
Hc2TBrslqX+4OOg6HunrDG2MDWskkrXIzf4IGZe5zpP+4oqs3qzwFz50/VjiegqOOLGIHDVrZfhE
+tsUWnKp9Xc7Fgo2JcNL6cOSnp9FehdsMYHe2TLEnMgHgxp8JScTnErvpIyAPo+b4ZOU83g+ro5x
rJghgRgqefkGITOmAR6WacJH0M73QQAxuK5j8Psjt0qZ6OtdsBrakz8fSW0juLcgRgeSLh1BZPTB
NcJ1YnSoEhET6+rd6NkGFBvfu9aY6T1ag1ZX6tgTQQzarjCNFYMjb+Wx3KPbjp9kVvtgIiu5yOLJ
huENfqanB6rEZroPaJVdE6cZlNH95xuGN2QNcf3fKVvtiKTj03MDo6KzbxQaQod7/j5sf1YD2j+d
MU14iykFGdJH1tol5culcdbWRJ0rwolePa/tyF/q+5VMsQrowC5PWHMSKLxH0KZujDnqPLwMOeeV
Dfi75JErkIMvpl45aguJElal7qdkIbZN1ygL+uXkJ0AUCR1jF/sXUkoDg0FzXVfDru+JyNevqWc5
dXr0pv3huLo7EkvRm8w+DQlRx5EK/FmMxgB+iqxnY5UXtnDiCbjmCEz2s303jz2ao6xqLLYmoOID
dbYZ5SFtIk+k8XD1FOjJOfWFKbT/Khxo+Mfzi4yuNloEdYG3ozM19o1O9QNUjb2D+xOLZklOXi0j
tKUryiG0Hrfv+Jx/QvmRXLJL+7BOOu56TX/oZFIz7AADKPG6fpGLh05YkHWf0907wNqsg+G015qo
rxs4TUlurRkH/YZPCzBBG2a/9VgkNHJjasSLoooiLIPcgJT3UZFFgKYoJGShNRehF3qAHIoUojXJ
b7QM3hEgGl2mM5yoWwkylEAG00LPWbANyinhyox9tOTteU7OzplAVd0BgiWfnYLRdjvvoWqLDS9d
ABgoL9sT8Si1ugvGdKrbvC5xyAkHoTd0lLJDt+pkxumRa3fEUU1fItt6wX965cqxwbRorXlBolDB
ybLS9QVR71iZ0yiU48ZBpangSOheULQheMZgow01iH7b00NGacvd1b2qPj77dqgb8FMcaomZh52u
T6/AOb81s5xScHfMcJ4oksSlzjk5/Ptf7dS/zqqvj9nUecH5LiQe33EIEAoWaEkzZ90K18fhYLjv
zzfeSIrqs44DSqUVzCfGS++md1j/SAUXO0KkBJi6ioYE78m69N8d61YuPfKWd5AlIH5uuvEKmOme
12t8qPyBgFq3YiLMB1mFBGLMDnGTt07DOlNqvwdiwgY/zEtI8Tf/yL2WRo1MEiTnyhcWc8oj/+9V
joH9w9Rl1Khf0ExQldFt7rg/RghzIFHXNzbA4iJbCX9beR4YPng/KhG9R2NSp9ZwiDQ6eObIPiUl
msHSEyrCE7L86IYHrVfQVLUoUKhUFGQPM/kNFfnsTa8Nfnhi0YQPeqX5B76AiDck/wAbWeystbMF
dUxQHnP/se3bDz7wVDlJYIn/10Pt2ITltbNaaKLAWKmNBBcB6QwB1XHyvR2Kkeou0wuRhYXUWOuF
9bpmrxHPex8dICtSzFGKnLuVyspqOCzVV0mnH8vk1z8oyfZxJiv8f1ATPymv2cp5s5qz3nDKn53e
UAWvh1VWpT+1yGPZ72+ZmoCxXyGC79QlY2HN0JL+uAy4JgvesG50Ix/1R6b9Ad2piVB9NDE9eokt
fiwch4vuwdqRH0PiBIEqmTVD5Ltt+TSHEPdLXzTGbBeA2hE9kQy2pGmI4QU/c8QvpjyldpYLAVUI
atRpvRC19SazV5KJ2cp1zaM17jItVA9B4d24DTKzsWDgKjuePOFvajSumdg252Z3bLEkUMx7JIOk
YoptjJCWAFwvHpRp2olWr4akifVdqr3GXvsVhy1GcbyDyY21Nj4UdcaefNG0xwhgkr9b/d5YKs2v
ADxOH+JkEEMDKYx4C+X2bO3sjgko+Aodt4Ddrgon/7b7GvYLlaVPLh5aPT69Bc9g2OyhkHAo+YZw
c4QWDPZQn22zZjOf9SaQX9YFc48Pd5p1ywAkeD8K2JT06GnPIJ2VStG5NZp9QwgSYifRTeZOUOrL
DXpSgWA60bYK44rIzmvMFBlNDBzoW34VRTdCesPz1GiVS5MQkALZMpd8MaRZmtTT1Av1IB7a1AMg
ipDNwiaYglS0j1aaeeqhKszKKAQ/s2XQ0ZylzM9cM9JhXCCXIBI8eUES1al4RaVDPTMOL/mccknQ
4L8DbBMVPEhmcIncZUIWZMUxmfRBs+v5qC7OWVs2D2yPKBNSU+aYZ8g+Zsaz1a+Jgynui4KXSAsE
zTPNsyDcWmUg21ZKdZIFjhWGxbHfRFaP7PZX+S+dSeEEso90XpA1UOmvGGJHaiaAeo03bbeCSmR5
xmA5mR1kh2XddTfwPwqnX9brAv844MY318NNY+uz9Jk0VwjBliwgVO9j0U0/hHSlOrwSCCjB1uEp
/4Xl0X3xXiUH0Z4u+sNUpGsLUxvngWqZIpHS/YPBMIB7xHRXaNHBG4aR0HMczupcNAtIog7jZKJr
ZcISqw4xc7GTq++bJUcZepW0AYKc/oi8gOaSGd8VGyNt2/y+A3ZH+eTYL4bp8tDqdY7cO0OZwFjZ
K6PICXMNGY2JYzioogiZvIhcJu66/RVvvNC6Zn0VcrHi+6u1VmqTmDQaXMKUxHwVptjkriZBZxrh
y2+RJ4uDKd21oFk8lmdZNoRGiMI5d3obQM8+DNXmhHKfnPCoEeKa9XicjKgf4UWgkfpg/rOFY6wx
IQUzWK25JREhRm2mP3uU0NcqE49/D2ojYpu7OJKCChkmqc8UMnXykqYLaxmgmffsJWcoQfU361+e
CGSd2MC8Tg7OyUHWR5MYVFB8Cm+OU3/yEWFYKZMzjIq1PgQhkOU7szhq26y+j1Tb9rKItKE2f1oP
7qMbalcGkSyuQ+whQcY6mihBOvXApaVjKJi6LwdV0Sw51fP5VvSnF7/7Qh3nFguST3EAr+HzBGb1
3cD+fE7F10d6TKEWBV5gPzPtVvJfgHHdxb6iZio0xw8quFR2M/2PgBjd9MwOJSJvhKIC3S0Yvldj
JQyzX36MSn1VNzwwmAQ9yFK7QVNaitg4p4Wx+bdsu1QokHG+O/9OpiQVNWAFTn4COY+kF4ZllfsO
gd2jd+ral4fNPkbne/za3KYSalUKQCBifxscePqSLroxFGzKpFAXPuM/c9GpfAlf8PlE8y3fBUxV
hzpWz/h0g6L1RSabeb9DOEP2ovBHFLAXHl9cLksmwZeKau9PYVqNmifPBNf06ykx158Vu8zB5I+i
OXk0Mfxvh0vMszSzYVXWMC9zH/TKrUCadqTucRxR89NtM6+xAgb66Bhk2Ffw4ALBJN2272HiwFTy
qFKTjH+HkI6VeJzbQjm51mzNQab6JIUEbEN6ihXRAYGyKopyoQfR4HXUl6oppTiMSCHfm3GoMgBp
f9VxYyDTS5W5yC49iFe1pKVBdHbDdDYBP5/R1bqNexbyt7NGsFEI+Wo0oox/45XCbVHvceiHTFXX
4gYGXFOS7Tf9hK9xHz0DvVWRKwHohOCRkJcuw5VI+McI/kDQOzjWMCxSK23NaiY6c0Q/j29171oc
gAJFaa6h8GgR6vKav1pIlhStY+m2ma0yo+n4MUsru7uI+afoRTUpLKYy10aqAmmjTVzQtyGk18ZY
nMwRUZZ4IG9q+EVMysK85DCdigeD/SgpYIL8/4VXIbITfBCBHSfWO013ajvCp4GcyxXnChbP2d1n
9ptQcGizl6Ra/nRPAtQ8GCj2VA7hLymAV2CL7b5BbivZ7Qq+thn8eIoI0TvvtZLuJkWOU9maWHDD
HPRUX+3LQ+IM3vij+rROjDdhON9SnjN2kl0q6gDy9uixr2xOclAAbiit2gKbOKQ+nr77E71QSCuO
n7tY793ZnIFNUfq1dYZ7RZ6AmlRZheTDbyIr5Vfkbu6XRLfCcASUZJwDaGtmbHx85pEywxUiTuTQ
Vm7rkbjZ5hIcFQI6yGv/8t8h2fizyple/QlOLmcl4jSTiqZt6IEZQokR0XkOmWXBWLylPGj/rgVw
/WkD3CALRC+c3ywdDyjGs/wVccKWcT2B77pNX3b24TLp0GLpA9Uop00Nj9NNYTVEZQ//4h37cfBE
fTuF8nsNRRwgiSIKKONXGmpqk0bSmOLeLw/jcqTH7OMIHgNIYsU1864RXlWvFAIsweihFd6Ymy97
yIxOreoDUObmfFA99VpXBDoFooYw8OEGCKw3/qpZp3ABwdfFKZghh7oLVxdV+TV4ephE8/gYr+PU
KeSllsFY33Uv1sgdxBD2ygGjcxA9wPXK6DTESGJBdJFH/zw6YQeG73frfwqy4wcyVJV+xeYxVwoU
JL+ijIYmt+sXF5McHYik/t/QJHItpfJVzZ7A69Yfk2CC01Clnmd7J8RW0de/MPlryVaS5Aob6sJY
aa7W8DNt8b3yjhsSNV2/GIpNZHxaFh20P3dgszrPuTARXW3nE4ZRLUYEhcBJcptqLB4/QKxT3EAi
gXBZ0GWzSuonWWX4rG9ECoDzqRT5RuolNLvVM1WcgXbmHno3T6wuFXmOL4zC2WnRJSZRDBdTYIXI
Ne0YGeCygAHw5t7wshu7ZrgoOeoiDMzuc/KhPjBzNeG52yZg2bDjY+d7+tsRYUFJ+gO8FEx4GJqf
XINJXLqov+A9CBzDkSfrwBGSzLh7mwF2n01Vyv24+atw9Oq6duhWmjPQAVf8X99gRAHQebeXsQvD
T/7W07Wjoo+xk87rdZl3HHUciTtO3Unc+C1vei7x+PqGvV1o7qHNJBOzqaFXILfrmiXSKrwMxbTB
KMB4nswvnZ0H5VlRZRdKcfGppUyztifBCRJAMLCIhpoxJxem6VAyi6m7kxOoxBRCc+1CjItvKJnl
/z1jmzt1gVBHpEb4ULpN96PjRxRO9SexIJw16ncKO69SpmS2cGcSG/i4DANH1v1UlNXWx8O6Yr9i
Uon/zUEsCCiE7EXSob3voAWCxIZTqxRceoYbYU3W0MDOv29WPCV7l3gzWOlP2dbj/Jl8F1edTLNC
3AH0oTHMazfBj55zog4xG0Jh0PG8QKD2BsNTJYh+RbRqgtIHhR+bVI12tSuFbyxwOMO3bkk43CRM
BU7aI86cZ4a2jZ5TzDLiW863emoGPeG4YDbx1SsJ0g9mWmkoqz6s9NW6Fgb41vP9wufRauPK5vMq
A6Tz5wA7Ja9GUHkFcgTHJmgIEgzszFa/aOnizliA+p/8x6sySpmfK5N82OP7UGme3RNAqIk7gYJS
vrhX4SpEbY0gQpWecbsYE6SEy+ck0qa6867fIACOpKRt3EJWhkySXH04svV3RH7r2AG4M7jIub+1
x84TKTprTOFKdCei7NNM8dnQj0lBcaiwCu63dI6O78EtEEC4ZjBKT2PY4BQKgWC994dzVD/9uK63
8kf8i9wZRrJwLhVi8CimLtfDapfDQjy1jcFQcf1ifwg5ewe1DXLjAlpuAu66zZqgPhzY69zQiKkm
kK5X0CcoNxPUxzSTsYhU3yKz3Pp7Ytm/5NjAGu+vuTaFeYGiOUOGzD+ubVYZSxNg/e7bivEYOS4G
wq1hR2wkHFE0e6QyTpKs5aZ1PgJG6y4gNv5CfqdVNMsBBOm6CilvR0SJDo71/OGc2TSjJtveCT21
Gy6z8ZN0dHW/QCsgK09EdIgsVpIggauF8U0faAJ8fyO1HJvAGZvusiLxT51xMuGmv/9Dhb55hwyI
Y/VtZEXpSLpYPeqt/q+BAwDTRDSKV2DF9kdsXAQEq9VHdGUB68gQblEJ0ERfUd9oym/kYX+RPVwQ
eAaI8Cg3Aj+ITxGevtbGXlNXWyDRFC9wobe9mdhgws7fsG36Ovj5J/mhVAgjTIfCjsoJ5km0QgDk
eR+yleli8RXFZvK2MqAX1g6b7+neBGxmcDZTYZTHdh787184/+p78oKM2U90PCFBXPmX1K8PKwBq
uqnIbck08BkGks5S0w0R6O9sMe8nZUqUmSEqCSEcu+doodFf8HeR98maXEFyoaeqg6WLF5/bcDkB
FK4EEgKEu6Qs1IoqaWBD2+XX0MKj7UHAz+WRCJTteRGPM+eGlslBhgDG3F46RPZHy73Bw+G1cr8R
kPBg9AgbGLo77FDhoyAfBAxQr2QPFdlOTDAUGT6SqEqDMZDcVELnwKhLPFeGcVN7hwurILDtvLOR
S33N8IqmDfwCeCRY4OoJv4n+zPyTKzGEovXociX7V+TCnOBjTSb/h2MELZ521eS0fbDH3d0KlTtC
E7pamyf4MX6tdhYlUTdss/AaIolZd3ETGHtVYYFFMdxq8ocDHYlVaeQXx/FW6lfVfCa9HHYWhLqx
1+ccfr9fwrAu71z1z+EV13pHxQ8z0EoFomtes1PJrBgxPtlzDATQUnxMhQaZDdzSyX65bGOThZcz
tKDrLLjH2xivi004ZhgzmRAKD/uGQKguYm9nHcykYYBTavqZTWsIqmy7czkY4S2v40HG5W6Ghw7R
XvFnil5C5i1sJ954rO6etZLI/o/YKbyzU+STdrrDxymVlhQcA9ErVjQQApYM7zpr7IP1NmzybF4t
qDhGYLIPi/O4LFn9BuBax+Lascz8QW3+mFAs6fPCiWY8X5V4E9iV6XRZTEw2dxGQpvknTiStkKYA
kigz5Td6A60Wy7DQLrBYeDMy6HwYE7b+We3Ctc40CHU3bJcpHbPDSAWPAvVbOGbBWEoqjsD3cq6o
LoHsyh3hUCy3Tv0w+kdnw1509Wc/siYuZiVe/8e7UHc9YLTQjC7KDUbKjPpSbm5dqhdOxLxysY/E
KwPOcLPHPtQD2i8C3+5WYD9uwW2W2fmtvN2Z2+M+QZfOrXMZ+ra4TDiZfaFOLPi3xpTRGFPVbB81
f8wnIDKU2Y8OAmz16wfWEyoo9G3uTR8tMk3gV++RhUs24ST348deuJt5niXndPwNDhwHuAGoDC7L
EHlWMhihorEdWgUZ1dlTgrOmyRQqkFhkBKUytV1aMHj2ryPP0snLkz0HeWWstYs1v7VKiZwTE/89
HPtLXe4gNhgoPMtka8nMSlXrukJf8OCK1YTU8ZIOlxQ5D7VLNjCb7zH/4XK3rZQxg5sNKemS/I5C
4POTVXyuTOqomq2lVkarHamUzHGBDK1SGb45cMKrJlYRXbC/BYZIdHivVSh1gbmiAFoeUdiXKbj7
UOWDDsyt8ZFLd7DSVObaZ7jGiWmvPcLV1CXjhLuCTIcVA+nn3QI7tjaN8mdP2+ftaabmBhgJN+JF
Byv/2U+uERJHTinlnxMhpx2ZcigboFD3060uXDV7yahnXjFAITkYT4FwMBz9e+Y7F4vt5bIjftFl
XYzdC+bVPTF//5cYSQgpDvjgF8OJebZLWCR1wGiuNdyErr015hxy6o9s3691fiUwyvzxTGMgotce
G83flHt7sI9P0aqwg8eZEzmwIiycJQuQVsAdD4i3qh0VKa6iTHcYQslajdje6a/6n4ksDm5ddRgO
AU4+YLgsQLtaUoa27KTk78j801+img8Uz+c1fAXnJ72mqDgohz71XPTl6dIpqZAhEvzcr/qnaBBQ
JanpKOv92VdzLNfJYN1B3INgCD0C+u0wesfeivoVuEH7Az0q3xhhWwKNnwfBChGpLBDrAwpexeXj
2EvIqBGzMnPr5vDlSq2aCbKsr1CwGumeYYFu2iDI56s3NmSZxceFMA+PK2qYwTN+/wSXYFhySREx
z73KduQ1W32azEFV6GAZAafRa88lE+lxnXtUgXHuzAbnfYquusKYT9jH3OXaKf8CNxu1r+zNgnx1
DUXNKMXeatRoTjxfdqUkznrNQ8WpSEYNptCwgOX3p2Lva9O6J68ECaZknzWngsNN1ukhSlwISx0d
2WYPuPPLhzsa1qRvHBK2RoqySpSYP4phwP/RFWHt7q4QAwm9rESu0x5GwLnPvIdUZZpUEPcKec7o
/woLcwtSgiG6ohk/kHkUalREV9E7ur/rxCm9OjcvEEd/TxBQw5GLsUXT/EQgBXSfo1A/lFA4NLb9
+ir4hNy/wUVBvDTuuCL4lcsu2V2IlkrOmJ8Df5BEZLYXG7LJsnK/ge7A49Ax0CYFEqxqnV15OFL8
zmDncgGaXkSspRNWB3YFUtS1zXMfRc6hqUePbaJK8Cc/qflhVuL4E6KSJq44KWAWN2oxtNWvq977
IELzUFHjPqrK2oLBsOxtU2M6t+1mndLRLbHYwuYXRE63vmHdSa21L5oP1r/UuX+nJb069EEoGnj+
Pht0mpCfMLnBZe6hnOLQ1kngl8PVZe8dSYXuUMBbqb8kPmrXAC36wbjyxjf8c00oxmfpuKMQB1Jb
AFk1meQfmP8rJTrW0TVm95sAImmAtBzuKg5hIynWxqVKC9Oye8Uv0u8Bls5wP8A+d9Kfyi4ZCWTO
fQLgYSVHzxts7eLfgIf6igrZ7tyKH2JThzbfqmxs6X3qdLjxJiApP2tTHSlY8RhvxHKpJFRqfeNb
MrZuPmiPAo5F1k8/b1qMN9bvRirJk4wTjyidpFSBXLVbounMXwOFhobU0y+rQIEaAqpHMO6cYBFY
LjPKvX6OJolrc5lD1FLKLUpxc9d096aICC5CuSD0T7ic3hnChXT2BZzHsQ8uDR7y8NHPbrWQVCW/
2dVzC8nLQzCKXdDtyzq9t2GV4Py5ok75jtgRvJv8KXIsOdnRNsi3ceofJEQCwBIicay1jMYfttq8
08tt3Ihl78AjRmosYS8Z4Hoft39/Q2T6NMLQyTuN+8hCe2noihY6Yf+zWFpniUZ8gDbTPYQ9w8hS
x278l38gP+vd4o7/l7D0phoZj7djyOrT9fnOrNd6QFc+BKrogAeZvUXW8L5Kgukv7TW311SUALDc
/Uu9Y/i6t+bfb+iDYzUwgWuvAIdg7JCkrss+R+6cXspW0AdyeA6oBgqgZmTKJpRtv52LTTqedENb
OqAQBRGeMNvcgTaHSHOEs6H4pWx2OGfZDhsLbedo5yjiyzw1PMMjNw7/T6Km2Z9pZcHwh8xtbi8K
StYecUVjnjNVVLUSHMcUIg8USDQUEAU9WRiwqaMfcbJBbqy2kQmiztD7758JTm8jAeYm0awp03F8
OaXDRlnJ+RJHVetqm1fPeeXuRuZ+AXZx6DRcOfd2WJan7wau0VhKY7C7MoWG5frMs1VfFDM8r5A9
i7G2iAWKtb0b/k4/X3cKCYbi6Z9NuPol1ucx851kT+f7gj5Jz+cIyrWZWedeqVPQowW4D/YP+q9k
QJJUfkWEmIOgrnl6ClkGE7ByHxn8yVEjRN4VAkxkNjP2diL0zW5cBoaApOnkIo739rV/gST+SXTz
l1jmde1mdHhPrNfJoIOd9Ca8IVU/Ch0Ho5W3QL69JalZjRx6VN9GNWrjeo6Xst7HXHVefIyJB3rv
6Sdg9I+Sp2wpIDXwEsQ2yuOtkGRAhrEGdAuWvcwNlnZ6sFSx+muUvXl25vS3VYvgMVMWFv6D2aY/
f3AaYo0UXFecJny0jmR+XPZGRA8qJdQy2be8HG/xFtuQoLa8u/QZXd0H/wOAF5EGTH2I1P35b3jT
NR0hEfPbrwvG8NwIlvLx7ChHjOb+wfXNCwliHi17U4KH8kBJe8JiVVT075QcIXQmYzCmitynYWXa
hnDwI8ZNGTvm+ABSRPVhmrPXTOGKUi2VtQ7eUVl2Gm6kN4GOEfcUhVBac9LvgLsQfgalRlj7ps8b
8H2MO7Mai6enZ2vNjEuzM05Z7SRfeqYcaiLJaYrL7uhNWCYO5ZOYINv8mm1TXlb+s0h4pnx9jwS+
oafbEOfWO50RsqyD9CSbnfyPQtrHKbgYJqFyC1mta4JMUmZvHc2a/w1WDEA2uMC9uAwk9l0VRIaH
0w5pcTW1WCVzS70bMUETOmCRcY2CUe6AS+DntTn30CPSoSRAeCx4KqRMbWvqh7xyLi092SF5F2Qa
i15Ai/NPQzY0fjhkNHi1OrHiPzWuR2EmKHNYY/q6zumuLz2XrlslRzB0AJk1BasKClFkLsnVfvCU
Xuk64a4IYIErnzeUg4Ytu121H7qL7HpDGgFjGFzgIB573aP8YD1leJovxoIXrY9nB6vgJ2MrUPSn
ncD3ysB+2CCY41oDidsIdgmNjeJ9shNvWIMadNps3bnP/xE5B69KPxBgi++7KqKa56SBkhOxkvkh
pvTtwI6LjS39jFFqbK4BFAzFw+FUUgZFQFPARpoiju1E/sBz826IIhJg3cprn61YLgWvw+jH21i4
cEcCXfniuTVJM0Y2Gc4ZeZlvl1CoZxMhWpxUDFzx7vG/lhSz9vbJ9v/TCox/vLBwxXRbkaUV3C/v
uP5887KuSkInPPcQrSMRjloa4rp3+PrP65MxV4omAQTaiNkO2MOb0Edu29Mvj3Y2J6C1tMoI2/sK
WXYXotJ50nPlVXN4+SrEJEdP/lmfh1uOJY80IqTSedazq62ubwwgjmgeWIYgwQFkViX9IlRKA9Eq
/7pNdjpHFo0qw0L+sU1MGdI+f9Ca/QdVgJhdOGpagr37gUN02dNUFwqwKVQ+B8qGXEALXOlSJlKy
TLx8UY1mq1PdZugRQkJ4btBRY5B6Jg3WT8K73wgv7YN5lLgcFE1WJGuCQgtgANv40vUsQC27JvvP
QNayK+4JA3wGFwWAZ0FFCDHGu+wE9IMx98vnVV4uOlV8YLypyqi+mSKGl0a5QBQZIeQK92+0n4a7
azeGhohC3Gj1ZvFfq4wNDIkrrs/k6kSKvuARZOHktzZ5B8NwDone445UdvEqJxSQyu+LsNHChr/C
Cz4RXwrfCxLzPmWR06OuO4meGyaH/Ct8o3IiF8sFEQrBUdymoXgrYilaNzHsd1EMEKikMZ0bdGwy
xwqpRlJGOrVi9MteBRhzBGF4Eao4IosxqOe3SRTaa682CtsBwh5cM5NXTuxEtdpPjp7MDNkIEGmX
Vf9hZJEvEGtk0kVkLr8v7dFfFDCsYWsXpK+cXZoc2oP0SSq6tscHDHtAigZpUKzKSk5b7D/feAU1
QW8uzhB21G7+jbbGpeFswdv0+WVwIWDTV7yHvcKjaIuTaPOp/LuQZSAwt7dY5vRn6Fq9ait+GNPW
32sam3rSd3Zheji5vs11KGhLc2/d/ASVbDiaFYtXNSi2jJ0Zp7R3CPBSCSntLGLCTju4leuHFxn0
8Um4869HSUGTvEhnbIHE0DCXWw2Z8Agx92yKiiTTJeGc8GYgGffzuG2YBvI6INtMdrri8RkbBLpq
JCqPEf8o/2WBARA9B6L/8unldeELS081R0MdjVfFER+hCv7jNENf2aW2q+ot4edzrXIzh1ehi2qz
D7/SbipBiq8Bs4mIDFg7jQwVZnx3cQpjo9f7spCybwOxQbOByn74vzCUGYYRD3Ixy7hGtYUfgTvW
hTkIQlEVol9Vz3B0knEQqeRfbGpg9YedPTpuNudSq1rE1b68v7C+JNL/QbiMhryDzii5zHVb+qvN
GEhU9ZkVWqHPDoQH2cbQjwjpUAOBtZnneVK7zpd9a26S5zzxQSGVzXOighzlytFf/xFOaIh5/kVd
+6/8laJoBPN35NHQvXBYWtMsaOgz9eHN3hTecJekGY4789mCGoKFytNeF4nV1/Dir/Wt/gmFjQBp
dmB3PfJpJYjOkZAaQ+GCSec8mTET8P43rv3otwEgJv2wU/O68LnW9g6IqGYUIJSfxszpKhQOLyiQ
mw+ODTTjjGNq9tP9coGgLr6a3/wmPNAOg+5pWg6LEwTEXwi9zh+CiEj1ZOB87Uzin5Hd4vOg77gG
dU+67KDV/gBfBtDMIld+PN81ZAKQRnYfHXv+GRZ42caaiJ3DRDyRE1OuuAuR9cV03O10OeyuXbMb
DWKw4zcbcqStnzwj96YDXkbFFxjZACgvRRgugtfIjjLyNJXuEoASjpmNYp6jjU+c7G30gOTt92/C
tWLZGfMOC2gQ2QPeF0Yau+f0ffe3nPhxbFcIFY5vqAnQB3FWL700FkzZLRzzVI5k2C49Lz8Va2U4
4nAKV4aQjIOKC5MQC+0S2FCK3WrNlV1wxUNOb6hkvasm3JO3UkYSzorjeRgyj0cI1weOMUyVbqDJ
0JQw3fAgnHcg9GdbiA+mmEsd0iJhCM34PI5z30u6Aez3NWrWdPiOZIGFHO+vaf5960JbViJaXNiK
AeneLi8KX6CWaROpZIy46qUB2uTysurpIqBq/uDh4Xo6QbqpqOqoKGaXO971qsRaZat+CREvJxgK
n7xqpvVSSK5BIg8mcGwJl+02G35VjXugJO4JX1uIUXXm+VYo0i3dRVYmrcfSPRAtitGNAllPzlqp
ORwecU9wqdNTgDnH3tS7DISJQOPhmGMs/P1al1rr9ZnuJN4oTUlCHw4PdvWzHL7q7lsTJdHI8dXJ
qCg/4I+IaFjkqdapLVn5aTi5tQPgbUtHAqlLt1EmOBFgyUqr0gWHor03Tq/e66lNwftAX+5WeTlS
hcw0tFvhE5ypTulJDgnx6XP5oFDSwSckCoJqp+2zYYzhaxBXa9debPmLp8Yu5nbKDOjwOuLLdlQB
oniZb5Zox650cEp0DU2VzDDpmS+aq8XMw/SC34E9y6NlgjiYvB1EzNOtPquKd5DhfHPphfoJ5EZU
Nu0LDpuaTjY3vMi+B61ZKyPN4O6kj9IStK+UIY5L5TSX3wMRaK7xCZYLyJHkUkJQWHl7VGpQvGbD
5INlde4WeBoYcR5txYWsozfUmJeirj6uvKgxJhgxoqIKREVeGChD4x9oKqys2y8gYtOFjYSaOz7P
zYOwtqWRjf8r4Q6dWwkTDt5SUzsSRQSl0Md7cz3dQJJVw5PhmqVZGAjlG/96Z/BgsdGHFZ8MAIFG
Uo8dOzIZUqEQ74cJ9HtwHGTpC/zZLM/3yhvhawmMOgP23thdDWbuDSfyU+mTKpEkVkdhuwYkZkBT
uMK5JIQap7fCIJyNczPL/QmrwDPpJuNoGv8r8rrYZhqBngtrAVep83ILaa1rba3whlQUm2TR4Pkg
NOsulm7kdnBIp5ndeWRFHv4y/Dk+7g+EtXJ17UmPGM3gB440G5lnl7ePb9utCHRV3dkwotbaJQlZ
KeMnCBBQsLAwr0+mEDCA3n2FITp4OQvJpSPZul/StnsuGhzYSJn8VTt/tiGExzczZCg9fJll/ZJh
VL3xBkiL5GE7t4IYHyB3sbKAFvPNtXPmG2VcDskHTlNzyDee/wx0rqIuk0wsW9+0cm3H/1AQnqPA
j7SnYqnDVelySv0rJ5wsGPkIn0sbof5HrtJPjQva3vY03vrfDyuwj5kIe6WCP/7dkt888Z2FG/kJ
4o5oCN1DHtPHqcvFNTkIEkoLbyEoh0JWAAJ4/HxiHCdW2etgEiqmw8YyoaY8rmtl2E8qJF5yQwG9
Ui43LJoFB18lIlyVmDUzL16mZnRO4C1Xdmi2O2OF4umSDqfImxv1gSWB8HlfjB9eUJaYJl0Uz4z2
OmNw0CHlFcqO5tIgX9jbNnefe4naYOJEH0jJ164dLGGffnVlgoZ50g/CY+6LgZABkMLHUVyefJ/l
ZuDjzJCmUDYt9dLJcqaZCFh6EXVv730d2hRQBE5lQlZ8tanAoEnscBD4WlsIemySka3UcptjwzFZ
/fh0/5sHNaCgnG2j8XDVfpzt0G3gr8mTtFBgrYVMpYX5iffkUK50f+OwCcUgoDSxpbBWwyYVDyb3
uOv4iOm6Az4TRMKlaV/yGQ9pyzpqiS15pb+pfVyNVF3cU4aOh88vOqdfDexZHPK9DnXwbyHCclZw
k/7eZEpSZOyJXwRW3oNm4LhljHkwnWuHxhgiScn9rg+M+Me6S6U2VWGSUUQ4lCUUI6sY7B9Vb9sk
6lxO9yCiDizJZrA/HiZ/lnX9172sFBcuOHdFEiZcYA05YnSO3fVwdPZrrl6lReAghW6aEqFTX7oi
3nVyd1OC8/rGH5KuitvzoBCdYrbuQqTZTCEpqb1gZCnPQsurHdW8TlS9fK+ZGRHTP76Z4zXtummz
ybmBPP1lwHAcQToj/+1I4S1q+KaS2PYa5Oe7XA/5F0pI5d6YNYt1hzzcyUGW6pKZ+tQPMGl2NUsN
WqhIAnBEV6UthSBiFofd1LAqFXW4cK+jPdrJtKWq0sdx8lsS3EuQhQu52sWVs49xX19R4UDIhSkb
aA/tJxtnRE73+lVCMK/HCRz6Q53q+qOgs4YpCJul11azIkEToLvEH0NIJ0xXhrnIsPvhE7ZB7Jf8
9P4ZUCjexJVE6mYezYULCgqWTClbnWkGuXU9+sb0qd7ymu2NlUT4fyvxIb5RvQ4mgklBix+gXXVD
tarTBh4IvkZGpFFxwf5pQibuHPQ0Z1x1TWiQyZk/HraYMs8Vc04EDYWVhXge5zcRK9/9rZkeyhRw
88oBXv6cpVqK2zajcgh89KMjUtdtc9lUvBsjyDaGmKak7Knk1QqW8EeZklsN6BrwTVd4RAFNuGyW
9fDtGEG2NAH2XldzUbXCxzUXl5QbCoSY1vdJuh57xPT9G42CjlOhMLOzsSwLOYzSf8ZoaAr/lPlo
rGIIP4dx0qRVf9GlONYrOXQF+nrdHOahj4sKhcKj0314NbJzpGzdl1UcrKTltoWK12pbm04uTkBK
kNmxTk+/BVcsYxoTjWyrRcmruuPXj73rT4rYm8o6ATHqidgMxN3Ex/LWFVVd/tTAHT8MUCYrxDyY
S+htwiOQJAXOgTuka0HcsicOqSgOx60x6CsWRlzCLwksg5m7bv6Q7L8XAk/degk3I/Aau0ZBRmXa
hl65J43OM5gC6+sYgosuqOrx46VwfruseLHcfjj2yYULstQ+ZIC7CAKZhWHASqxhgkU0C2JNiFfm
k51E3B4NInpXh4cBVYq7uryqT+fjRMbBQVYLDXShcVPWjtcgXfV2xlJUc0d5y+uiBaOBM+KN9hTd
XFyf9Kz/erBZltWbo8iOU34getKPYJHJlWbV/avBP+MxstvnmPUujvgrMer2+L/5smwbe+jKVzuG
zjD/Kk6EfhveBAUgu7Y4rgU9nrnSzaNXDNlHXykyad9sYJMYdlofhldRZ51mbVWDWYFDBJjorREW
FfX1p9trafw7PKFygcQBxN4jhq/8v4diAArhH01L5vAiJntdV4MxOPymhUS2T39ZztAwlmiyIoOR
5qWngGaSzja0mlm7HmeF9Dm9ziHYU1x+VzLgS60+VF7w9WSByT8g68EmWPtizGi++XSo/Aos7AvK
5XTksqPeBNU11hAd1husP+zdED4NQ3H3SbR726XWto7dEV2MsxCG4OpUMz9h5QfjbJWVsE8zT1bl
9Di3Sk7rejWZyNbGiX/alqAPWxvRSksriQu1L1OYTpZ9yu1orq/ebEWVKD4UZpnBWT5ss02lEDdc
WsptHVw7DIo3AvzcytwJy+XBkrESRsAjI+uJuijh+4VC8ifKqQ6gKvJ16/QboMTxgXVmVPn7OEJF
cDYksouFWVCZyukTvSpd2xXGkE2frlXu4MpseAVABXmOSncoxC+C8BvaV8c7Uq1j0gUN/w1Lf3g9
MKMV+iFLDxKAMk+BSzM00t89ZTUb72lyLs3zN6u69942dzpYukCB6LCq4jI26s7ryEwJSv5g1N6o
DxUiEmcMJoHeTbStMQtE5GjPqQ8jrT2xxYHOdHeaMpGtGEtd26OsW+26Q4TwpUulpxLbfdqHFIx2
kT/Gqo/3rKziifb6yaVYJ0PIuG11Ghcns+bzL2W22Xgks+6S8SDSQEnJd2Il40mpUx//uM/h77Qb
fnMe25K5T5UCT45h4PcyMjZQtJuDJDQD/PimUFttNGahQdFEw+Pv2M77JUjC41OP4UKZjzuJ+LLI
4XZkck5UsHvQEe4ZjNmgGPTahcKcG+5Q9onBGgaKj7gv7qd6CAlDCjLsfy/ylyNBsnK8A9FWka3p
ff2pxMTrb0Nr4twOiex4Mtyvr34ZkNwa3zNi14pAMzhQDXx0jWyX30hN4R7q0AppHXS2OLChwZjF
4CaNIQ9pbclUhu7Ee+Jzgk2FxCygyLdznfcj3JqhyrwLKjRDG/Uo8E/jdiulJmq14+KoS+TG9qj6
WMDGRVvkrCuiA2TXKrHhZw3aWgT6IcPMaC/XQVmEJB1kwrQYaO7BQF5M95qFV5XGThnX1VvmnQjI
sjRevh4JHjHo8akwRu+AA74Jcilmh/NsTFUvTboQbhmLZ/3eFA72Z9AtmMpkRDa11/gVrC5q2VYw
/jU13Id0MZf4iJD6fvVAACfvqD9v8z5I1su/OtGR2LNFsY2mzBFqGN1kiP8+JJTavRzSbfK9bIWA
I4eBoeFF/J+8DNfLBeXYC+LTWzArDMIj9JrqIdYflceWQPMGC2KJALzAa7nFWwypnDWPudyBhZHa
HJBn8eTp8nThhqN2h5HFAG7r97v+lYqIvTLSrapkjFqBwM3VFU2p83oOE2b/KIc2mwU3cMy2Nau5
GziU8dDoFGxH9C9tXpDpX/dPVJHz2dZtcLoLEBJ8K0SFVcfZBNYNXewD9VqVpppzh0ZsC1EBiUR7
0CqQcY9wAVuU/Gqzk2FeyRdLVqvs+DJMUwWY5odgrfGyzqfMv5ruGkhY/PUWUb4Zs0Dr7GPIJjIR
dT3w4KICWdOT0h527Due0nacQNNkZOUsFrNoDQB4S3VOBmPT0OacZiiKK6zPmJJkgLIB9TMxm0iS
/IKZk5ifIlaT5tQXNf++HNmMaBT7Nsx4HOZCsUVyseEgCWcvjTI26SXStqsWVgjyT+jxBx3nK3b3
/Cf8U22m7pTQ9+8uE1SNz7rv07c6pRdiSNILu8G7QgeiKl2K1ypQ8t1C4IkWCXogEHeAQIZZrNZO
3Kfg36TT1AI8NJLdGW1bCpKd0RFyHJpe9hZ324em1/Waef0vwHbRhlalS+BJa7yXyBttaHQru1QI
gCW6CeStQiJgdqlSCNCCSfa9N4LMOGDrnGxFjg6OJoA0UwqycIxjqEbz12rTyi6MBOiXJLZ4pPij
V//XesF2RTJguIbUvEFyjMK81bMYaLmymSHANi9Ta/aS4HpprBqhBA+jIADCExkPhzpg202CvbNI
jqSq3sHQkrAIiDppi0Km8nlk0yRYck2eENHBbiTo7TAeyi6X6DAHC9lmC9UBru1TNRjY6lNmTFHI
dalk9eZHUj7xGZKJJ7NW6jM1VDf/cAQJkatEWUjaYElrsNWyKMywyNYNR0eSZ7GNn0rSFvMJVLXM
noVzDYE9e1dqNtt24erhp8B64bFtpmPGLS4godXJ9RPZqZk+W+jvy6xwjDeLaVCdhQyHRPsLUjkJ
yV41ec+aZtfP6BOA8nf2OLoRG+91onbSvI5coOUFwtTxP/Ubo/7ib4tuNhyBp7f82AO7S4z1hRCH
+KeJ2ROetndiRwK0/UmpZkxjLVvwuKPwuOCgfDYoc0e5sVFo1p7c8O0CzWhFeV25qcX89NOfOFi6
xeCosfU91wgVC/7KqUBpN2Hkex9idoMDAIIxGB50LX+mLlrBv1AKQFuDceEUIwYGhspzNKtLNspP
zGH9ZUIouXBlTrP1zxocQEaTo6fStBjSeW+MFFcATOmi+L5MgLzDiJfc2Rt7V8e+Mk17A6jHg8kW
VzhsIX5OLnzXcrPLSZGIqh13p0Y3WsTNWBw/HvMCY5HIT/1I2d2zBwQYi6Cm1cM2ucs6E0zfGhWX
OM0GRryl/dviSZOImMzULG912RMmaLX2axsU3+n3fp8xM/+F28LgQy1ZvAcIOQK8LIZh0f/7Vn/S
ajeUVLH81AMIgmfeWTG9KkBICJ/ctAcfoHyTLqyOAPKsc040wKjoOBS36M0fDZ4pQ9AbVDGfYwyf
4ITAN85hgeAchmx7aPF8+hWPGaa9AvKF2QQrFytR780EFD2HniWgT4vz6hicgU6oRhq4UALi9EDQ
VGnzYjI6iXUaC6/j1LcsZvt7BtxK6VNE4P0VXd6l+/MV1iCYadc/F7VpoRrBdZTk8CqOd4OVoQDB
xqfr/KUBgqh1snF6J7x52oAvKV4k/huLnXVFS3ek3OUfOGOnGqehNqVcuC8dNNAqFSHG4xsdwJd6
As4fCqxTzjFYsW9TwxzGAknH8R6ioy+pOXuEr22axv2BTdSBXrYNcltT16F88TXX+mc6tpVAp5iN
G+wVLVjPv3SH9xDm5UCMzxwMxk0/Nl9Cbsg1ZNu9VePWmCUT1Bq31ZiUDGxZv9pMZjKxK+do2fbA
jfzGn5RHVdutdD6IqpdbEGYARP8ENdCHBEv7LFI+thACIykGqG4RHmTsF5bvEcaECb8UFRDpBKJC
8CECebcU7Qb3Kw/DwC38WROjCmuF4uwZNBz70VJGRg+7G2t9wcFArH4A8ghH/ZaFXxvYBINvIEjP
nsH6Yj/KnlZRY/apcWJyv7sI06IsgOIJBBGigXniJjMe3B8J+ZzQkXC9nnlL4zX3i4qirA3mhdlW
0AKURBqalntUT3UChvoAeHjy70gzMtAt9vksjRCFcawUXn9IIO0avN/PEjpbB9KUMjXlvHAaCh/a
pgoOI8kef94/N/PH6D4EWdLwnWJUgzNWQtYMYr59AqCdF9xMmlCkW4m3gZSBhL3+bIu9iUFurRqF
GQyS5IfzT6tESm994wUPQHAguUpNWKHvzy/tGn4Q/V+Nyjil6r7oaoWpE4WjrQD3XasSzQCRg5cN
IpQErV+pB0DDDHXDxL0ha6RRMthO3LBuG9GBjOMMRTOWtdz2fs5KwdxxFQPyRqZ+W8X3ICmHdy8G
yidq2s/U/Ejz45pUCxgCOFss53f52ZGrdE1GlJRJSSnvUUzSP3ucEo2fE+7EGXxhmNy88PJ0Wzsw
neQsdD6+RJC0spgc4cCdYBcXdRl/oPf6ZDZQ730gVM9aSqmI/o9RElrgf0dXMSXvZ60brdQSLb1b
q6a3h2rhTpmGp73rIzXAiEgHppHiRHvpfVTP1VB69GB2TH5LJ1NQdKN4o9Ht1TBhTGgoFG/IW5C0
VyINlJBDPFU+xZ1dhZ0HlkxepX1YeTVHasq3cZ4WfW8G/xK3zgfP97HeZdk5UrMeJELB4EdbAgW6
AFnicH+4/K3EiS+3Ue3jEMjewrRpxTCjYBK90vfZYFCU8ElZ7P3E1bRr64X385kKT8VBBKbt+MAE
yvsTtY2iwS1XX55od8g7ETVYchjMqAF1CGM/al4Dmqg62MXX0R4j/qVSY+7hTKMytRXeZ+jidNm1
CMzJ61id60z9dM2rw50ogzinO6bHi8IhqybMDOQMg+X11cNJO10gSVpAO1mX3vOjr75tfPWJZHh6
Sd2Hy+5XF6q3hXE/hnuorgqxKck4msD6a/+ybOhcvnykeitlalooecEAEo74/DYTmYMXOnCcfL4W
rASAwOYpLlApMrqUVnyMMzNPb3W0DWxwOeD+r9PbySFaD8m1IH2rQeEWkd9s5Fqmog2hWPo7To3x
rrd5njfo/5E4vYV2Ex5r+fwOUTMdI9yllDeomKDVTGwHqS4/MnQgP+9Bn4x+p/+y/TVCe6VGnOQf
408BBLwqyteSal7nRllJ+Wlw17wr3yb9n637bR1tPpbsFFdYVrCuJK8W3IXnhYQexDk4oO4MUu0x
9Tl2BjsUM0QpuxJeTBohHi0fWyc9PH0LnmkBV8nZOieGhM5+kygrgV/ecjkkxv9ZOt4ch+wz4x7z
yBjcRs3xhY8pm18pD4xkDGz22vN/omdaxS5euaftWVAnTLIlMjvhsy04MgMsRxZ5XwYzi/qouv6H
3cGskb/x0wbmKk5uQQs68FKZTtf6VN8XFqjELtAr5izQhuZ+Ski8xews7m8OtnvueEmeFUONusrP
CEYE2tC7WopxOwGexXUGEuDxanteyhT+7wDD5237kK7vXTKQXGkqyYWL40PPKGNBg6oXbsBSaOvd
D+SIf6L5XMzVV8WEd71oZYu3Xv9Yk6nD5PwDeomYy4CatoZRDsv2bFi9cVvhPzSHgEbTnn8aGm9E
12hcw4dJcePaN2tNP2zxaqPgPZ0nohtUKYezbCs8pZGU9IN7QM/qv2Qk6CGknYo6B3qz92tFUhSq
Fy5YxHi2V2N2O79BIG1ZYLUUOBXk8zGv/lroa0AE3BMukyUIXEgimP8DL/X6Of/7AHzHXRE0sdbl
hV70U9ENUex3UlW11DDIJX3W+GJ65ssMxDVjCLCQB2jmoHuEH1QJHhrhDJwumh1doAPnSkVqxBUb
XaUzIGErZK6lrtSORNmUByOh7WddpZvn5+XYeFVC2gUmW/hCi0yKqQh9JbV4Gxtm48+B0QrV1vQz
gupSb4bQsMUduFIjUuQVgQSJebSD4xPh18bqd6GXI6C2pVaSFASHNdAGKl4z7lk4uw6a4mtB7a7f
S6dRPNbYeLOGd2sdke3G4m5bJ1R01SVfDGNuM18HnAxnjRZg4w8qawaDdR3ma/gaxrpkVteLnYS5
rQPsFUs4Ojbv2B3IJUGNVRTUZayeAo/dA9JIAwUssuvW0nRVgq9zl3TwngqftdjPya5NQUy6pzkn
JD3DvxQzOjaYClkyki98porzWAsBCyMbPQy5O1GKfVko8s8nt3tvMJ9B98a/1FBoUc9smcuG2Ilz
uDi/kIPh9C5S+WmnKyAYThgQUjfPXJVP8Bs+/4orDxK1ndYk5O1Zyh2Y9rpbi+g+IAouiKviavZI
Ba5eLHf4lPvV2BxAxKptNZeOJ45Lv2oDPk19kg+D1T/p6DETkbHNJVPHLDpwK/F1lKOJn8cNjbae
LQziHB6FmjIniPDpd+6YaiKl/xBX8D0gegxA29rVB3Fg+/JT6amjjNxskOkmxKTSoDDVzoAgP3pX
0AVAVnWGcA8yN5vbbH/UGc1PdbTK+0BHvSDMOJ6wq5h6KBI/MWP7n/QLZtaCiI8CfDg/s45BIpnB
mOoomIjGgVhE3F94SDuJFOSxb52ja7mLsSpvkpoek4ZImvtfqps49LkN/by1BECLZyz8Fl7BPTwb
wbUNpBjEFq/zCs5SGJuu/n8ZsKO6TN+sMs375xGz/yrvHBzIpwdl1vxVJhSAkGq9iE/j7bbxQJhj
TyRuzLY13JuGJLpKiLR/luF/DD1czfc0cww9TLDUFrNvnQOqKhCQ0LfRnGiYtKvArWjhiT6wvt8n
/WbykLW4N63ZYgAU2eCx48sq8sOKXGedkwrge5My97eMXJYCF+4avSrdlM/aYqieJooWRyyiq9Kd
eXcPZW3qgIgTqFcBWAiAJ3w8YM5s0dEh7IUG1pNWKHbEoXr6lxniOFN4AOIZmbvP2QWuCbL8lzYE
wRvPPF74/ltjj0/aKVm7PU2SjNvM+KnbCXc4olUVATYKU7PKiVlJg+M4w9aQSLLg0IylUMuStjRY
MPpVlEx+zZRG8cVLAMACvZeWM6q7jFmpWYM5+Tw/Uqb6+W01olLKu5F36Ol3BRSxXmaM5A7b5qGN
yf+tr0NKEd05+/N6GbEH9qkn9KAqBuXLs/C0mrgkWycYgVagJC60teCZH9QABpHZs+8COSvroXT8
ykaDIHSZ7hTx757P0gfDSmk6wdmDGzC5bXq6wnuVRndKC9HvLxO9svhM5hCqnQdi751SpWvIcYQ3
qbc/qSBOtdQ121+WQ5KAwn6ogexs9e1XMnb26gjPB2ykWYAeeQIIFKmszCnm8kCMrW+IbDzx5G7L
it8O5vrbUutJWm/f6xLaBeQO6akfMkONlhGRHe/4wLbS8cYeiE7xZDtGlNb7VRaQjGVL9cYpzVbh
XXsYwgJwFR5bt5bRfav9/4xS6tjPPupCPHuvPwrljZp8ELENd5y9qlNJJvlV09gHj1RydHE8/vWn
qyFKntxgVWIpNPMgpvgNjUzXHpAlYFSheOt+eVQKRNQLr7lnLdiTKM+VjOMEnhXnMwvg1hM1zJty
38bB9U+U9zz+4ylRsz8xR3wE3F9Oiy3lwjyaTEEuTsJvJpXPFsuTPi6/4O1X6Gk2jk8CzS7gho8e
xIxQaT1TlagaHPOaTpve/xji/9xwFgUa5Gt5WdqRRSuB8EajECdGOYVuKWUyQ0gbv55ohS4KZ7FE
u7f5AZmIfQo4kU6y9ix/NHGS9g7LLullSai8/LPdmn9A1n0sa9RNi12Bi5ABtCmAzrRWiF3F/nsO
NZOVROEYy7gIKZUDQGTkZ1OsTybEGji5xHDvKvfLEjRq7989s4xrj4XpospZRxdtv3zNCAjdRjIB
n8CMcy8pEH2cGdRbI2vi5twELRKbQ4YxK64Rk57Opxh6LOuJKCYJ6P1pa25q6ZVCKMA0ug1+26gp
dTMgVRwZL8H3JJ1pbTRapTYJD6/qxabqVwkjGOGQq6hsqutXBCAcb4bDvSHXwaKuFn3atHcsFStg
No86fNlTi9s34XKwOLyCB6tUCbuyH5pAXN9v5Yxoqr+Mfbru1RsjB5ZaQ9dz78ZtyX5GFx7gZ1RP
EB6UUqH0YWZP42TnSjnDa5TmBeGj7RL4CTbxfFQVTAWuhedKTcBu8d0Y0RsQwa2w0zGNcOr2bBXp
RxlSueAd7rJ4L7a4EijCrnZoEQP0LzJ7S6Yq0aeiSTJCaeUkLcyBmELzJw5db4nzPYXQgjeQXlD0
RzYBwTkFticK4Fmhe8fh+UjsaEVLT2rvl93peKoC+qh7R2xqzTUmFFpL38Kg7G5txjLMB015Be2k
oLHXzc2ovIZwr9ib6ULrZzOsRPg8cBaV5gFWD2IGeL7eHg82eVS/LQoGcDuOWKX8mUOTcBqoOvnd
F7GgnDyyINxS3vP/+buelNFCtBjwPyw3Rlzy5K4Ht/VI6RvAY+IM74vuLePW+doxynNfVf5Pq0yE
11e/4Ln/cQ/Wi3XweFDg/WeBA1AGcu7jyFgLoM9JzK0BpU53qchvk7TdZCFYnqdFfAWxzBO9niMg
nr83fMpxsZ4nFpCe3czbAkW2M/3KwJONRZsb6iiP5H25PVR2BUJAuuve28CKHrUS65489YR9QgTC
16Ab6En8c5FDCbC7x4SOe3gG/95NmqA2S+VF59MqSkn5xZSYoAbD+Ch/aZmPC7io2dYCNb38Dugo
TaoxUTpsZLDbGrWt9P7RxLOWIkdsU/O3LalMeF96lPWlrYlfcaSFFaa/qnxAFZub+5lkFiDO4bl3
LY7Pm8tgJWzC5ZtyBLCpbAVu4BqmI0eMxUE964zsFKay5q9xlKuf0Pa6qmBZog1hAkN+HTXQrI99
ueTr14bM5EE6ECa3RDYt/3IOy7rHl9iyRGpMD2bq/Yln1b3xObgrVGcVrH90O4JXkXrewvz5nEP0
NoWP8tRxqAHgAAg88zeUUt6jXNxwYYN8sOIZFVa2EPbextwj/4XE3Hy3+14jFvZxaqIF495NJYhC
3LreiI/OlFF45ZeZON7mytmIj1eWZI5Qa0amc3Ck1dQbbGchkdSqXpWVY4CQcMv/J4eh+dAiUhPZ
lUXcci/F4qXJVN2I6tLoIhZtocdWgsRIKX4qbYm+ZYKoRMWHRWTWgI7qnlnAim18Kgar/6ULTcEn
YWaD19HiUfLCHpLaMHkznyfI38KB4Mz9af9tNWF31YwGUs8+ELhpa1NtcR0WECXrsKmseFT2gTXF
K6Zrzoak1EbIcUsQ7rL3XBxUWD6pMHds6rN/8Hg6M1NWkQ4+gVmLAaU67Ih8EQ4ltdAkv5TR83rx
nrAt/TaG7rTz67PkVu6pcy3D2lhJo4dBo+nPq3IzYAgOnZ/S8JHZi7cI6FHr1bGuOIiZkwJQUPSE
1HUornvn/m2a/0klvZuIm+UDUDbUibQPHCkc97Kg4yN8HiAN5uryPcF63MLMXu/kyMphzTsZ8SJM
Knq2erGaIoe28YDJnkvu7fc2zdiUzE4KqgJtVSkU/Jk5LkZmVrCGHH4q3s46Yh0eFi+9XaUNgWZ8
7vv6AEGqt+XwSRg/bPU+oQFUlkedMPborseHzErQwwOsG7MP3jdVcWP9zR6Z9a5rMyWOfAFNDWgH
htgtGJBnQP5KOfC+gM/eixbESiyiyG4i8XcQin63zKvEZIfUy8a4hrKdNiaViQo0+FNorr3VCxVc
1Lp1MwXhMTHl46XnWE8aRgkgryK1KHBCG/GRFd9WRUXXpSfIY87g5mUtk6Ts3yjuz/eWriM/4+AS
bV4Yb4s6GBSt3cSmRjRGqJtLzwiWClPWtjEbAoNrwc8FCGOyaMmwyWJlpCul9Ya6TtzN0LqZI3ah
KluQLkrU8BE9n/mpN1hwr0ZzuNCeQXN+c0Ulk+P9bUjkOucAjOTubu2XhMvWq2Zmx6Q78bsWytxD
1TemhqGYZ+4x+nh2r7jZAaqSnQcFwwTiIIg+ciDCCXbEDlrID1XGY72UseFhFewbL2pDmi9skqax
LIgPNI362jYMLLtRH9VTPWAJ8NkJnbZSmJsFW9e1ObNt5JGiy9zIZzg3LTi+fYbZORN27F3uEIeA
ncFneD9Qg+pWZg9riGRUMoG4bKymFjbKjUmwKL3Evs/+Px7WbtOWsXVTbG8sJtJCwnbdlbIh0mVB
chWwXtCf/W8Jc2ZcJCV38GLCs4Z5a4i1/z+D8LEBan+slWk2S5Bc5PZfDMwt+dKWbKRzmYMvszcM
bf52cj/qtuiqlLdyBcqWTiW5eEsEQ2oK3R90mYo4XhAoPSKT4b+564TqB/lg4s5PT5SE/Wmumxk+
mqb/pHvIjFPde3PYtvwPw/5KfNVFowVx0VjqEjb+OCqgrGy7BzApW2ea2+5vSjCBLjEZ3tza2QYF
zn1z6+ud/EdIEqktcHfl4tBLM9DE3keZlYqpzUFwx6HcnxMB3TfHqbr+HObkm2uyCw5DFlA1NjBG
7kKclcb0cNBHEeHdOZRMakLESiYHTF9vQ8SQNLU9G6tJMIegegqYMpCQ40xUKkIsguMHIzwSiRLv
bvVzBhyn/vMUONUQjxAM7DCnhVizV82XMITqplo9D65RaZrSW7GY6qNqerrSyZPZeurByU4D9f2f
7DCTDDBijl9NX4/AVL4hNzGTn8HKxuivx/d3o3LZul249T1gldwotrZxozKzZ+oOBGD3ZtN2y3XZ
SVbHY+EmVB+usBpC0a4N0sW0qHfymD0r8D+I7hMHQnU1uDD2HFujK8gMtfXkA/RWU4237J7b1BUQ
LT/4z9G5+aaPwyILdms1yndpDNpVoz+YBH2bfKEmSSOqbwbs8TYGVfYOaZz1YE0nc5criKj4Gl0r
wX2FSTM+HN6OWwWt8iOlrLphAT2waFhXIsCyzqXwRdnouQjzxp85DHFxn/Z0SQMIl+dpm3l4e2eS
TqEhQA8TbEC1qNntZjHAmCSeEVroG2kgHZove0M4CB5YP0gisAQIq+RgZfFq679OElS1en4xOVSt
L0GdSUZvfaEm6y3fErHiAwyDhHO5YtVGfmM2oMzLJJIXrOuhVTIBcJnNNCDz14h6aNogNY2Eyhg1
vLrmP7z942YakCuhra4GlFtBhAKjWsWeOonVk4qwDDjPDc6cMlx28kMfJTaHWiPzr/IszQ5eAwDb
wCjWlb5KpmdSxtJmpviVKnhIe45PoqQvq399RRclKdBC7sGq3F5MvY2d1QhIEzEDgN61Et5BT7GL
IBzS4VH3etURB3HckK+9h7c3qVF80wb/2xXupV0VYXMQHpaNx2HdmYDHm2yhY6zKqI/h4OzFvb+c
FhKcIqfrQ9vLXYEnBy1zOy1N6nLax+83Nf/3oMBL0umJcr36md75FmEmCRpwmlTKEKYCKHVOEiDO
CogCcla3rHOun9Dso/VPTDWsmyIPQo+UB2fU7IY/uqqTa7Ag9evgT8oX5qJKUJQ7TSc7tfV7xnuX
EHE+pjngH1DAzoXdRn+FJtnz0/5+S6lIr7+Vv9KURp/0XtgZ+CxJ9HJz7JMZ7EUnuVRGVoyMSyjd
GphKkJrHO/0ANuJtAhr09gh+7KrCGEV3XIqU4GrVmfGb0uy5gRvgWJ1GWC12P7hqcb26SH1hfVTd
EcQ2bsnPQHtu6C53/lHitKX9REkI84SWBhhDvGEUnLxgJjeLKXmOevEV1WW31vOZpm+DjsqMsDqR
AXROV80Hn5MYPhUBSeGuKl1nN/2GGKpUu3himtppyJMOTnk77L4ukM54xH6lOBckcYu7oXsIYTQN
ZWWY86VpkO1XiWBdJ7+zRAtJgL2kB8lGjFzlB+yL8lSjCIUpDbd4ZEFvsuaYyA05077RWtJ27GF4
032tNZlAFVLBo1S4ARaZMBYE0OUA0U8xh6Nbks+rYo5frRlg9p4sOLvowXEQNx5kNkOGThZ30d9T
TQWEhbkFOshoa6tyccZAa8OT3OZ4xjHxGT8grMazf99DW86eZD0rHT1OdyK6AtzUUDz7/o/rkUNn
QVVXwsukVn4LkxeDBnsEfJt1rjsyHoV4oMapi+Nk/7oarhEHLzfEpDHbQWjhhm9fUgg8s4fVZwlk
0RqUnb5kJoDHlzl6sNLHv7HPLSDMRgF9XXt+d1iP+FgKjFj+1cLGIdFKZHcMpFYYTcTaavRdnGBS
3whebLTfH6LQ2Kt/pW+HivYSgoSelKJ7/3ilSzcpHU9v3qOQ2ir3y7H0pT3LtHdwIWmn1ZKtJK7b
snDUnxtWAVlLxRozwZ48EY6BcMzRITE6sf7a22XZy/GUxBDpsIbTb+lgRBnSfMpG5dJ2PpnB6w/7
QL0QxzOTk3YQOq7g6zmMlUkq5uBv/SjqCZt8NHDpCaGUyq5Bi6px1ZbXgZcdhJ6NdUdgh5/TuuVx
CXO7yXmovrojQF0PnYlQk1U68ttK0hBkL0ZqZjiVEYxh3xFY67sPkq2xMSzhQrGjDNilMKKgSfiL
aA2DL68KJmsD2cU/SfwsexyfGfRqF0SVSKj5GjY6xQRs6nU+s+sy4NpRbBUZ+CQV1wwhGJJDK+Kd
HF5XRPg0sOAC2f0WoQJcYt8u1cqhQRrjmcI/QbhZGzsqMZ9I1uvUw6WThpVIYEu437UScsz29iAT
fki+pOx6vFosnqESoNz/ozUmNPe0aMKuF6dGtnL7+QErrVo2Wz1Wcl1nVV14aNveSdtyBrCirzrg
KIXJZnLpxvu1H/EZ9lFm9eL0YswOQOhosB3uvazdgcGl+Y8/pXvbsv0vGI8fDEZRp7u4Jveifpjv
4keRde1VILPM96sOI9OAdkHltCwgsWKNG+DiP5wPxKYu2YzwKoHTMt0SOXZBrZHjWnM9BMVMt/zc
x2/B10ptReeu5qTVxpW6AyPuDikQPT+qcb6h44YXKTHqrQz9TVoG/NSBDFGC6a1kKZz+Df1mYyl6
+RjLF9TqU+MHcaHhER05l7L13vTQinsIPl+DbHFmKgFz0VoACVPJYVZWI2aNPfDl1vE09RtGCYaw
Lou4iC64ea9/MjRBSZo0OU+e54d/LqymFt8iLympTAqGJLG0pvZX9niLZ/0pNAsk9Q67TpuHhUMV
BZfOpy3OHOrFBeFdnKKGrVEkOuWhXBTDX0TLoj+vsj83xXnlf9nleu2d70MxM9i9bGgv8PGWyq0d
QgSakE1rExo65a6aEBQ9MOrq/RsQ1KqgQ2hR1VKVarABkoMGH4S4LjAVL2mYVzCv5odubOUEZThq
wPtSzvJlS3/SYwmrngvde0zjVno1FJ2zDGM1d0HdocwtEGVpsPgtMEW50J//oqq71pETj6htLHlB
IMZf6KCNNSc8nAcFbw+IKZ6A+blDfvbFVt4s2XwIg0EhCi4UqMCVzKMl6apWEN4YHqaC7wRWsdqc
HewulvTm/cpvGm+DYcJvRKI6a0pushjcD9jxaUUFNT0d3JeaTBL7InG4s6p5j4PYJXJMFHDRfJai
T2MJaASOzZqiuwkUVlYc9xdMDLnjd3Q+1YepwO6NGsDaQtkyAPvmXkp7TdXWk8XZYcakKPPFS+/2
glRpNNwDXFtVvngqIhaUZvZPDx/Y665ftf6h1fS3uazNDvkIw3AdR6GVbBt3TuBdpiUITb/8TpER
/ct8R9jbE+OabnZcfh3tv8mqZjK/rV67WAHMz8L9MVLI9E7t/9hpVgp8NpPL3VYIKIkuPiliZqDO
IrJ44NviBGNmDyjTmLAzk498JXNUGRPTQnuifkG/PxgukLcadv9SYBZxWR9hLfrvcammjs4eQUOV
RmeI5cNG8JH0q6KRODUgx+fULjgRsZWn8Cue4HGxyw0Y1OxZA4dABZGXzfe/y7R2ZMUUuksWwldN
QQvKYCbrqcOLYXTLYuAtQH0493GtlMRXmcZByGL/DZcpokReeDsD3n4U8dHypkuNydNufj0Lx/jT
BO6ymehup0PxUtfTdIiznoLWf7Ot5Pa23oAstbYhhN+gQ5S5XEsbcZ64/y2/3Ksy5MXpUvvX9pVH
4hWvzqXWJrpE910xC4f6XFtVFpOxKmRSIBZqN3LoQHIVNxEa+5EkjXzOe8A2fjNBpyOdguxCpGCF
8jSrBD8tM4W0BKvSzBF+pMP7zu/gZHO7M6AEuE69MHJC7VRzHTunQIqpayFvqV2AJuZyjO3GW3er
cHPYuoZN68Sn9dAk83+CPEWuCo8cIhmhbZmiIx+ci/vlGkpeUiLa7lH1f8rDkiic+0zUNcuYi3Uq
0r9bN+l8ceLkSjsdFtg5CVHS9IPay6nr+l6u6CCwHoE3JnMH6Ai9oGmf9/kaEXDt4c4GxF+3/Y8W
C8HqqXPnr8EdLIWVuYrPrUdZAZbkbfPqhWfZuWBY+R5obzZdWvfTtYs55JdCkSO/v50iEhdp3i5K
sOZFJk8gIt//8Hr1eebnUG+rguCL21oY73ZkSvlP4aXusITBJMN7YddcNZFOJHNojGEB8bfGvNQm
NEBd5hqLxHuOCGU/JYJCnFU5uUPQgOgbaa67VndtaD0Wu4dFbW459o1BuJi4smQhaVyaT+ZnLaou
3xM4WXE5QeLPLwvD0s4AzpcIvLbe20ceqgHjIdzdzaf6u5le6obK6qhdoDX2rCjOdVbBycCfY2Up
GrgNtNQT9Yt2DzBuq7jzBACIvNElDK2oHDKT26EXi4yHwIDFb5ej2BZdagIkPrcuwdWHuE0Ch9tr
iNlGX4rMIyyNm8K7MawLWUZO+ZV5g+YOYfQ0P6aDK2uXIWy+2mx5DO3hEaGWqrIBOCTGk7BkNAdd
2qNSLxtx5ihoAGVjmkAmnM/5kenrhNvNJZP8GFlkgaocS9KUgRuW5GSIvCJm2+veTWyFejRvYzaZ
1B/MB23jD+yaYT1mz3W8h4OtgqxRvwlQZ+gWudDkCJ6wDkVOU22meyHJjG5GMAaW6acIhfhC2WLU
0dRnPfofGcqCQJehDoQRK43gq7zABUCp11hPaS6gNlRYxdISClMMQ5xAiFMKhHArgzjQ2h58fYJF
wYAY6aY/X3adMDxN8Y7qM+/x9t8jAEVxZVCIehVIzTjUhrm3KNjcerZCWQFBSNERMPgjXEUdt4o6
uyUGynU+eXWxLxrNBHo7WxA6PyzDr+hafvMrtUYGvhFnJIqT7LQVCs+RBpUrNcO1Mshfa5e2oItQ
VPXKupHc9KMhUzK/MQkFHr6Xa6193qi9s+ON16bN9C+QNjQGFuSU4oCBlOy8yrowaCsfrxHI2r7D
cj63AyNfMCfMT2opPQb7kw95+rUDT3Oxc4TWw9Z74KUxYwH3JkjbiPQBA/o/s8W3T6U1GXTOmdXm
jZtgAFulOQ8Vh0Bn6JBSaaexM8fJyNEbzEHlgwtr6OQFZlDuLG8aokwEeJ+EYWkxTj6MKYzFB6NW
rmZo/dKN+wPzSprRCZfI/ThDhHHixmJWYN5uNdDJ8OuQvfubj55PPYdN8I803loKsAnbYUQtwYBl
2Ex81z2zNuQHHsa/uyZm3JlH934tdOA9fD5aJuyoHqLxtsqwg+24AScvzb3V8j/NlnEMQ0dW2tei
oAomZh5bRbkR9xNWlP0jhRIR0p0w7EcSB2cxk5D4iZbr9MyHtfTiCUtXKJ0mO9VawIM+v1ws3zME
kpO0qLHrk6kn1jCN7NItZCXJVUJpnK20+PRNsfYbnsoSnsQfehHJqVI1D1fzbEf3xzRjd6c1ArzJ
ZaUnvAW86SIxsg36BwR8iK41NWDWHK4V41wuO6cOXdjq/+rU29D8f9ovJ3cm6itG60Stzyc9o+m0
RK9zQj/EqLgYQWCDAn0oXndqlKEErMEqDx6Yh4D0Rn0WozSwTj8WBnEAg9wETAqntowX20SB3PSG
QDUdEbMrtobK+zWS3oos8ePEkVkKblvms/0zbrlzNqSL4OqrvW7Bc59xj8vKxCIgBmZodiSLqud8
n9iBrLng4XuRaTzsm8W/B26Ydo8DKz4/kObxLB4l7rmE0oFI617IK8xkyy7zIMR+02SExr0A782K
2gagl7giAAEuUn4JqZ0unfQHUV/W2J+aKHtU+/ksHxvUBwOx9vkMxLvrl5VYztt3VUqQCaTBtZMe
0Cl6KLpqPdAG9IHwrZsPzzrx8+vewqDqvTvBHPmKK/1c9YkirDHQvfE/98hrHl6yRaGHpH2rF7Pq
oFJrqeOrqRLSL1lVP9LJq+HUu/P/L7S7oh4vtz7wT/lGs4Q4o6mij5gNJYnU/lT5YUAqyMEHHIuT
FLqg51MRgRVQW8b68OKFujvUy3Jy38JL0jpqWBXTAA2cEf/8PVqBjeeQcPriyJvzPmbbuwPOS4o+
fbPXlFu6sgNiHSLXP/gSSZlSIoneUnfyA+tpmeJkP95lcPydru09S1uZsAUX3UtvsEq8RnWW9bfP
6jVJIuWFEyIDUEHggCPY2j2Sxd34qeXWmmATyDvmHEzEQbjcXRodNnTrJi06Qoh96yaehR1XsGx5
KnCzEH+qyzUdCbGfmplOTtGga6VxYzIDc2ws2IH/NacWQxRaAczzOMYl0pXpWjsfBj/ctmi9oDBj
7XInB9x/di2zuD14qAaz9D2Rm37qzodtwT+/rCNGHwlMqriLhS7gJ2nRfkVVciUMaqzner/sHZOK
5dKHhWCW0qjFnHBkmKcTQdfApAaDOC9jPW0ci89OutQWqy5ZcI5I1+81t7tR9440kjUAbuqVL5bV
jCXk1/CNdSUxuyN+cP9Nc12bzqAP0NvOJleF3S42YzgtCkO4y+69cw12W2tAaNLdvBGJzQTwNmLS
A3XOgqz3maonNEXHdLS6ori+1rICTpkfQ9c7quZmodxt0kwiMGvDdSoGV1UHKnUJxdnRgUiu00pP
rP771g16nieB5uI7ZdvlXYiMn5H+gyLUfAM6f4Yf4ekXay9wdtuQ9jSH8kVZIK26DwMNOo9v74wB
osc7FZ3b9KuT8hzEW8IYJoxnmpIuHPmQD6wenXm3TWL+ahLquJZ/7ppNcVrQralffVOozZYQ2NZI
afMcHMvappFTEOrb672ktNKi7UQxA4TbriVXIqs31JmdnDUm7ZjOP/xSdZ98mnrkarQa867RIuZT
nBd06DvP9pIu5fcknwLjImGM9ADawlLIypEhymNolBt930arXvGozYRkWoEjguhuPNb6XfGAP7NE
u3i4+C2afdvHtNkiylj62N39wBtt+IVAvC7tlx+XSYIJ86qqanSDOvuZyCp4w2DFJ2G+0CpebMib
GHSYY1Qd26hZG5M/8W+wgL9c5HmX+nVhes6d1gOLOK+84ajO/yiRWkAGsKUr+4WKM2a4WRqBoALN
Cwbm9xHj8YSnyxX57t1jP9/YwRUumXcWGnL+17s9RH57mHwyreyKBJu5jh+9RKxavu5P2BEx3VJa
wDYwaxxRRhKICDpG3US2heUR+ZXyKRdEV6peP9vbyS0TvEhB86qQ9VIWVnNwzx3gbUJ+M6CxDTnj
0EVQccICK9o84tSHW+GkAZhTK9N6Ahwi3KtZdblv3HJ2i0FNkzGWhW0n34tH5OLbk9qh6Vox/kdp
48qZJscBT2POjmD/wZeeXns2Dby9lMmeOgmT1X5UgFAD8dze3SLM48iHKLpJfN49099S1YNE9YzM
Z0xOKVhwUxGUF4tfkzyDvKsUfyLGS0qmvuQuQVdvikbtHuoE45KQYNQt7WE+qRV5i0VKV3EmNa9e
ytvTrDjrKIkMyUoLJxQmrI76vO7G9mLHLE90cCLLgoV6r3xHuHufHA2uvmZWKGsnxTKoIx1A6h1O
8yghtmhi+axJWtPlmuZWMOoUcgEjBZSBsuY2LiRKCHnH6lqeB0FmKq4SZ2ePlfOL5eVzzXJsxZNy
N/k0FboY6mRk5fcM3nuPx1pdSlUbnXzDzhw6ytkTe0rI+b+cQgOcb5qeivSyNgJXGAtixCk3QbVE
Pc6K2JhuL0GY8096Aa7Xh1jH4IFL90lFS3M5fKqlC2Y4E/+ZAsBhZp6FD7ZM+1v/0WRT1PGuye7g
4fgghoO1j5Jib3yoLb5JEqXnpnEc14e0sVdTcuMKkVAqe7xjQcOmfhNx5o8fNf7l06jQmyTptK3U
edalPqAuXsL+c0YDyyf5WB4Py7zLtt8LiG8xvw9IfAtTIlNuysKRClnBQN+g4e9Upr/z609ZSeYg
6f3hprJPpElhnSJnnqAcQMJnm1XCSdit+xaHm01trRRHYHSMQ+eQWDK0gB/RxwzJ6pk4Vmgh87Qa
J9p7WkVEa2aQNXgg5wy6X6/g0yKxKmLK2wX6ulkq8ObvJ50cedIfkL4K+vZgLOXIDg0zaK0NYBC3
71lQuvOOP+hinXKJDchgEOLFiSi9mEICE3J4f5GQhDVMkE+QcbIbhnIJrvSZQSTBMVeHEzW7MygD
o8b/bMvnXRPGMcNqZ6+eak61wIOGYD7rNZCHpQtNoUOAc+EaWtYDnGez/ozq7ibwh3+8H2f4htpR
9AfHcbshPTPCh0weseWDC7HoaLS4rcoPARluA5zFXe1bruuHS2QYbe++30LTmsE13EG+vAlRD0SF
JS+glv26CP1+n5qAMl73zMcAjfciMtVn4wgClrW8x8/FVcyGG7uF2XdD+GVJGrrj/i6rFhe4DGvq
6ohi6iRSXZQ2JecmidLY9fgm6oXKYs23pPSgL3cv8vWbg5QjqPUp+oNB3Jk/D16fHAtujEyLklrX
uAJpm24HhEJKozT6U/k6HsG6VjlY5rb3iyzSZBbxqJuDFHeXBKJAVw45l1HlE2bfx3FJGyABTipZ
knR4rRfnQZn6FkszyavslfqgvXhrLlP6s9XcWYoqT9U69VUtzW+WaRgjk1xoQDiCArZjj9rWy8xV
IpIbKnnO85aYzf632LO7blCQ7s5auf21PBQIzVsosZH4EkIYZZXgOlVG/rsw1cxwR1hxs+4jZk3m
eSya8hFD98/TvD55CoJncEDdVKKkCcBHcP6iKCV2CvXwWinEBzaYL0nOzSB5QAWyZ0OvlI1xPSnv
lBNpqKZOt1TODiiqjMX2QqgFX9YkxQc7Mw/Txr0tDowOzx5l7ljk6q+xaT+mrzrVlTSSVkMg3ZR2
2eSFHo9G6hLM4ZY/aGFJhc/iOH2WE9BVW5LawYsH17klXDCG+fAiM5LLzDbFzThFDsYhKT+0txf0
ObirEFIld6aiMoF7J2Oh5Cd0S+8kPGno/n+xtUgWBYSR1Yh3rnFJi6+N0NO3DplnxlHzX3cysw2B
atjxvGzmLS7cIuaTajI8Kf+ZY5lLSqmc4SAmPJaSa6XCspWeVkt6qD2cJq5G4uUrRYPPi04tpT78
qCtGD3ztTA7LkzKZiSg64eLJ5DaqWeK99rAau9J+GFXgvP6bECjMx+Lg1sgakGPQYk+bvddmW1wM
HhYGJUv1KlkPuh0T+P9cNTpQl0ioN3/tfByr/4ndZQKqiwxVUrpSjxjIwTUidCQcc7myltgPa4/W
VwvDkD1HM1DIShqCQ04msKnHUWo4FesaFEtc82vxLFC0a+FlnaBt6BSRvngUMulUU08AQaDh1O+T
iejpy2TXsNgFpK8/qNIEJc/0mSo3kzN06SDF3ODWyuRBFEpC26OrWMmVlXjJUHBTgOxJPG7usyPU
Au27nokld9QT7kHC20NZFSZQf+fvdljIdZfYAdUjWKYS4Yf8YOVCLMBCTz9wovXilRFBN0wAUjxb
mdGJwpj3jCn6gBuLHsuD0H7+xHlugyivmZPOLtSMxJOwyUJ+auoMa4u8EZdruZlVBMzgUwjEOqfL
vlAoRNEG/i+pBmVRaqlmWPi7BOU0cxRUGw/LiUIvqeCu3/rSdDeUN5QPe1wOkafh9pQgsHNt/4/w
b2030wlyRb8dRcHDn+c8XmKj699+lIaxRDn1hPk1HWZkxay/LqxILQS1E39f00wa3OTTV1AGL8TI
QNfS5gWBCG1y4Co3w+vP4B0fNEfizTplIUVmU45c1FbY2ji4h1J/lpCE2PQ8YmVCaS1lPdf0T9QU
isBV1QVt+Y31ffBlDX1TZoSl+BLejFJdSFzFarTw82o+husems5KJKrpMcjw2uC4meh602ub6L/F
wWNqtjXezIvBKwqlAZD22jLwXyVzcugk53XGsP/g1KOezMDPmgij4ffEKZl3S6/93UgXZRqd/v0P
hSAdJEQoyt3arWZfItpMwQVRvpWz7+q4iagZZaxeL97V1jTE2O4lXUDJCDs+lu4XiqWDVpk1EyIP
ymklanHL16EBxQkxcLfIcCBnqEoxCJyht3eDKutqW433QwRTZB7/dXZlHvysnGyp7K/WqntpYInv
rCMGYyj9FlJ/oev6cQAyqJvpTv994/zJEJQpv9NkVZjyu7qGIOlZJzVa7B2xZPrfLNKtxjcI8Ury
gHmoyV4i6gPfkfZppG4boeayS8kUxXqUF3Zi3pevmtSa4L5ucQPp4dFx/uVFmtSABt4gL/2+Jq1I
+VVBerIoC+7xdieJWKMF8VU6G7bbymLKY9gnRfm8TWdQNlPwfY8zWVQF4wHNdm1RHmOBI5fD6p1d
uy3zIyhQ2yFsnifnMH4f40Fnfi2yRIUbuvRqHuIkesQztYELodx83QQe0JBombtPTYMWju2t+2M9
kxmnODyO9VFs60zzPYL6lKXw8FifvBnFpxr4dhnfeThZsvp/KLvA9FMfh9ZCG7DOG7xZ0Ks3CZJV
D2tVVBv+GMxlS6DmPzyVguivDeS+OzlrWLusDXL2vq/vhAE/sc6mHW4yCRIVGSAaPSGkDYj2s6GY
8tSPajxpUdD6wV9FfSr7FUOc6jxpkAr6TKFWUhD9dcGQp6+TjCLAast7kmfkft1pomD+8A/qZy2o
0mf65EPXsaN0faYeR7Y4U/rXQ/tFcwwhxUXOa3fZw5NAniCCEeQATb4MYIrOlGkf9L2nEqKsMuht
NUhufZC/r/eIqhbGcyX5PI+jdgE8AyQ1aPwMDz/DFXuRwHkAOVh8gtOB6PIsyQnrBiXYqYpxCDwu
HEM9+82RJzLfycpb0GvcBXavNtSKyG/7WoHedi+LOXb+QHLWsRZGWc9L0vOtU8fwYvfyduE0JbV/
OsTQ321ZU5c7wj/ePdCgJIakAmLJHnh7pfZkAcDABVgllrj60UcZBM1OUrItLd2F1HzaQ1+oqkkH
fqWum4+rmSiL1thqso58LI2deIZfTfiYI+GjXheC0DWx6WQXEvBPsLZQCtaDGDatThf6ePET+LW5
Dz9QxKjSbk0J40HP37A93+2h0IKYZUMIci0KlxkhIAvOSVeOG7V+FCvNE2+N/ggq9sAAldTxYvyg
upqL9t7xmiDrZpGI+QbUWtlmXbfNKV2LbxHZCDBGOAMbwizTtS0K5AOBtsqIW+4tIFcTevHgblD6
Km7VERp980d/UYnf5lp4pHg8KXE8JjJLMLN/cqlpPpNclIhwiALFleQiNy3Vek1b0NtRvNigStxq
+Tn2z/w8PdYvxeHRfvok4BlhYCG7VwC1olUuIQRRsQ7PKygUueoFG+38d2IGfveuOtfNOe8i7/uD
2HDS5kJJDZZuhWvevJf8nu6QkTvOJLU7hL/DlFZY8CfxIF67lkM962BlkcMC0OyPPo0mxqaT+46s
cHr8orRTOwdNO4QqZerQu1udZbdZH7eYYtg+Cj6yfBkcykJdB16rPqCQAKu1eubYIshk6/aCnj18
9jutoQlymvXMmN2aGl924Px0ajNIWZsXMo2RVBMkMEgcd/tl+HyWvkLm8nXHOm7M7P5aOIPq+Jdd
VDb3sAYCABcOuyp4zimKzZRnO74KMf8ntMrIYhBIREVdjYaNQWf9PTtmm62johNbNbxL6heNl77C
p4zedzZ+o7rmvGUMhr4OBA1ULVqclZGGY+MIxhp94G3ook4RIw3LmMnfAGdPaAjmDW6fpuOGXV8w
AKs/6Tam0hzzq92Uho2Xx4G0Okt+4+gsGBXXTHe53WDk6I7IxssK0EahDVbstrtzWdZju1q6+tVO
vLF745lgi+Vx3KvohUtoimgboNinWVdyx8PdtW5vG/EMxMFhg3vASniCShf1QnzudqcIK6/YW6Ce
DUlDHbtNecsL6zeo5sPq2Hgxs6HgVQCN71B2JNqY9250qp/47yL/Y7mFV6/kbSHSposBvXOx/9AR
t/Fnbjl6wo/aNvCWDRrarB1Uadcm3FTkyJadHS1aw48tXtGIUg7zAR6pfpvDFt5SVCIOjL4IKVue
SXkkFcccF8v1iRpjO6+joTUD4G60HABQY/mM/8z5tF/7dzR8DjD3SRWdfT1msjv1/XGK/+jvqeqy
xRqtotQIYXX6mAWZM2mvlh9Fbloq+d1oWUDx4qDBUelbSTI00fL6n9+8d6kw7r4FB0qzGhaBAADE
N0+EMsb2cpsG9rIkVrYcDuotKkPOePA1j8yyx3/6CdIOfbu8KBKaVdbu5nOq/O/iLay/z7cqK9Ko
2JtMvr3Ig7FrEiQeDFRHjigABGCBVw+AB0uhpBMN3rAu8O1XKFY0FhAW/FjsCMwR3cRMd0i912rE
XMux9ZKPzQ1RIKLjoGzjoVkFpKbdZsENOcc0Zt8tPguXzS3qjH8wdcrtffADeYqYwSSmp1zGQek1
7bLPEJh3JVZo9oLttqYGY+c2wEU4NGJT68vpdBptSlsb9WbbC9fCHrq0wWQ4cxt8pVxShrEnyD54
ZHCZjQn4CxbsA7t7H1K4W5VuG51elgr9VXr1kRZPHzBZ3pAIyx9OKi1J0wdA1YoA4NNf1B2Hfo79
i2Pw82wq9g48CqHh1SMaYBwpYwrLn7Q6phinD9hBl4pUZsUTY1ZS+3YZiY4k0kHMO25WEWLjsAwr
LwJhxgZbTsMRXJfEf0I5drk/nPdEvZMq6dmZkyH3dO/3I3ZuSpG/C9rXoqpjf6yLrD8w9svQXK46
K+RN1ICEw5bsJRGy23COo09SS5yUy1DEjll308OTPLTxxC1ZYupMag0QqCQiZAPxu2cy2r5+1k2A
00gZqbE+iS0Aqm4aK3rG9yMDPurbRy8J3r+UutmrXoX7QF5dJpqzWwDxFqF2DqMk8j4un3T3y894
SttJz7rYv6XMGk7Tf1e1KeSO6+OW9FxVS/nLQ1pBVZjGt1ty7daq0TrfbbVyNyVjUYYx5beOFPWt
6RyaA4Fem9AIKg+RAwUucwGgNeQCVkaarPV0d6dcf2uIxR1vDGLSj1vCVJlZ5hAutmKLr15QzNrH
CTr/hYFprazypNHqPo1FowcDaM9/aYjR/AAOkwX8XU8NgCsq608EA5JOUX8l4it3FcJNNV48+i4e
XxPaLBD0PbbvNNH9bd0aKISK0fs18ps6OgjUTVXAhLbBFJM6HOetGD2qwSEi9JtEV9Q5DVbNvkJB
bI/CWE4svdtdAXnvU5jwL6PCK0RR7p68vw0kNdRK8z3ATF8u+sial/3/f/wjhtuUt5f1R0alSjri
nh56YZ33OcL1COj2Cbk6c2FVN35eLEXjgsybZb5dJ4r+0k50dmABKb22Hr0bpfFmy9Kyg0a6w7sJ
Hc5Olr4jP4ejCmGMqS4Ka88ZRKkimoszB/FZUmVtMQ0drDbHAscffCk2xEpWuJZwIaRokFgMrnID
Mrzjn/WZL9vBgiUKsBVoOlHfhVyQ5sa76im7MxBCmAi2clmiYJA69nR+aWlq63E9twUw1+AThlIF
Z4sN9+cOAycSzQSpVvK6Pq5jqLHxrHcNaCPaUXuZOMG2yumNk33zR7Uj0zULhYnlCsC2pRxea3V1
zOUaa/t39Hx448uYnydAMGC+gOkF5wWZWHqRXRk+9DS49YfP/WFJ/mzj1v81xYoC5IEOvi4LPkAB
DgBqHVTpDSrJ5UmECdtwYtTMfY6D4Nr8U3OZHylYfFsVT0ovFEeTnCCRrjArCaZr+tbF9y5lS2Q5
0BSg/3IgVnRyZmgFO8vypObOnVz2cCzGH0tGBnsif1LmD8vhCg8BXRm5gBDb3syLGhELmG2r/XjE
HUO6B4AReBo2FEqteE4P1yodC6+I+jjZbjcKAOx3koh/hONu6ImVjtQG48wvYQBolfWBeHB2PG8w
Fs32S+K+BEI1DZE3j9Ij2zl6K7Y08FTz7/kIC3CkYOVptSliuHTXZjqsqPNPW5tp6eRlaM2zy11X
EghdNaSSIZ6qcEMrHiwIAWe5RSLECybdJraxNDa7CYMEhSpePza/nQDLuUGdWdXFx5GTgPpoCWFn
Ovj28Nv6jYY6MWOD42ozjeY0Nu1nqQQ6xq88rsp/kpVNgBOOcCW9R9LnHKbJEsqX79G6rYwL4zH1
ZRQAnJCF5ZTVEoUcsMLH/Le2s/Z+WWXpjUk6kphPtD+r0zudAhqSUH63YWIiKCPFlU62W8aV+WV0
e3Op21cyXyIpWWhqZOMoJnJOsqoNgtezpZNFVYzjGIoYkvIaEXM5s6JsXbUSJcsLlMLMWpqs8Gf1
vNGPifsRkWnoGCKCdJIlxbY6ytN3O3YbcMnDwFe3SsINBDbBTlod2hpbu0WLv2uz5FeDzfRueE4I
mrQpzP5OkCZLh8o0DSmhR8RSmo3d17ZAlqD60wtl+N24hykcBmqjG03DHUc+/RqeUJ45BujoOyaJ
rcUK1klWbA8sqdp3mobvaqjJJl1Rg2/CMhZoXwOhC8h1SCyCiOo1aerEk1DdgRRcKmDAJOuaGzW7
ZwkXacV48oYFi4JyN9ZolMo6WW2AmXYC0x/mnVcSFXrtxgmmZiL2S2dQsZhzdPZKAk7I7WoFswW6
K93drS0H0n37ON9MntC557oGf4n8vyrYzbmpLzPL9sKVn11tSkyljPcCXokwElv0lwPvoPdZh29d
0RszPCD6BG+otgsoNWJugURCBfdXGR8vh+Z1B/Z80lDZQ1j6MmSU6l5LD5i6DCRr3bVoGcQSwtKV
eSRybbHZ/5W72voZ0+q/3gWVMMHS1S5xisL/Kczt6nzzbC6pCE/KL6Dn5kGSwQ77nJ0oA/2JKOEI
xrZzkmhVXYMPh5rxXNUVR/myczotZenZM3nnkGnat4kmkNQi2/FS8QAQkd9ehBJii+ceeDATD8Bx
8Dz/yPJkIrgsR2elmB6aS2h5rpa6wImtCU1zU8OdqgqiKQzccn4kBK9/ZMlkUlpKvk3f2jx8O1Wf
IibQybc/4/IqcZ/IAitwFJgKkvBo1CE+Q99dbUH2p6SqL51aAMPLgrMdVGY3XrvOz4Jfy3OY26QK
PhV3/2Sq/8Xv2tGC+ltYNz8XFDgoTdeuODW7kg1jOAhIOW0azifiU6V/yG8kPMB7tFzipnyW+ChU
inzBaPKvOZzdkMagCRfaHGYxDMbVwlkckH/WWWFRH84+fChIzTzfkmEBcLNN4qPYaInPDgiA6JJI
BWuP5Ua+4Q/5gM+ov83y9A2KCSrhIBff6hQVQaMfDVnDhh5L+l8D/mV4tZyhxSfUsayp+G0RontX
VEWI4EOoWbjXHHPwqXYcyjN02gcNacC4xnFQKaEWciCYXDGjWC2wKJhlz571XeSjDIfG2gRj23so
X3pZtpxVEtYnHEmIhqrWftEI0/yg5TRSB8n2tJPbEGhkhdycwH1doK/DgROICMugeOOXezdHBWSM
MsTOwobD50H32G0gW/t0hGsxBGeYlCn+G66ADfBWwTNwGQaPOjI+XP3qexPIgEGNiclVEFRmf6sp
RdBNAgPJOs8Ni3LF0bpAmsJbRBUQqT3qzbdkw770YUe5TdX8FpQdkjjB5QlyT0Mgzl7ZVjyz6pE8
E9ExS83YjprMmG1eOHkxflBOjL/C3MI6BaASLsgrZhOh3phOgjR9rvdVbqKQsYfO/1KYjz6b4zng
KRzlI8a/5MoQ9uheO4knZwzTYeDboQjII5c/ayW5Tsz1KOCdUu4IsU3PoG+2dtLT1SJWsKlX9Vms
1tLkpPSO7U/RpgXW3piU88Dw4U6+fNEhIlMyQSVtD2qqAbha2E+8sCxdMhPuojB8YjCsmBGMZIJU
R10HZWe9kYEORXAbMrIlgCC2h0N3LL3OlM8nKO4GjcTOysmWHAmZmgb77k+difoM8iXJrwW0HkJw
OGo9A/S0ffTXlu2GESy4W14tULpwWBpLczGzHyy3YMdli6y3fN3Au0jvF/Ol1O598Vhi80jeVYzc
U22VJoX3q25Q2fXPjXu5djVCsbVjhWqm+PL60h+maJldFZ3tnZon9ffjsgAg0jEwwSqt3c3FSk9l
IVKHV6NVllRlu4mUn/RLBKXzR6/Vd8xzhyWMSGC8dS6mVer71fK0n5jpv3bedOZgpop1p0WcWG2H
zfH19qVDk9nDVAZ1oJyIHGzBaX6qUnzGDHOoV1EtR7J4udRstCsI39kYRYGvaOOspruqUgDYsI5d
rO1Yu4hsK7TGhYnyqUr8LerQ5VqvZNKs14BTlfh/64tYdF5UQ1M2MYnj0GiTypWHFbTtJIsE3MeW
t73OzP+LjjzvbjnLXDgvbVstrwmchBeLXEweijrLe7+llUpETIilfeEq9wI7Ck6wlJYdB+IlBeDB
c90qVzUIE1PpEh31dCAlJyRjXa8W/2aRFAC8FtFuq+F6cCzPOURVQuhUoh6bNtGSfZS9HX4j8l0n
D6Hfb5gD8PfnGWS2+bau1uHag8/zMLEitm9Ke8wS13Gf34y/mr3ls90Xu7+eY4BWsQp5S085vjZc
W/kcjk1XLQ6AoZHRUPK6j9yYl2m1xir4Vl/nJ6H+3VaSdSnuhTxT202uCjQV56lsp+gbWa6kXah+
ixxLPGml8G1e1aJ2NVM3xdoKbiotd2xzg3o253zj2+ZLJAe2GDQJ752+PpM21qP++ZWp0YX4Nv7d
7oQo8kUzfgMh+FO54fzXF20WFocyG47J7CjRlTI/LYslHPx+M2OaCCAcoQSBT2ZsPVFHSB/q+8KA
rhJ+OgoEOT6YRm2L/NqbMSBNDGapgh/AelODnC7yskV1vmPwLG2dvWkYny8cs6l7MsWXF7u+xWME
ZDEJlafVgMM0YA4GDEMg/WdDu3Gn26t3vfT9OXuB3OuDOoYw5dcXYUY+4+dj0tWwKPxtNZwoeHIl
jp5mevAoWf1YnEvsGSZodguvHqIk8e1cJOHVf0CrDdniEQbt3E8Eni0nUqeD1FAFCO7fP/D37vKo
zUKpo9vwUfdyAsBFw0EelClsr2kGJy2PJ6bJ9UIgTeSCtM3W8p+nEZ9X9ewL/sbYotMG0yVk2zfo
UbJ/b4ZEbxYToC0UWHrSV2o5iXdKvUIWmzg3I5Q4GLSs42CckzspAIRCP5VBKLoNTvt0ZY0TgphE
GiKluRU0JQRjVh3Dvb1iWURGfkspqQPCkIuZrPLg59CratN8DVDfB3ocPulgcdZ9faKms+EP8yjL
egAr1eryC3CHFK494gLd0rZ66/pI8cpcPvkfwPYKvm9Jf+zxMPQjrHtbxg8/w/Nz4kr7Cvw+gJa1
rC/9ns9i/mwwc+w9V70FL+0o2dCCyk05Sw139SGNwk8ERNDCuMLz3YZTL0I3eDcE/3kvhMYR2FRj
YFIgerG9cgt+rmeNWpjVxpXHSmDmPC2pTbqsTGMMsl2vvdJJFhgqRABfA0+xzekdtvbIXMcPPpWd
7Q12Hk2lwoa7ga0pqxkurwlxGEanQGUodlFc8pznPafuGKSED9ip4i+fLJbtr75+NItC+m2AX4h0
7JI4exVOTqRyKEHGaLDGFLetoyS//5gzWvgTOQsqMHSe9+Tsy8YP6HMHr0Opw5KFt9PCHGssiPoi
pTgC+rwszU6clZxAw3RTzDOlLT3CHH5qR9LyTSYU6gBeVrhWnvLetyz3K3NrTCNmESw32gm+8tx2
ZhSPQvg2rhYIao7KeRDOhBqAIwvAv3xAtuVUNixQQM5DwJscP2w/m78yygfoVDSdA959ee41LBuu
mowx4UQui8cHLOHSBO83BjreqPBxBlEYhLwwLRV/Xd2BrPWn3lXvLKX4w7rau/KJAJ8+GIXjdV7h
mbtw5vZUFOi+LgqZePjr2EEnZwHP2QfbiKiA6q3NxrVEgejx4VAt5C2u7vg/5xNchtttgzBDart9
UZfTpAPCyEu6h0877SUdqWJFTVWTf0pmTKZ1Um7FYymkQjY/k7lCA3WMFLL5t5eRRWAaAH+aWfYr
eNspQdG51jR8lw7UuEAd6RWpn1bXgsUbdTPxacxT7h+6VqJhKJGsj6UYT6IaEYK0cHP6vdcgGIFc
i7aHWI5ysgO5bOr9SgA6fVYgirIFP+gj4AF6xwLbthZj2u2TUDl06xG/cuFWG6xRaReEIWAH+uQ9
li/FPDpdsZ7zBSpN/o22+ollsacbb/FLr2/TZdQJxhIuJz5PLGYzbyen8VoKUOkTUkOiwmxOkZkb
L1oCVnVpERckKLZo7FokU3ZVhdhdhYjSd9RsHF4nIbxR7rWldDND7FQHjlkx11Tq4qIXM4yFUQyy
d/4wcjmSL4WDMHEtJMZ77FZWW/BMbFOlYOM7PW1rPu4gyvvmnR/ElLxf/MThl5VUnWruy79bdQK0
1IoZAIPBd2zsTruaWna1/BDSu5miVNVsXJZ5E+SRUf58ywWaqBWesDqmhclL5aSa5sjK48HZftYg
CP1SfiObSyXtZOfhOSwylW678FZheXt4ILaFMQyS+RLtNBXrVCcXL6u0aNFKM8U0XJY+bfwJWLw9
b7e0KJ9RQhdL39GdK0jVT2+D8oPaXnH7+90LrQXe2NMgLyMfTZYWtOH5/aZ90Ql1/P7KEkwWphWO
cbjy3htGfkaEhbpeGfz+ESd72coevPsuNreJHN4aZ0BtRr2BrdCZts2PLUF6ph4mh2xjJAmXCVDF
38kQxG7KgQcukDnEd8a72C4YXBXG/iYtoB3NvgrXas8HWr4PS8xvPzaq1sKCqstMqGB6h2bnZauK
2JZmmXuH12QcEq01ElUW7JtxKAM++WcEuXhqVsyeIbntVCcMExBzdIWJW/j5uz7v2WeGIyLbLBpz
rGlVtaz9JwhyW9GFl+eGQQT5i46ilRiH5HwJTV8tMcZbmNWucSSw+izVpGPA3F4zmmh9GgyWN6YC
cZhIrLjeBGmRFtMeY6IcHkFeRw+xWOwe6/DpTUn11bAw3HHqkYMJMQsii3rKxlk/qZprUlRLm+hE
ndUmINY3IA0mRHPupSv5+meHncdQhkyQIjydmpybjXtAzNkzYVjrXe3Q0C42K+qj+DQWxpOczR5N
39biqqbibyDEK2A3Es2JC7l9mFVoLLy+0BZ7yR/X3ttvyXfeKYy3FYYeaZ9ZyIaCwWIlUFooTObS
UYYj/ra+GTki+c+oDz/t13rwy8HYlwJrGrG9ztHVGz4cY0CQTigV0nKGxT4fCypFF7F+JCnMPwSo
oQkV2Qbe7SdzMHyLRs4JVHaM2+l4+CYTCCg17arPzpQMcsQn93TH04bDvHUaj0pDUWYmW8/aHlCJ
2+FLTrGBK6ZtbK63G1NCU2CNhsVqnQtlAKOGIhETtzJureD5fxUzPw87XxQzFqcSarCZmU9CPCgx
Hx/AbYSsBJmfQsYxCu/pByCxzXPAQx+kBdmz4g/v3owFfWGh9KtQgACVj0opmid6/5Ih52GMDmqi
al9jVgTh3I9E1noyV5cE1PTVkwYRisOGxOm8EpJFMxixDHYrdJI+5HchHb1E9uNsQduwjR0UgfvN
Okg2XzRl8lbL3WX48lF+MF4uIirkPF2VSXff2Qx16gSZIftemM6nsL7mbV5K1w2ce57RrPaiG07D
cA/lYMbMN/L0j+1Sa9DE+78wR1FEsCe2Fq9AA2RFKIZxUU5Ql7KD+fHTqUhtQFg5uyQ8Bx38qclM
iisijGa28v0skw/jmlNbabYzp+GF7RetNJUe3RzSfoQlc1QyUDy4XSm7+v8VuDIl96T+C0vXkjc1
66FWFBg0LFv5rm6Y5I48IVlkLdMt17hBpXxWf810YuTSDxMJjqIaOBMhSUp4YmEmtmT7q0zZl+PL
UKR/5gHxYGana1tPzttR07ZBhM+kuG/FPFZuJHedoQho3jY03yfksMTXnp9B+8IF718V/4q0KKDE
i+OQO5kO07lYTbAL0LukYMW8G63HAycwd4FLOUwOin8EgH7BpiS3d+T7QgD26GlSY6LwyKIwmDIt
ugbhIjpYHs6Um+FFKuH0YPJWKj4cztTwglfT+DYYBNBpT9JwmnlvmdEJ0VAbfNDwUrs6/3lXPlI6
oQhnzfafKRL0J40qd4O746nZERU9Fz+W6YqZ/7uge0XLca8u7NtfzxREaA4aY8bvo/GigK9/a7o/
3Ui8Y/B8D3hx5rAkeuDJhGkYSJjL3+AkOe588LTmaqNH+AbCuQ8wJ34ox+u2p4ZCmcls7/m+w99i
eT1dbR3Ac72gW9BsFh3AoPdQDzbAxXvv4nRse1I4sAv3na55mUXDD2Py8vHmoQfIsl9lti6y8TDX
j0CzzpbASWuIUd5rt/QzxYKmyxL8jLqPIZfjKt/y3ZnoNwuKmh+YeyD2g1ngXUZDktGw0aMBdDNd
djfhsNJmr4eLrxKqjiliAkIesVvImqxBDv4A22Qh9Hk9zifTtTeTFo9NiQ1inv8gox3QG+QtsXVQ
4aMbPDPZvf7McsUJX+eI8PJ7eACXeEJRCg0sBvW1rL+/pHzX159aQnnDokk0R/5dWYBtvodRM5kf
hMeAUUagxocgLXvT3vNQVq3dywRW4PnODYwG0OU5XtqE275mVRHSE9IJoL9phX1MESfCax1U0WeI
hkdWVYq5HHVUnBLS5JCMN5YG6QWDMwqsB0jZhaGtOcQ1sapm4BkYRNeyrnj/EOK89p6ltJgDTK3N
HRXXHhTox/nu/J+iZwQ5WoFz7wyCW4bHQXbR9TX/GRNEnsPZIW+TfUCqGkpYXEjF0mzq6GssUe+C
fv9s6qh1U8TImq9xTLSS6eg/LZuDUAWwDlT2g4Ejdu+GW9iZHTACbBBYQ7mXLk3laoCMvyXIZu84
wPhUaM2NatZAgFx7pXV+UuVjXrd/FPfu7tBDcsEa5wTx6/kNZ/Yhnsg+5oa8sVjAa7VzYkgpvHZG
6SL6K9Ycwq88Z+6ihC98NKB4Nc+x70R3ouP3ABLM89ubfgwwSYlFDOV1N9DlL1J2K4kNDmt4lVy1
KmaHF7/OA5gjt0Hen9L5i9NOEyvahKn7MvEpASkUi/EHNtqXsL/5UKQ4sW+gK/F/y6Y5dxwOLlJX
ZBPvRzEBMsdPYtGRFpulh0vc3NWUWOICkBXAKeQcH5paEkboeOW1Y2QyoRfsICBDTs55iiUZVRP4
AzER3Ffg7PRYlSZbd89YfzWB/5aoY6/Bxzmy8FV57TX8e0rlO4477EZyfrWQBfV6LyH7Nxy/kf0r
XzbIWLgwjpHe8UlyzHgo3sZTmUB4QtvxPHgL+0j+CoaGjTZjZQAqYgyoZ1XWDMNjPBKAQnitjbK0
XJCtrRidJ8oldMRTidCI/gMi31GDGnaDx52FYPgliWmG1oEWBCRtbqXRm8I+M8E37v7FYpOG0kSv
YLAeIu8XMCJJtzLQBVucNf9rEnbmjRflZeKU9cvl216kneD+48iu+2ZOVqks7Z/lr61FV6KJjldJ
PjrMl5bHSPdS/pEBgWf5iGHfM55V0ECPbPhyx6yilm2NnxbXIPF8jknXUgVuHQfs9nyRgXc6SMeH
umL+li530EdGoK9Z5zT+oQyWVW9t1UA6BqMyteBBTe+nSUtjHXPo1kOOrFw4BgE0u6+jjiIsCJPZ
9Lmr9eBqkH6SsJrSrNgK5r3VfzYtOJanDfc6UB//YNTj464nTbp7u5GU6Xve2Q6K6q0ZBV/uW3X+
3oGcunsE2iTbxRcmNrUgn6hN9NdGppT6XIANw9ApaIAiNL75NkaFR5sxjipjXkOdW0VnmmMMDL3q
qvUXRKs0C7RgU9ALX7/H0DDUf1RRT0On0Oc/puw16SbwpHnuzt+sLDJ54XUXJ2ANZGF9GQjg7aCR
ib+VqTO29tLUIFcY9MQ7xOT98NOaPKYQM8Q6EBYDF10gN0LQLbzsEH1Lmufew8HJEuphw9WNroqa
euVxMIOIg/brjcK0o8Y/XIeYbsRxqj9RtVs8kqy0yAIzm9ChBx/FLH6MtALHtRBqI5sAtI7CAHMm
TPj0v8NFdD8CjlT524FA5Z32oCAFVcIq8BInaiNr03o9TIT9WWeTPfA2o2/UOZE/UvW77cNYq1PH
qfrotA4MAb7XZYWqNjXGJ9MGdTHPrMAiQaU4lHnZ+NzpsYpqVPikt5l6Eit10sqsjVwEC67oNZL/
c/IdJkmD4hZDyrJynJ0wrMIfZqIJkvhBCuq8AGF4pzVfJqWqVNX1lLfRa+ftRS1VDQFWki1ibPzT
IzQD7uPdQBWqzFIRb9YjzMJ5EIMLNjHiYljZ2n0OY6B/EqFmiiOPnutzV6Sq/QRLISqlnFTL4Xuy
kJEmKkSeQoZlvA3ee3Zsc0hn5oj1bWFFSg7ItVHcK88LW1cUec/VmFTYlJjA6PMBagVUfPkjusXT
/C5LhsMzN6epyu1g8Kf4EcrYiJlnbk3Ybx8oROQ5oIWp0dXyxoNtAqE2nYNdZtPnI3epw0se4ITj
flc9CGSq5DemFJTeRR+ZQsYZFtJgx/BJCSRFkYn+c+hT7enpVvR1XXk2koDlWX8oWWi1YyPqzz1V
saz2Pt1k97KLqKNnDVre87o6u2lF5VULChrKjx1XfyaL7y7hfwHV+QRTlHKcEMV1cLiHtcJZs/Kc
zGAZP2iRI9Hp1bmzitWbSzavYHRCVvzxskoUZo4a4z37i7LMGxsu/Zp1k2HYhCAnE2HRdtENw3CC
vttk1vPy/hAm+0Yq1+hsfa7Pirh2r6yz0in0HOWLYGuTCC1Hd7Vlgfq6CInrpn7fnmGO/YJmKSAD
yQxoPKZl4OKw3x2QVnZv/UYsKk+8BW+PK0wIX0pzojpQLSwVNQyoD51amifeWreTQEYHiScpBjh8
+Eoakwu7lt+FK9hVzlYsba4FuXj5HYF2IdGO870jOYdY0dlzS2DLwxvXnmyz4GwgYGLSilTB0MUi
QC8pAGpllFkb/ksjKXoDko33JS3Ij5oTaVP1gnSl0lD9JlDtEcImteN10utxunDQ6j7P1UUFmcwW
hQCIwtLozhiLzb09zuXyAOXpYsgO6JwDvj7lje4D4tPRGEQDAz8l82b22la1rRUV4ZYqtLtQo187
rUWr/yHA/P5cDK+fkemBpqL+Y5O3IloE02cbjHKGmBHgsDmSG3Uv/BcblreOukPnsToXkoXP36+V
NjHJMOGwAufjsO8HMQc7fCCotrRjJZR663ZbIw8KZ8C0+yo6A37Z59TOya6PIultbICtQcqL0qaw
sdtf2i+6cIdueu4CH6nLU9NnalzZKTLhDWOSy2faCGHCnJrL2N5KfCCBM/H80qDcOjnH/shjZ8ww
BFgpXD5SWR3gyc9x8b/mbzRY9QLupjLLDsv8PsJqi2/759GnZWAKZQTZqUGWe68IUeME+uBTjQ5s
8j2dKHX/h4BT9NBqvP3vzoe2v7TCEFR+UKFOGI/KqmQKcFGbHVrs0mJW2s+STlCBdjNs9xHHbBM1
+DtEhdtqBrn+ouYfKdnDIZeo1C4HYZ08RkgRz8cAmH+QQI8gRHIn5vdvejZUcMcdly221OF4YlrF
Pa6bvS3z/9zAZYJO4iOFojMhtpCGS9lfg5lTalKf/Qq9NpDQuuOXUtQHmKV33XFGnV5LRen9y5gx
kEYXZbHP0RhG7VzqKkRAnsmeeIpk40aibNuoVoPWFkZvj+Wo/1WeYlRVvz/WIm2jJDJ0HgTJu954
aX/5jL4h4a0t5hJOFm31TX/ai6yB0fDQYu8Q1+HnIA1bL4Wq7U7QU7Kl6Z8DB0A1IxYyOIG3+A5x
VSvln9BlLj2SavXeHF3OgvAOwehITPmzP9Uy9YHkCP0aXiSObeR9gUP0Boq3CAWIhHTjoNKRQInG
o+Q/W7cyKmXcpCUj7PNioa+vplvcW8tbn3ilNRfcUpakKdWNmx+vKL1FrzsVtTN5wLkWNDm8efUY
5JV5NeOmOwMcwVrAy5dJ0oFcXlBAWtvHJj0cGcIVRfY6iHWnFiPyPgeqf6aQzwHR/P5uGJ4/l0Rq
0kLSmAYJx0R/d8QNprP58NkfX12lA7J6l+U21kBIxDURQVvoUzSqDPcuoVDlTX+ztoZE0W6q1hn5
NJDUWsLAdWwfoM0Spw/rxVz+a212TjMmSCwdC715zpmN0z8FUHspBXrdB4zHzVA4Kxvcb81lEOqy
mA81n6LZ3Fp2G3PwvwN5v9GwnMK227V7UoYQ4k05wAgKc96e8flxe7VleooUMo28iL1bASD6ldm+
Hbub4TbjFg65qADOXIyzbPD4ZyH3GgyDBbEwCyyj4mu9oUxFsvG3oXQF5wiIPN8rmGZZqow4J8rx
MPEWLBNMLdCuSvmjVDOSVrMBCPOJk7kpkd5lNnHav9/Zsz60sEeGWq2p6grpcC9fcB223d8t3JTX
DKckugiTT9tfwJkzlUmVA5Q7fjZMK6nMzxVHBT5upQ2Xzc95/MqtnMohmtknBh3HE1dhCDac4ztl
WaTReJ5rf2Mt4JfxC1d0ZZbkhknfAvTNVXWtLmRzx3xqC81UQG8ZBKHWCH9W78F+T2bvtIFSXlP8
6CkeRkfiJLBwn1a5ocaLCJJtYK0rdVh7Ke5V57fBHqegJr4eXWU9tBF5OvBebjIX0WoEKbDvvvHG
6iRheVWX93C5jNlmIcqfmlfXe2Moepxt3sMZtVSm6PZJq7D1BwZ72P1EBAEGSk81t6i+JO+ati2/
/HWnuTourrU6v/E4JQZnUHckigte18mDDK6ffQeXyiXgpNT0TKDIDxEOWfwBu1B6eVa3atuKNKSW
MeJT70rPoGlFybTK1DQ8bZqJK7UIS9ZhavhK3NmxIGxakG/tXKeqMMDPEE79qfZUYp9zyLixcttq
p7XAVXYej95LoO0AZgpK3EUTmiG2GEcktb4an31MdxGjVOu8uvLMoeaYP72Hd1QuVjGIv3VHU/MI
VNQ2lQTWQ9ugsCiDJNZ7HYG97vX5RH0uBg9GLC2iEt9IreSnDzTRtS+7Ph+gvRZ5ekL8KfQqqaZX
LoFqkdQyf+6MFotmNIiZyOAiQaNnE82NvaUOblfLvh3WGuHnWsaRPjY757yqtkGDEtcXKvlJJPCu
3/Jx6xrMvzC8PbZGLXQEXt2OwTZ1XdNxGtpFpqc1h2JQAvz1JgWkRxEXlv5pMMBcvgT6yHXrISUD
ITFeK3XIlUYfVLOHXe6a02v8ASNilK/QE0H2FBmvWAn8SQk4N3zO9299d++bZ1j27l4M2DAgHw9K
ANgMWLGw56GZhefOte+zKJQpjX+xIxJguXa9ucplyAT7k+ekB8rwW2BwZU4GAiuY5MjSoisA7gCH
0Y5vRf8+raqxHRFJXj0k8dqhSXFZPa1etQiZ1JQa95nLTBXbwRVLe8lYy/L2BkVmLfZF9iNiWtsQ
FYwMTH2wc3G6vOvXEo9JRfp+f12iGzNANrBe3xE1GZr/r9Z1pToqWoCgIDg5pAXa/irzY2YD/XTu
pCgyQedokOecNoN46l2WRUyY3DWnj8Tjf7ncGP550x/WQwiH1vAXtNw2QtJywXIVgzP3zm8S6Mxv
lnckDaWmlN7chhibeXKDKJwrBj3/vex73easU7Zyi5dgRkeBFU7fSEJTl9BB8lOI079xcGYHHIsH
3FwRp8JWKd6hQAuC5aiWwNRtdblyIwePb8yxvdf01xNw8C3FXdB67BA80LhUNmjbL5gUPGkkdZn7
QxB6Pxwz4DTDxpkVLFwTUHuaZVl9VWpRGAod0deWZ3OVnGH1VYZKHq7h5cm6MbQqFJnM1TNK1pPh
rBLU48vWbj2nGzVqbEb0wsyKYQwauphBwIr7St+MMP5o00lFOBmOo3h+yp1hir6f/hPJz+Fu740a
+a4+jG3pWKUm9I2izzvrZsqf5L/XuuFf1W9xcX3XvTEyth4gaqHd1/NdLOrcu3jXMHO+2sgyewA0
uq5Bso6oTzov1r9TKb8VNNBfnS6UQ3Gn6wA3UKAhwEaQFsJ9tfVaVyCmIGRSZ1Vfd7j7TDX/gSaO
dHuMfpMi8PZh6gWGgzxq8I2OsIWpIZSBocBXJfRpAjw+USYNJ6LKiuGb3YO0SVq3kDSdsqcA1II3
YLiLQP0PnDY7TrJSTO4a6pXGXIR5sPpz++EML6QIa4zFEYlF0ESba/iqYVu4UOETSPbRQRHEVBcm
jxyQ6/nJfjxbnoTUASI144EVpvnyqt4kyvg8ErIbMqKtwLh9EMQTlDsr4WXkqFeAHNxqNGhKUSjK
H1LSdUJ6NqSRM0TgLtX9nhlUNfDhXPSomze8nvjiYfm7bwEQ5XCBZEvY/SBsB8hNQ1s2882ZL1w7
A6/dgqdgzWXdJVjTfy3Hur/coAq/DTkHjUbsbzPZxsmDcbh9BKTvUUElrCLZ9h0E+MEP+en6IXWA
AadrnKMcV4EXZQyOSNiTpF+rvxpnkbOd2gZy3pifbnzF0ZP2cVeo7u/dEw0c8gSwVoniWbBYc60y
N1TAiO9hdmlGXaIGKpmrX5V8sSEW+yMRP7mS90BGN4IY61l8wc3UrD8XTC9Chbn3DCB6kgQvvfEo
Khc+6awNI/v6VXUQFlJ55/ZIIrLS1BlrOhpSRtGVB0LFRDr3vJNg/HdjJsiXrBWDH7FwrD7wV2FY
ZkgabpghyCCHkRtANkHsh2HyW0tAofgg4Sq1h6efQzCz8OMYopf642ne6xMJNzGnLYC5R5h5cp1T
5D+AVH/iMncYnD9jfN7LTh7uE+Cqe3feoY+XdxLnkb8HNKd3wqfy7lghKVn5ofZOHlxJumvhNenW
VBAY/u7nBYfEI9OKNE2Vyn0K4kUkRSj2FRibpGLEWAiE6SS2DEjWTj6tL5SlOO0Oer++fYG7dNF5
oI4VXsBC3jyFI7KTaPEdFgxdc+XiHOERENE/hEqhQavEreV5M6GpCm2bDBgoaqX4BpOKTActe2XO
hiBZbdItHX3ezeMkoSCT3FXDX5lldpXKovIiAi993o0OIeVgyZcL+m7+n1Xor07wxCL6Awv27mfw
Qoeqcukb/0fG3EwTZ47FPdrOES/RuofNM8pqaNR/xfn4E7SJwkUp9Wci6kCYdtS3jYjwVDgSjjOb
qrRZ/4zJpJSNj8gw/htGmA0qAeQ1TAAERlt6e6GTLJmUbRw1qywRafcAP92ul/uEWXlJ6ZKNwHp+
zjK3vYdZpzQCr6KfrUZ5W6IPXe+StUxtIlf9akwjUwSV3M7j4vyYxC/0xgeS8sbq53srdQMezgsN
0HLRhGOeTyqq9pbFax40+a1SXJBVuPL/yzNeIz8lvde9HLRJu/TP2yjGA/Vh7Hxacapv+kAmWyQE
ZFeOXAnzp4YVWE4qxVBq2xc9t5c3TILgedYQmAit2wkTG2OtpAn3VEt5FrkSFGl3mceCm+NmrtmG
vvsZu9xBvLBrQrfQ9qIaZGF6DjwCwK50guwdpq1H6qYnYdvL200pZ8nxYkDN5j/+HbJXd+2Lub30
BRbQRhQ6a84XCtYuq3rQZU66ELJ9dYCzFnwCiyZXY7aA7XNW+CYt6Us3t3rAOkX/Khg2suYPczPR
DR0oIiBaf8/OTCEtnGGLxFGmvYh1pGHYyenDas0SN9HWLhrMy1hVNA7rqD2JgpCH2Bzqh2xnrJF5
XBLB1CzQv83XIohC92Zo4xqBgIS9wJXUrAjh+YQBm22mF4rdwqzI/dD00K+EwIkglvOX19rs1odb
iE4wYUVOJzLdpsYZ/+e53uqNzkMG1NZ/cc8zFqOWODQMPa3TDp81tme3gE9lxrsyAxPhqV6LDcuO
BgayS2zpH8PJ7YSoLy66IPor3mr8tWZiHvhZyJNjIWwvgZNSvz+QYAZp7VJq9EQtdcJKNuecrR23
zMz+obekc85UJfwrWFb5DdXkxZ/r7vy6FE0FqJVqqomkWcbR2DumRBRaq9vkyTU7fXi4e/PsQNc9
r9QfA8y8T+1k46BX+kdrDnyFBajES3zN/6S0Qy1oRD9AGojMDmhqbXx+vBpPiF+RhAjo0i6V45wn
rBeIAZzgnFtJVmoedxszPIvT3vyYOfJvj+gcZnnO4XhBz8+sk8N7XBFGeuJMu1jCv0NSr25t8YWL
uEiBpbQ0P/jTsgy23BeJZOYVXt50uYQBXZPSjtvgZTe7DZ2FLu+CTMtXB3EOQJivb+zLqpnhHnIs
mXJofODMvL+Nf1zLb9f7M3y6L7rpOhVqxtddM3s/ZUJuhn9VkYSdw7/MC/KFBm+K2K0/iiuBkbjC
payyaYru7+vqCaGw7d+bLcKY6FQmFjGt6AZZMqXrsYXDvqewvNTawH4Nf9x51imxIRq7a5kZ0w/b
EF2WTDDK5O/nQqcOTVAZf5F8oGs8Xemdm4U5h3sIw0xRaha8m5ErLiTmTeK1Jy/mQTON98ReNGMs
AJ26LXkiFo/PSmCTc44hHnJQTrtsabFMaix7Z4bMdsmKqxc67D/AbJ4Ro6n7JaPjhS8Mr48U7KXA
x/JySLzEPUt98wvMTFmWB11VBvgRrV6/9U9RYJEatrxLdNaXWJlMIA6XNiUFiHnzHgEk73XkOvMJ
+BSJr3vjXmEZ4wkwbHiLbRRqHFDJ8hwVylNIUB0CtUg67PH99LCSISHfkwN6hCiaDdshAvznwKwu
sPf1WcHUTW7+O8MdxunnSLmtYLdqoVPKWhRrAYlptAMPG+SN8Zd6XIc+LoniCzoRJfknNV3Yqnya
RAmTh00rDvA5PEBHW2RTwhaabkzC7XNXOFBcLRSMyQNWYo1V3lqgYwiHi/6ebdMIJfEDb9UZ7u15
HjB/s+hxIOKeDOWK1eZIjrs0DxKs715HQR5dvQCqwTfo4zQDHtNrak+/1KZwNh/fh4qlfj0wmHtV
L54xEdeX68auFUAWtu3OH+027yNfmX1GfA2PlkRVEU7mtNIUpjsFASQdJ6Xfg2/cyR4k2J7eqZZY
lFY0tNBsptHBIu71H4V8+tYFh9M6zwGhV4ugdADsjhXuf6xD3uexTnO9BEV2E3avjw7tl4K2tRUH
LwzSzbZD8gyCIPgNtSwQsK8/Yu+CmweNty6c0sgjeE2/1M3PPzuHtVmgxdBIE0OIM323+mPJXX72
Grzh+Z6WnsjUDoKAu22iy4gJsW51ABZv6ge2Lc7G33tsGCfhM0I35D4xYma9ris29WWMaESqZcyw
sBo8hSpAdGmUI3gMIIXQpSUWqSLSuvUSLK/SkBa2it8BX2KgMXchSuEXeaDBgTdlUKQ/tZmrMgYd
wLy7c8tc3lbmo3C68F9RHXt3+KngthoZKFdgy3fT4ewJeZWmLE52t8bmTvGbjmj4N6Tp32x8Wf7l
EcM0eefFvnVra9bquxIjkddpz+3oCsI93Ai78qSMSX0oog3U8KU/4hP8sPeRMGHd5HZJIhoMDyla
BtX4Uol6X2U44RYINCc+yo9Hm/3hgg36WePlJ1D0uXoW0SOYQFW1S6KPg3lKNvZKb8a/4sP5Yq/e
HLrDKLkUg/Q7QTc6bUA8HKyukbWW7PHFzJOtfbn5h/QDLvdaf78rzF0btORw05k8cgBO/q3NzWfF
bxPP7mvZV79waaIQjWYRHPn0Nrd6VPn1QoyrKWhwP0ZDd/8R1qfRL3dfgoJx2u2lHkTe6Ck2XOID
MfnTa5R9nD91iT6SDt/62y8ZBqNI0ApI334NbOI1LRAA0ujRiEtdGhMtrYC3z41Wxn6T6WasQv1G
+F2745NK71NMmX5JYwdt915Rha3JzQdsWoE2Nz9MMk73y4wNKht2I3WpUniOiRewWGHRxfgCJTqz
Wx0aucEO6gCWRKg5FocMeDUWmuZgK+XngcFO9VaOmY7seRFNNy0HDfIO9wT4vox1oDtoqIOMHmHE
H51J6MQzxPN5iGIZiTAHDm4vNA9RWdIAc6zvFomt6MgoqINFga8TytOLbBcxG7oDH6Nw2VBMdFfp
m4ngZEKqxd6DM2Ki1UKi74Rguk87M7PrFtTwEnPPCM5y8mUKvDVYhUdOLt5IObqVI9Qjyj+8LZhs
m/peC5ricvJtc1lbMFbbZxZwKCm/3dRrXU+WTZVU10ohYWouLfO9+9c3K4KMyBX5Ui38r6lpupMH
nepxMXehPLsAm54m8ip37J4ZI+7Cq31KvygeBAyHiqREKsCQm5xaXemPYlc4BYhabODz7NV0GOgh
ow3VKG3WCjROEOwXeqcwNb8CMmJqQGpjApOs3LkG+7TZlPkNOmxRYh1vuOOjSaun+jeztD1JC69a
tHq3GgUns2CjcEiq2hoHMDGgnYGfDpb3mpxvF8ew0r4TWn2vvbFwe+6vM/s59yt1yYBXGP+vUqrk
zAAajJqMHxo0eqh8LT45dHBOY9KfpyMCf/YsG19ECbVG0vCRIigGYb+dKtirsW0Js1fbPVAUWOxB
MIgq5Ly2P31xcCvl0e0wM/KKt0DAku5ubKt0bQB1pdk+083e5CTb/rXc1eejck5zt2mAY306VzuA
EEa1MN2iHIe2810OWe1iXEsoykE+zV2HedGccwQ1sfsYXltcJ8Bak3Vu+FSGJHeOSb8BEwBphuGV
2Ei7YnIehpPV4t3gsiYoTxI5eQfhwf13K1tGD/4H4LfP0Q/h9TncYOfH5+RqCxhnERLplOgEEAft
PxR7X5WpZVO7Sd2p4ASHMlqz/RRquSk1fbh1Gxv3ngU5v3w9chp5iqARi/vlgDh9gIayPzebk81x
7m3oKi3RijARw37DdnQTCAUpmQQaOpQLC/Xj36+5WNce4sRMt9p5kIfNVgHjuhxz6lQFNkAqb7pX
cnItyzExE7ekH8Lix36NHttkHP2SrXjvJEnbDXHo1IdVld16CxR1dsvdg8EpU2r2kTuwI+UuIlkI
qvQuDDVsliZefCYaMWYtoSkD7Ajt3AGfru4WiRUQ71oDGa5cBmP6NqF0AXTZNufSbS/XJMu0W6TN
pSe7Y/whVEIqIbEcwRFnCf8b6tt58UweaatdsjjGalBp+V0edtxim15aj1FK/oSuoZqS8/i8Wz6q
1J6YiC2/N7Aw8B8PdfyVXgr7qhQQoTwU8RrXhpkIZ2W21Su5ReByc/YhJoAaNIRJU/0iBZtIqMNo
rxqFRV4E1OWkykc0Mie/wvKQYhJZT7vzguUZ9jDqrOXSxDAeNAMk7WRpeaL1jEAEJemFXPVquXVe
U8DNOozkJfGU5osroUeEIHlBgnADhUheS5sHbjYxb2ZnUSUqR1DOzepAxdLvstTloG63TF7y7aQs
/zCadV6m/6PZ8Ak7wo5iGtMqaSZG0GjVlqksBtZDDn8JhHqknEOwHol8hKtIDQ0+BEg65ALekbQH
MYJwuIfUwCK6O7QeGBvMhuT5sZewoatgPzuvYwHhXpLijBAt4/9OyWhj/zViHLuPs2q7bHNpvmVI
ExRItC01gzo+NumivbNXuFpYGwEbrhYVyYTctS5zBmRKXBCDDSWL83yWkqeRj8M0L+RZg7GnOMug
XMo4MULWbHw9PTL4nNYclMule2OEW8y52j+MMnMuHJuHO5YEOWjeAmsdhmwTyGw3SAjPZ+jofGaD
tkiinjSgKKugYzhtDiajyVkxeOz3i3uGq7Y2PkhV3267rysX0hbiaCE52goyC3HQ8fGbwbXEACEm
9LgZ8a5KEdreNQ1pNHY1spIFxrKwpmO07/MbVtlHKr+Ra6AG76TSHFobw2qH+BxR1f4v6npzjbFc
ufZCsuMxfUYx0WZ8ujHJDcqy5ugAuJD5V5HlD61/xThoB9HluO0D6/w9DLPkcZyHXPABR/FdDqpH
VQm1ZChVALzgw+0ZpwxTthw1VX9RAZE9dDsloLl3m4S6wkKs0C5+GNK8ouVpA9J8b1Ddy6YKQJcg
jgQkJSO6lKIWffV2QnxYi5yDLrGIN+KA20kwZHVs+gePUknmOF2nRAKs/Yli9ie79U8n+MwnuIIO
orMp3rS439xuedYYACCf6/tq0wPHa2VUjwors/2mzmlRCjUuVDGuMdpmoUqsSMo5nm+MRsufBc7E
n2zw8URJI9N+n/yA1fNnOHz+QKBsN1vrknPRKNDV5Fa3Lk3vEteILcYexMVUaeEiRtPs6pfTWvii
G2F+kZ/Ywpy3mly9JYmzW4KjUh7zzxuN4MQ0xdpgDky2PoiudZsI9OaWlzzPplHRTj1yjzVDLHVP
r7yJzoeLdnLkZCRAdVKk6Gv3/YuVUHBdBu05Q0CtIeAvlKYa3v90eYEjWdoFVsTSEjn5bFszP41P
JGNzkB2U+tRBp9MnlXjMEloh5nrykNFjJnVdv/DzVnTOkYQg4NqKgMQ1a+8ZGigVk1L3FFGisrO/
9a+we7kCuoCENVtdH8SIoNfNBGuO9/oF8QB6hM8pMQo/YnVnJQZw4+p9hHnVwmXBT9TrCdpO1pdM
8mErNYWyJNg00VDPBLN5EBdzxIPk5Y/n4tm4isHqOhDZs93gYwejetQNccszp0IWdTDVLIt5OJSg
QO6pknO8Bw7ORQFwMr15SgzZDStysNCXZxU0lsh7dskWFiHr0O+qFD2XNW3MugWABdE0IrW+vFsB
/QBEsynxzAG/3ULoPx6oUoMrLPgsu5e3UeAAUxMpoRHPRGO6GGO+xSOArFcaXIekNuZEEePuqbOb
76HLQBdXDSZfQEjWQRvujdp3B+UohrmXxJGF9FJeW4v6AiZcTJV+xU5WmS4A2p/rTkutvhbtkUl1
9fdZ5Sj/5LFS0dlVwWbe4g0VKyHXpdUvZ9Xvv7ANFXKyjGyGeneD10duLLD5KwZc/pUeebk8rjkU
vnXUpLx3ItbbJrLtEdU1z/CIUa8bTrhI9CX9aqEDq4fL23e7NHDsWt2+3e8F3lhpINeHZYQ+AZXp
zUDl/ahOw9ORWz7WTrua/lw2G/tQFvf0raq7Q7zUGy2B5E4mMInHITgxdb2/nEiFsrtYtsE9tI5G
gI/tY6KeAo4mG5nivXofwbIXusfRBNBMCUbCwAdI6yls0A0FevA/+PjiQYPcut8I2+X2Toh/qJ1a
FMaDlGhKKF+4Ic+sfRTGx9yNa5IIEyqC1Jc1nn81cDniv5OaaeHsrzJmPrxroxhZDqYstBkhgwRk
kMebrV3ZF1gN4T0bPTxDyv9UOY1uOOB6hi4egwgSIEwXgEWaCLxY+7CZKe+EszGpq1VbhFAK+RNM
0OgqN/XDe7Yk62Gv0ftGt0a9Q2NHJXHkNrCoN3RGEVAoFMEhzzc5ftVEACR8FS5PrXbq1++91J5L
WBNSwLk2xd8EFBmT6X8DrqYLOWY+LjSKDjpsrfcvLyFlurP6BlSMydzyCEdzxFf5W9wRZmcGE6SR
AfTb6SDnnKKoXC/fpcp37hgHUqoTM3K6TQF6n5IAMpYeSk8586FvvaFtPgZ+5i4C7iMFLb4shX8e
2piFwW9qeTYngx9O9XQrGSEIgOSM49rP4khniIQsO649flrmDysIF349VUVhQ6wSketQTQdQwqq1
MDEGnSG0BcK18w7d18zAe+uGGYrUGFzmaaAbE1dRNqnt/Xo8LmikTz8fpCr33aZbW1lQiem3Kvk1
EzbarJUFs2tq8UsH7r4zVDa17DslxLdzMp78bBWdSEvMLxvtnipnMoDLqE2RT2trx2RcbevQhmgw
8gV8Vq691ZtubQ+91O7w82j86A7vA7i3kwNO8CnUpHi9AKc164F8tYwJ7MAKwBpQVi5BIOweGtpO
AOfVvdjhb+cA77zieAk1eBm40X6EmK/NtuyuNcp2JpwbZukz9ZofVheCkkQNMQM8w/YGaIZydz5w
HDNX55DdaNQ3iEh5eU+kXmczlUq5vdlXqBOsFlb8d7twEAUtFTh06mJFMDLzfU8YknblqvG+2c2p
gQnFZI01Amc70l4nAuP7CI8jkImj8+gHNgVcUCH7m4eohuJCggXa3gsRXd9yJDlZAMefQueySG+l
K/Yegvi/rbnDrnQV3NH7V0HxplO6XJMJX/7vhS6CDwX6+PSWGKDtOMzx5RDcBzUZfOUQjTQy/dIo
lkTeJBgpP9ouSv8ciy6iugqeoIP3usfNZ2lyExtJDJ2z5oXobsIui+TZh/aIW482raM4wKmYt7uk
W7basARaxWX2S1cyy3jmYG0GtupwjnmBKjOhux8pgSBko5v4u4WqsXKS1xf+86AaVKnPSsXpgHIl
PkiaeIQfMlnVQ2oVzs/5EMK2+DQrfaghKCUhPygfzQFrnKWBVlgXO9xB2OzDJ3Q/omEJSPpdRckh
9V9iAT8JG6NS3L09wgN/Ih88ZhfKz5yEtv9vxSUjkYVc331sXQ7yorGRR3Zt7xbuKDJdl9bWuydM
AN6RTFF06XQcDmP3vlJE1YaGQuWM6IV5M3d2hlQVChoLw5lYKbcUIoBtFN+e7yOI7f+mCvaj9njn
GTV4UDrLBYtkRusK8WNbL0Yi4Oywagvf7FDdm/2gRdV5rp+ezfQi9j72w74YzziYVT5+ElA1vcwd
JKC1y6H34gjzyhd3G2Ix/mC2vFDoTDqTsDNrEWal668e++AiPBk+k3qfq552q3vxfbN5ZRfoGouh
JBXSowUbUoKxOmQgQJ/8IsrB4hWFW08zCBUIizX9v3cZbso7bfvFuhP/KNBbk/mILDdeCNkxbrPZ
bz39MizXqfCB/r4F6GL5pqYxv48o4fIqiWsPxpPLXH1jt1dt26UyK66e6V5Ew/gGL1QwRiJw6xU4
ACuknClLa2BJXwAiiIhuizOkRik2heBuGvks7yx6DlJbNeaxUROA5o5z+QqPKn904/rDUZewrs1H
yGjmK7b4naI8S9dwg2kLrMAaDZdouxVIFs4g1Ye5c+7MVYtfD8FNww6kZTd98wNWRy8eBlOa4m3O
jzDZxEmL5P3XK2Yf28IaXH97GFvJz2pc3QBcaWxPHvdZ7T8DvVYUZSq5Jc/qMkDSiWsfyTeAsBDI
1ajFS9AeRCXgmBfQRoVoDOKtGF7h0u0OFm1VotauadNN0JBbbfgHFBQ29H5xb/+mSMm+PtdAe34M
pdzV7xJk0YzoDNW097aNV2k3UiLL9HFoNtS2IWWZvJmIThy0zE59mqwE/EVAvZAW0nZkiNWoCyyC
suo/GvT1mJxN1a8KZOti5+ZGY6oo0PHLtOfHpRs5zreK6bxyrxH3PRKb6vN6T0zH+dzm85VwHY4/
CJKZvYzbbN3juiN5w/j3LLbtLeaDlpAqUDjeHT5dL85vmcIDEwQPSL4sW9rkW+zqk0vdV1GfonZS
XeXSlbHnHMP4f7Rtre7z1H6eZUqX4K49MIr0iFMYiIhSFObGUOxP1HsFnux7BhQxsFhsGJXxwd4K
vuxAK8bE9FYJYY4SOGx07WqQFhvKNTunFHAxPf2S/LkybvahKq9khl1Q9gnKB02M/ZQysYofx/mE
iTDCDyWptjE+nWqLOusBGabh09l1QUn1voboPwKlaG2LrOX/SDZiq0f/lI51F32t+tcme7dSXWNR
Bl2b9fwwPECxbvgT/vxDswnSaqITJP3ul83GyBgO+FW1H4I+9c/jIrZ66CDa2GgdoiDJcx2/I4d8
ayUgIRCeiieuPXuCt9HJRaSwEg7dFgdq/Tqp9yLWIsrl+jSVdYKRbidhCQk3yTOz9g8AqIwoY/Ex
7GGVxnMrEn8ZFYp3/6tjAkVqmEoDv8ui2AF9dwp7K4QBiqndysDhOkW/AG7bdQViXGGiUfgkUbcP
LndgidhzHUICuNkIOLXpSKfdp4vbGHWJqrdQu2ykMLLUYmpKhScqzIsyrRoS9ryZHxIgSAaVAF1E
9OaV7hKyFm14Dkqsc//HBYeAwDkohOqL+OWPB/1rC4KHLb5aurAv4GcjfTjeuR1GzEVa2G/N1vKl
E3J88E4hlzz8Jqi6penlKDsyf3flBLdVAT0m593PrcYihE2H6qt9RXkp0iSejykZuN5fDUYqvSEO
HngIS0yB+GPqMQuIcufwTVFLulMtD8nYPmusVAdRmhfLD7/c4yYJwOFTOt9bOjXebRN6xBP3leK3
AV4JM5NGB6E6NRfe+YISGQhM/cz7qZ1s8S33TWMKQS1jwV1hTkHuPhOS9Ca/rnCSWuknxgaNyLjP
HAGddHOISkXWhkRY5cZaJFcSDj49LPqe4s7sIW0wDRZ+rreQbaQstDWZBuzhZPmv20FxiylJsY0V
nwTZjUHc97j0bDUiEzVHr8iPJSUaMRaC++AzHxaCFb5nLBFivy1yCDyOCv87UQWj6rT9Qop2v9u8
OqD53B/LJpQsLD/lZawFZu7oAcC18a0G39EiFRvs3Q1mVrfd/D2o6yZFsu3W0VvkMfsSjkzmfeaI
a7+D66y4DNYRDGFs11qTxE+q6z51IwXqGjMKMJtrYXVsjitXJ0KK1r+5sOnFjPHXQ3VKbXmEZlh4
HDF68atbD6P0sdCdlPI4QXSjEwwZoh4HdlNa1XAr/6FUQtC3E3zffjnxfJ+5ePtE2k6S68I3rleR
2JgGhBsvVsFnHABWB0XlYNHhauxGqLYOop7cSMH7uvDixJtgiizymNV7YWn+FPJG2bH41W2Z4wbc
tgjB/zr0EBrVFJaukyKKaXFALxTeqWENgwuktyH7iXdczNcHKiZ7A/rKEBDxW6fQTRrfsDNvpl5l
MufIDYSi7OUZABdqQ/EFFnh6AnvSA/JXU6ut4txW85pYO+UV/CJrj2YcXKFkmRWd58q6xNfnvW1y
7T7IdmL129Bfkn5X703HZSElymvAguSI7Ki1fe9NzPLnO2WGr7skIlh0U5ebZhLuU0bJiB52Kef9
X6Ef01M9gIpgsiyHGCkjuW6fL6e98tHUuRgkFVPoYAuNB4CrkyF7fSabVR969ySVypP3DpkuWEyW
gGnnkpg8Pc86z8MAb0OpozAcv+hnJf/11/ZvT/rJwvzo60RttdUkRBlxQ/44jekfSsbDH88mXIgA
2hGyqcJ1Mz90KHhVwDTMu+5YSwJUE0eBjCLJiVca3wB+sSmUZhjH0MveUtYoq9aTY+DbYx1f9U/K
D4pCDESY+piodpbY6y2ig+GD0PeeWzisOwpwSgR3beRNxN7ZHTMpoNKSWrQLrUwBiC4ns/iTSaiZ
U2sShepDQgph1Ql8l9JE1+TMsI5zgzr+ybn6wsEVzQf4ThqI4KHlvDz1TbCbsniR/I7CC/tT3quA
z+267oiFR2R/Ngg7gxFbrIRL2q/S4I1L40NpQkunp02sVfhB1SP3WuvNL1hxmHqkDrv5apuSVP/O
6KxXNUp6ECkFLhoHYT5btf/SVsa0Ejm3x6/Lsu3ULtRPmWQ7jw1SzrhN4vSDc4Nt7MN62XHCkpzY
ZA3oOMeYs6rJ/+B4vyijQwU01s9kKRxypmVPdbyJ3fni6tQC1N3ET2nRjmzKj+U6uJU7rgq9un7u
8sW5a1Nqjpuuheu35qS6gz280lBsapcS084DuCSUsxPvNri/UoQq0h8uxD6H130HjYhLtCeB5sTU
SBHhqzcFnHCluibu4Y0/CFcWetnaAo1hdZe7BkE+XXr0ymorJIUsMeRsZdhCy4/f/jZyTAPof/j2
uzDcx+wX9sRCqr2BWU70j/OzynCB2nh3aME0lXqrg01PqPrKqI3d0MHypPykuZ8XgAfMfMAPuQX5
aO0cceYXwQfwBZ9/4KMVVJeuF9cgs/o9AO6DG8LLrqezEaKAEuNpJm0QXSwjpadedBR2ce9cP+Q8
K0E0d2uNquuWMB2xlBHRc1aM7DdJVZzG97yytPXqXHRP+8JXvCAxt92tuzGY+qlpnl5jfrDjsgGQ
pCbBJ/fsQ+iu2yxZ84eqARfWcl+U6WbnFbxBMKGTc0ZsVIdnD4QIynPa9x04Ur/3nsYNDy5/Vc+w
xIv4K2UnTAp22Vu0V4vtmgFi996Ix6zLKDMzQ8OSn6XMBQsAUrJIyvNc7JzCh7CXxhUp2xIapm4U
qFGiZmPpReMIKAADxvcgS+ED5JfhXIiZNYshGZKA9lTWrPWo3LT7M5T4iUkgqxbJdbSQCbw+GduW
s9kXw3KAtdcb/MIpmy2Dk8VyekKVYpiCHyJqla7pjUspjCXCBFTy0iuWF+zc9KOCGnuSUDABUBRS
n7rCMYX/okyavFisw10nnj1Jui5HiPajd7jxpJLsbrIOfkLZ3yobe2d9LWENls5cV6mOLOHsiSYK
3YQnXeqlwQR8S8njcg44gvoxoYSTPLWWpiQfgQKNvEb/DctES0ZsdGMMD8mgfCgK0oJ3YAARu67v
N9ByYdC9mD28qE3AyrdnMRl8EK58U7tugPHasg5NqJpvDP2NBwRJLCaGanPIjnDXp1H/WBfeOiW/
9WrKNmYMB99ZwvD49EcihnPZOIESgZT7S8Qcd1/raZiSeQCxJleOzZSNiffmn9WIZeeMr4vBYB6U
WuFvx1xm8Qla+7bSAUmu6R5mikjEHj+FSpgxGiYVBv+/vR1tN6sdb67s3zj4KwkjMwwupm6xEPmx
L9X6t/qJibhpc/9lPD9JyqCuYy/i+sZ8l3xQLVKk+E8fmBkfnoRtGzqGZU4XiVAJ+umAhUjr9+BL
W7zsC1thGZlIuvJRMR7cVDWz19fUVhUd3X5YbfAkIJW0XN6ZwZg3YZgFXL/xX2WsrTFLXCrZ2yc/
uWX/T+pEy7sjH5SNdgxuW9Z3IQr94NqoWLrWjkFUYKgq8beur0u+HjMDr6ui3LkmUj4C3FWQAW8U
zB52zZeW9ce5Exc/hBXS/+fbglE7IyLdYqNhgr6kd45cEZy43f9ROWqzZ3upcrwzkemfjT65SBqe
6JIOb0jmnnvhWKnWjwtOgZN/FxAN+SlbgWKT3UiJct5XqvE3/fupvU5bprqnn02Mnej8ICwm4iTX
phOWDhGWkZGILnqUs0wtsrs/itW68oDpc8MSSv0ZX8zsh0YAUPKMmwdpFjSDBXCnwu5kh6KD/RHh
Lx2A2O3rPIn5v1acWQzJEW9iE2NElHt2Iaebd4XQ3SyuH2XO/iQ0WQrLxauOy4zhfM+Tc7ZX7dxB
TrCBP+VXYyDOIskbRxMw/gQfecSNBm3gGKZ4EUFSJYYCMpWINlZuLZTh6R/Si+VEcrAue2NlGXcb
OZqe12oIt0bwzteuyBnYPdcMU5A7YfRnhRg7Bik6OoOuAzA0Mf6k50joxlf/NhX8SBepDO3UJZr1
0HF8gLxy47RS8qdOV5dOvdvx/GOoQTE6boQsx15Ss9BriHBWY6otY/CYCx31vO7XqlIViZSaScuA
rGNKYoKb1iS10bjHypD59b6c1sL+5HgV40BRhgRjZeE3ezp74Ua5cJslX0fEqsaLuCF381KFDPDz
NJIQ24civb4NmcMECQOHGc+QeSDj3xXrkSjU1bbT5EA5a4kYyXRRkLmjlRitjf8P27e2d7SSGJsH
xRaEkYoOyMWAYILA26S6eoWqQ97NfWs5uN1HxiWdy57eGdHjmUlNA9eZJc/VwEO52UoQ9PPsIMWj
RtD586vJIuhIUt8lVEj2o5wxhwS78m2w/C+M9F8IB1ceYel0jKIQ50ol25jFd7p0V0x+walW/tSh
4qRVWqr8LjYPZlL8+JT5XgROie/MJWCjNOBZDXfFNaIslY/ver2Ate8upQEzTwEfixOoZVgZsein
zkU0cbM2OgyEUqXkJKY5O4NjqjplCqbrDZtu4n3P+hLFLFE7IgrkBAYST50WOoofPcaKN79D3Nhm
m9B6Tro5qDtxACy2imNOHqH8rOlD6Ti5SxqWGDPSABj88d9yh3Yf0iy10pbbVbEzpl26SuA1X1AQ
+70oFKvsqqOkhhB3pr/0y03dvQ5WuY7uKkCvkV/SkA1NbdU5O0yPtKrrCxt58jUm5GRAFP+DlgqB
wPv3JLphGq4e+mfr+TQmYimu9kkX7Sr37STv/GbjdqCQ1giyQM4X0yMadtq/tM37A4IY9wMRZ0xw
dz7d0JiqtsePXH1wSz8GdxVT97zobzcMaNZDX264n808/XwJFEmE4hl91Tqz6J6zU5qnsvjNxXJR
ag8QJVf6FT5yeouSlau5CnkdMxknR0cAXlHsogTv82xsR1XUMpe/G4aziGcHLtNXCb0e25LDS32O
Ug2sD2bfycBM8wzT/+34/A+kSnCbUCGEqvgXU2RTai3HGuKh7i/uVJM+Av/GWqqaihJpOjTTGiu2
ZxWqFCT9HPqOAgIfgllP3ANZAXsrX36CIjjwC6HhyhDRGF0SwfeiRVzWksSCTeiuUEs1ZNMvLYIt
l1w/Faz9oQaJI+S0fA2iCY/0qollzb2whB6EG4LUsHC7RmjfftgTRCNn0rzGzjxrJGeujf3cJpYV
5YDuOadO2nPGNT0xYxd/lOvq4WtzF5U+P5yMfNMsrEMWvt/2S6J1RXk5NyA+Ndvn/oQ68eSs8pEk
6IHjS6p8FtGXSHsAlebM6XvLPnACcXmNFBZlbyCJEkKbH6gy54woYNo2bGSajtvPs05DnUSkJQ24
XGTEtSrKmHvkBMS/nbyf2plDvKjXwzn/rvZbZeGNfgU+FmrcL05S85hhHvn89ic7hixYVeqcDVpM
9xG22xexCoZbxtnizxtR6A1Wwt14sMLFKgvjxlUfgSI7L8MeGNwo7IF12kD3SHDs0qr843OObzsR
duItoaZaIqF5+I5Z+0Ym5rKZq1wmcrEe+kolrGuciZAFeU7i6WXCBH9SGs9oek8cUDgMVYG6JOw0
6OaBZ6BLOPjObg1Qm+C7EXxi/zGJcpDqCmZen/uuUiQTHVp+ju/Vn0YQqOz42rWWXwzz5Q/NGz3r
FwlAXmWbG+H2eU0uOh6Ww3BvK4ox22njaAIdegUNZ0ENKwgKaf2Js9o4bbJN9Zj8vcd7I4VyNbpx
0pzBC39+RtGqT1ileleph0ewqH3ftNTBpTPsqSuwG8ZtT2IwDFfa6kYoRYaa0Zo3Y8P83QDUKUJd
ZMIxQ8Ia3erT/XZTT6wNFSOvDUqdHUBF8y8dCCQYj8rybfX5/6LllqTG2z+lEEglyJGy50j6yJYR
/3TOsBekmAqfGbrXOLpKYF2kRb1oN5Lkbvw0aATUO4GjuRU735eQwEqUvlMEDBJJuJkoeqHOPYN8
p5AoW1R2oJKFV2f6cyeTDzsxcJgX3dAOsgKOstfscsoRA9BpZR25oLTALsFSo92NRba9JQzl7qfm
qO/Iau/LyBuApmybioVCZWUsl34MRWmaVNlXgldVSqofkZylhrbbho4QiDbPfZn8AUfHTd7DqhtR
AQRCDW39wSqCDhwwwKN/tFbBnW8eXnOorWy4uMRfOenYP9RiR9ytQpg3LNFSEvrBgpgeXnzCxIDg
usouUrozSXxdNyao9mnPyeRUUUmNigzPgHfwU0ugN59z1db9Sx1aGZcziPdIMAT9Sb42/I00ZW4f
2+DJbnbaje+8RCw/MT7E/3x7yy33BTpV64m0ig1oZ+WDPIasqbAVV0DwFyOeLPgaGTyo/rLEXs8P
se9sZZeHTy1ovyCFiwcrOQ3rHVER0uz5uFKhYjQHddDyKcWvC2+VLcsyFGlCfwmDZyg07ZtMrGoz
7C+nm081dEyiK8dkqHSSt92OZcxsfyxvrXxLsmsFBc1pu6qFsp69TndmmYrPGTr5hUu5u6NBP+1W
lultnumZyROIvx32l2C01USJ5sQBGH76sDNz0trb/r8QpmMFx8ik48IvROqUVmJ2fixNDN582cyT
7Xzaf0fEzKy/zR7q6QYH3BlObb/0e4EFm/XjpqVz600hQrUN6bLCkc60UL0kHUPiWg+594fBA2o6
xXLghMigTIhAw+okU4QVX2dXajFTxLvCiftrTvSz5aeG/1wVb47eduI9DplpJXpJASselfcA5QQ5
6IcJ8DA0r+ATuCGHVb8l/jXe4+KRWPzc6Bb5gBTt54q3Q71tYRWczXxtKp80dNpSUUhZbwuGtrTS
HxZdIGHsWTDpbNoEC2BLi7gL1rs8Q9WFXgz1vOMDBJsQOa8WgvZrWWlNRBNDBh9J1pV8PZM9U4Ec
j7F1puZkliV9kweTlkq3l1M7emay1LJ3+m+yL8CqNAuN98mcywpDl4J2obofopSNaJiGDvKIEMZ8
ks8xY6pzjqpbllgklWq/tOI/I1RVlWK28LOAC0RBi/58sdi5EPz2qTDTPygRNyZQo8LWKivGI0yo
VoiTZy0ELTr28xS8tfayqwHWXw5cUccwxmgFWvKuUfce4L72zhdGX0jdlmzdvGU6/8Ybks3TXtWL
0ZXUzWZCQfjr3CwwZThdTEVj5UeSX68/92Cw6llvg/ysX5wE4TGA8I42gBy+WQn0Q0zRi9C7erjm
mBkH6/nrn+gCrlZL+vrR4S3tbImjzeV5OYMpE5kV4Oz9SGanSMff+yqxoalAVueOYqgMt/xUamWl
cZAJa84AgR9oLhHmXkCa+vRCX7G9VTIyD5glb00PbKfpjRL0jhvUG/5P9zQCkCepKqlggZ+92j6k
sh+BGMNsyE4xkRD/AvKfG6fCUEx9tpHnooAWulezB1JVL7Pk5YNYevpqP0N0t1PmzLXfYC7BH2wl
zAY3UAwRDqSq6Abf4X6HE2NYVXFtPX251M5gxyFNqQjxbOnK3qKXf0tVeOjiixb2JbQM8fsrb+mr
8xWi6Oe4U7JWAJiMJHViQvKuJ4ewoHfglscS0MqcrDpc1DIfBWwhcLcLQlytX3kZPuetK/1SEovE
bHi0FoxL9VnWhRzqBWXOBIJ4ZpzTW+g8pZruTb3JsRhQfcqpqRrZMrFOWnLXo5uG/2kqUNVwZTTX
osgp/UAntvj1X+jecyUlPOpk8CQpIhGORxBTCSQ3qrhv1VtsGFneyfTQUfio3FRuKDNgJesupPbF
HcbvTgJP/tcRjvd6kwJva1yaNFrM+RqhFN3F5zaRgOHfOeuX+5iXHGCtOIKtPkpFArikKjNdVSoc
vGVRFhjt0lIlqzJK97K+t8lf6pL4guo9cIVjRjG8B5rEC5IauQktkSkU5tjl0pUGmlaG4HZhr6ne
1TlZWL7I5gYicQ0MBzq6ypNEmjL9+M2oGw9VuQJnR4720wM7mw+aRgrCWWkkxvaOf8/vWZi/dpGk
CtRnZOcOVgOzU5nxntxJDah3+Jo7h83ZILQ4fn3wzERNJ/tPFly3PFQt6oeC9u8lx2Vy9CcdFwxm
fni/vcYvUp5goJ+JdLL/Kx6TYnZeDM2oFNFRAU6DTY7+zvlmEm45QuYiZaDzr9UYO+U+chlWUjZl
i4+UNyjy/sVk7VaAaLm1rz21Ns02LHsSJtNv16YCavTWVQhh3ZjVvC/fyfxbZSSQ7daIShG67Bxd
OQObIFuCmjd4YQvD59BBmuG3+jO23x+ddf77vkTV/O2lbSncvvgLbyCWg77wB4/5JDxItfqUCL/2
6R1Id2TvQ6RzJBUJeyvZVBIcNTVgDYQQ5YPrK5C70fmLPdb15pr0N5E2xCGNhqXnhJCWDYbeSl2G
njSNp4fJ6ujTQogevEIg5ZXxk+3OX3xhPs7AmeD8cwj72PpHUyFOeZ+K6AFRBRt0jA2aDws96zhs
KRNDf042k02NIhXl9WLGNHfFaU8bmBUNCwWsSbLDXwD5/C1JULrDhwq5X6UeVh4MMI+COW7V4VyR
mZLm1GE+bS8TZUIsrws97jKP6raoWSE4FCIAy39XHmSOw/FFE532q+LdBINFFqtNOfvJhCwi8u0a
9WTO4NiMpzq+kIUivuzqxoeockQC/7RO7ifHVF570lRmcIXiKmX0iTIviK1WUJS+XXhRzBFmVAb9
CCd4jvORcDxRi7uizTM2jIFys/zx2Q35KxUpqcgA9/HTI8iEz8KW+moKxaReV3BIG7afeN2+qEsn
PzkmO6OR4cbaF/nWB3rg3vjAuQ8EtcgrqhrcGYwe8e3A3UWGZCxfNmrOjxX/KgkHGh7z8SRXGEZW
GYw5yqV03Akf/9n199NsuULmOUvoTAil75Pc/kEi/3yTxFH/RkyI5l+3Sb+UsIcHabIArHgk5g9n
7r8fsk6LS1i/6oQiZVCb3nOkycgQoeI/olbg266oK+jKU8gCDM59cajBShpq5sMFr4AOkYcQMaLv
06zClVsLPXuSOPuJLb57q27zuNcSQeowT5i+eXnQWA5JEG0vIAici+ncccuZOtrWslKO4kzvOY5i
vs0QYc7GwsCRrbw6Zsx30qT9vvlCaWfbSAqmzW1kwgMfF8OU9WyM5uNuWqknp5YxNF2Og1PMcQY2
eIY4KbV8+m7fviPPkvd4PmaAwLXlT7yl183ossWWxu4/d+gjkFa7+oZNu1mv8u7FVCXF9INEn7OF
eHiP+5T3YET5fL9/2xCK9evzFzY492lT6vIjkKheHVp96EyZ4zoWQzqs86ZIsuyP9E3XcDJ7oplc
4cDH36Ar0Un9Zqa3t/lVY/tKopdjsbE1QnQvd8z7ysqAvEjPsApxP9TFpQxJtSzkTVCjdzoWdSbE
RhndPSg7QudR9IQ3dmRESATbu3FT6gy5VxNNuTbPxd66dtNC+EgF1dw5LNDTsrgbBtH/PL6ojMuI
KmBrPCd46ZnJBzBbk1SQ0WDBZi7wAYxdsyPFsmQGq5ydREdfr8CSFka65EeAOkv3jSDrfOd/X1oH
SUZYftPbWUntTVZet12s4aVuTJncP6hB0CmCgwrUhzC6UxW8unHPmakgSI9qsdeJT5ta9ys0PxvF
jKA7luTXy8co9ZSZXdzQdnT6yXS1Mgt0fL6SgHFLb1FEyfd5t4HRjjsg0dRzv+/9rRdX3tiiYxfq
VSvhwXhebVN0TBc+/vRM/SNbeKV2mWM157KkKSBISsjKJzC+84774CJ3J9HMPajd1h/gW2F+u0nN
ZDfkzIbVzd0Zwu8T3oA2Lu7j/dvIGoA2Ae5CA5YZarZh2Y/LoZcqYRGMyxobRF1PNu6ChUFwrmso
5WXONf0VTkE8VQOD+ex0iztNeFnRddpmdxv2zliGen+eeEANU96ZfwiLVLQ0KSu1wGl9iMvsnzKX
KqpIHhDA35+anTrxZQ0b4xSegifFhBaGIXf1bw8PXPE5VuuttuNVH9YDwJE8PqbOA6vhyhurIYZA
RKNar0vKG2lbQZZ+4KtsewhKrxivZMLqoE057ps9kA6EfFvTK/lw1Kkz/J39UWKQ7Pl7CU8cDsUs
8X+6fVc8AOVbbS/0y20j/705oebMWiV2/E6oQbJ3p4/KNrF8rmLMVfVNl1Ed7VNP7RZ6AnDYUoo+
olee9wVCraQ2ucVlQkuCYWf6ezn9Qnf9EOXyioLPU4TufFkDUdUSho7zIQAszChRudULJfD0J5j/
O1rKTWChKMysFeXTzZFJx8h+8gBq2h4KkBF7J+mVb6O4wv37sE2iQhb2cb1+zEFPpCfnTlPA75+a
qVxX4+mv6tkpQX02PTefOET5EXYw+asz80LTKm0YeuO73slZuERkswIz4BrMmbpzgmBqYN/l8U8e
8jODIRm0ltBI89A38/g/MQHWwDkqOQJ5pQq8efbRdk4aTsdbFfpt7BiOciVe/pntr2Hk8hPWOofM
Z8655TS7/9UIVTWmpogxfAt29LS7b5Ed7YGtFmfAXhhUaHJA5U7Seb1eVHA0i9kBxboC7aO0SGUE
ZKhwgoArhDYH558qhAS6z8NnM2BnBfPc7W4H+uHT9ZjYwn4lXfp0APUuChUddeXzH90YpzS4I5U0
ZN0FN8604wRiCznc18YngZV64yqr9FX6/N9kAYRbm2f9IFnveSbTez53hcFgep6v889Poa3XEFGO
ZuOH9cSZaAufbFJ1EdAYYSE9SY/lkIpQNYtN7lweMTcMdxSd9QE8LRAZ1Xk8+c3+g+FwwmPXMV6G
wXxTNXLDPN3DAvGjgDet3nP2H8qBFK2c6CVS0Ht2nevTBlQHugdkegPe+qLiyWH38vSpw+MiOoRQ
67KBOIIglJvi82vqAatrzqzRoDeXuXoGCidPgYOcR7yWMuc/UOqbqipISVMfAHZxZp7iolttr9+l
0l9knV2xalko8Phkf5iB/0SQU1IeIY+zDVQhC9CQbrcqcdjZDyRCAAcovCovwwmeGEQOWHqCd2Jv
QcwRdVv0dKacFQihAn7NmgLsHY5IzB8UuMfGPxC304xSJffTjIOckPzg5A3qnaH4LI5Wlcrgp/i7
UN1xlyQLzqF3OGhaJ/ABCkO+yXqXX4INex37E3cqrbLpa2VV766ExmFN1FdL/pNd6zz2EoriLHHV
xu8zVGOTk2Dpgviz3bxEsc01YmvrlNZuVFSKrCc7PejB58rKr8RbgBdHBakBrvmZYCT0UqWZ7vGL
86bRxduxNRRw4gWX12p9MTfqrpAHxSTKuG0xjrk5nea53d1cXwP3bkAFpJ7mluXYq05qR1evPBqV
ci9163wQa6dxp+WioB8NLnmCr3MYZf1Tk1P+YqNrtVCuq59Xoux5L+VRcbc+RY4/qyLoMla4SLHx
rcEO4jzArjZcWFlhPPAb7t3mw7AJye90N+qj5oJyPicd6cFf29KPwe7/YQ6iX08keaInxl49Rr+O
sxK8vKaIutbq9fyxUgd44dqWNo9ea0Jf4yS2yPGA+4BMR4Y9Pv5laNFs9uTJWNNxFxjO8EFLtITD
e7CIIB2HsrBqX/B8ZfnpuWC8Tb6h1SVarJGLUTfDto/zzU42jiqZNJjWcUvAg8fTO+o2ux3V
`protect end_protected

