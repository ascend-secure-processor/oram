

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P/xlcjJwX9s+lRbxifq85nCZ+mgGAvyLD6WIWoZKxcA1nS0F0NwLLZWU3B4OXUZU6YSF0t6vRPFF
mzlKafs+Bg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f+/bEb247PSbYNmMjfJLqmwJv6VpC+dDE/fwQS6bTTu6KEySaNh2a7n3ZPWIwdlFtMsB6GJxSjEw
5/5BTw1i9BvSAx2d+8ZQ3Lo5GG1Vk4dTJ1o+OqnP63cH7L715rHBjKakMXWMjSMFYjDqhfYuDu2A
GrH+9lAj/CZwKSUrK6Q=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vIciPaIFcop7yWOlf117qKTOMDeA+0R19+UEUAP7uX06ZMRgR6AF9Cm4mOAOyDFPWQ2hzMDnfwS5
7ODwVDdWIIm/PEroVa2PoSJ3YalixKiZHY3/STHroQEEmsV7aphXGJThhYPuP3+nRo5lN2aZM8Nx
smgCmDeL70m67flis2XlFWhu5dbE4khdk9SOb5bfPqXvul4ToPT4A3x/4GIbsujiCTnvf01IRc4f
nh4427WsXMjueN36F5P4iXM6sALRusteFCZuSD7EJzPC2hmGOs+QnE4RvDzplmEuSquG/j714fQX
PFjjJ0KZu++rZxozY3TP468UagUxoNtuNfoHaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YVAbEnJyFFlPl45LBlZKn87g7Og+C45oPK+Dat1+IPasApeIgL1YGNyyJAlERBXc3Ec59+9YYSwz
P8MReitbPpwVKvE+75EIp2ZIGRqBUKDimh4BMGeVCi/U5TRcE9KTzNR/5eiBib4yEJHgOcJ0rIuC
LH3sd0v7YfpdA94aeyU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VGlfI5KhBrPK9fz9cY9PImkZY5i+87n8lUERM1HUvHB0Se0jOmSfciUzcJjCqEiz67W8Deg5jnkf
4hwhQJqIrr2SbxW3Np9OmGsqeXhIufZh+e5wE4AvAfYyf6mjLwMAvIq8ypvk9LT+ST49vNAkBEev
4g3naEWky6lj3b15Mer1MP91RZI+jxLL3dTujvprIO2yM0ycprhiGCppPnLSI0lShJW6AoGybj0t
yH/Px7EGZ55p8CqXu77sIvpnIqHi0LVozEI74whmLGX3unQ4LWLAP5csWHz+H1SGxje/KuNZcozo
FbHkfyStJ8IgzMFP4lICblbLeb6UCwoSd/z/vA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45184)
`protect data_block
92Ckizd0uIEPsoGpDaUsMSvC1n8oi71mQnijcvzr0/67wyiVlIcC/2XamL7aNCCIUsjV/JgmjS4Y
qWmRkxtdaN1H9Vw7JfPgb11wOlc+NBlUSaqo7MHoSXaeGwH1so0mDR4oRsryFSC1xXm1P6L7OxA9
yo9FfezzPi8cTRc6y8sUM48u8a9lZXSS/JK5cE7uciJesc7xHZDbii04youm2IFpenRyCHc2dqsC
dP7fZZMe/mHrts1rD7MkbRHEO8q3GL/9B0WT3kSBi0m/bOjerbPeOQzLRsvWz4MVimrvipI2nABZ
H8jUiWnYrgOV2O8rPToge+ZG1iahd6xG2QbuBW4O1wq1Sk4GHts/m5vjNFreIF8/1YVVVTXg5LNz
pZ4KE1n9lkACvOMasuNCmjw2OqJNJYjCzW8sh4Ng45mIVN4Z5rgFPHhW0sigDlnXMWrttcFv3qMJ
E07o28H/JdFzJmBBYArUhwzeMidDanBbgKAhK2Aa0aVHg40g9fb3dANV2arWh8Md0g9NvZGDTWda
moGMKTPyc/CyecuGl/m4ViwgELWhdRSUu8tciupI08BL4hTQ+NFzV7yIh6zJqU9wxjG4uRWrZVyy
b2X84npHWmtINsyW0uGnIQAfi+TA9Bwq/OfAeQP+aujl5kqZEusc8JeR50TyuRFcZ02BnOb8Kj3j
W1iuqFuMMI9mH5C6GwS5zvzY0g+dIgYFfgMwv9Aij5i7MPBMO6WaHvlbxTpxD5rOfeQrTAYETDi+
8o0X08OTanpnnHzQ8PZdv0v3bI8oqCFnEOdSYjc0jTd0I+WpjIRI/OFJwvnUDqn+lFyF5367POlq
vzVxivHxJ4r17ybyUvZgLRMP0EXDPPonmSWvSknLDx6eZVGEsZ7KdQxByjop6jDjszANhOjzsYA+
xL5aldiaJkWA1oZ6jomTom+Krejtso9tunZsjjF7FbjUCIr9M3E61CEHQruzpavdY0yu3F1m1GIG
yOU+jIJ4vfhNdC/XW7AuaFHOKSfEUfTCidd57vwve8KdlDZLgHZC+VWq0DOy1cBqpDeWYs8VuY+L
uGFViVRJTRQrGIOjC/Og2KBKwm0H+SGiqErV8sJZzhEZu7Q+l5fuzJYhAG7Kx7vv7o5RyUDDQS3G
scrf8G9sapaX5SPmj6NzjjQRqnBFbBBKBxbqEWvHVmsmiDg3Ye2rjKXrOPkWknRt0X7ffQeb0z0K
t0WXw0O/JXvG9Tz2tv1eyxfHJiYkjfA0E74V/yRl6GoGz5FeiuVKo2GSOtHiwFA3LpOjtIhl0VzO
W5dsPbQcUEE/mx/7YcZsHCgMLiLoYhKIfxQU9McafONcRad7fq0PFgnMkaeBoHwX+0JoW3yXBwoS
HNrljSSQZfoj+Laj3rPc7HnzaEAwNK9o9kcxWGIcoNIFh+ZOWLSnu+iR58lfXJzyaK/Vl7rEPR9X
HZXZdbIfUTBtt/EES+d1VT+L25P7sv5N+CtsWwrzY9y3g3slFRSTIAIq0CoBVoOEjQMj3APZI/ud
q+vEhNwb/Yle5ddiArlPCYIekI6TbBRPdUo3AZFhWpDIWn/b97lF6eEgXsrLECB4uJZUVIPMTJcq
TCu5nZsimqf7FRkz+V2gKSzkenbUVXF61l1Qa8D0z8drLxY4ve0di0pWDAh4OV8beOha8NM2Zor/
vLe7p9RPosrOtuvznfLzocIXsG/65BKpxbskJ21i4JCrVVM7va1ZGYOXO1grUUP7gskqCBJZR2qr
GVURfNzypX7izjMUcNDZvDmZSqhgSWX1ywBO+kcPPqFIbtnppBPNQhBILQ6tRflpAwnNrUwA7Xy2
EwDCvhSnLhJ+ZeAy0c1vRzI2yva9N5P04N+++60kL4Wv7yTzZjzd6mY/HAMNfr4hsEdq5i4LXqtX
Ym/q45E5W5JY279Y/VrJIfE4NQui+skg0Iq6cvZa3Pm8fODtMrO3CBr13HTAX7AXIgmsc/vrTlD8
wi7NB3yvGOTOrlVY1D6e7BY9HmTsfxzrxirNuvKsCkCa4ViAWQZQTWtNZQacqn7CgHi/Th/IA48r
iH1qIX9u8FL/qJlKBLeFa8IPxDw7IQG3mT5JcHDbvusRZp6TELKFh5ftaN0dXRGnNRTXMQFgX6wv
MKCko2k7GR/Q3TZi3IYzrSqii93dWB25270xNe4mwgrEs04NsRfUwjRzW93Srpf2TgE3qR9UnQkS
P53VDtvROjLvTogEf4a7emEKY+eiXt0a/daySa4JEDqYuG6hT+Q3Bftz+hxyzmdls0C0TM3uonA5
Y/HUt1E63biqa38bqa7kSBic4GB+WCPao5NziN/oKwGS0fd3Mw/p2O9YLjt8uFVuMyWHhSvmhDdm
03y2pH/yb8TCpw2QUuhsr+mfdKOx3lBMTrRa6uKzkJAyaiV9moMjS1fn/Qkvp2JoEkrtV74cLq7P
7Sfc3/TdWfT7JL9vRJbgZCQP7zt05pWwFKr1GwL4g+g82I+X7RhEasXrYOB+WcwCRLkbHAuzFizC
bcNB5vnTb/iYdbw4QCJKYKfMH/LYxPl3pUdU3MCO0pOyy/SUgkaEbVtJxuortDrfSjwjNFfdXcc2
4Nx0/8jDudN3K1twnO5FS3/sfcBdoPXdxT4HBgJXL3JZajB09eE1wI/2VlxKWqjswAMAFZMOMGaD
v32w1J/0xZa1f8ihyQyllLd7kdg2SgW8pzqeA/KsrB5d5gJrFd5T9VScEORx4hrzO9BJZBJZT4C0
zKj4KUlhSL3zT0bqJjl6yMO1ellhuFbQZ1sv18/nUNW2Q3GJkxgtMW/QTvnPvH2ZHZ1K56KAuGZc
9+eyHmSr0uEqnNnnLcEeBsC2IHmRuHshVY+LpMyZlqDC2vIL5Xcd3NoS+Tax8Dfs2cJAjcpmHIpH
hFOyP5afimbLyZn1zLUQOpABXGLUID6eSImrecc3vOVAQEL0OJPw+S4bBy0vxweTg4+fmA3XU2Zv
MfZsDpSPIL/qYA74mq/UTPg5pJTA3ZWBTaDri716yjoKi/JtdsBjMZrOHp1CMT0lL3nq6Im6iYV1
iKTibWZLMDYcXZw6QGct7BU5yUAA80c6LrEGKnjMO48j40zQFiSLKPikHWh/w4NkSnRIpeLvs1zC
kbuSURgVJfPGDUVIugO3eXB2OMbddH7amtrNWYPJ8PEnszGUqmmTooc1PR8j7S+wFSPLeEzjnsKs
HzmcMm/n2vZvlVT5n/gI+w4dF+c6LJDj6Z9IuBAA0BQiX2q/dtCMpxdIOdT3awS+qUewkwTuP311
rn/u9YCAzeFdiYs+cdh9nuFtLBAxNKsXfdGvhFDnJyV8+EtgIhJB9wo0qi0WwIXj7tFwu1b74W7I
YgGnwDNCrnrOYuBNIdd2qKUqHtWJMPevChPOHtyI9vmS0xdz3nw4ESe68tndLnRAOE/BpUMxHRe7
xw9XkaVsF2T+UJvirEpiAgizxHZkNX+doxomwmJDB+Qvg+UJ9/ZC5U7rFgy42gXNZv5uZcv8aY3B
M/a0xk4MEXc5AmB3/De5gNaxpGMuFho32ycHMTu422d6+Aocl3KuXL3PfF2pbUPBeqfei4eT5c5K
w99f3PEwkO+s1XWkqOz7AlM4KrxhAb12qoRP1+Z5U9512+SzyaPmv2IiiqrQGf9kgem0NSv9/0S4
33gEXfM4C/ctMh1T5bnPPIC3spkVFp2wy63kbf8X9TAXeRVFaXlccwZiWQI2HX4AKGYeisjJ/okf
swFeWAKNhpvhMdlRidVxp0wYFBRshR3QW5GwFBFt+ybrVAt3lKnxZqee8nE+R3A1mFJE37+Xf+an
oi1cujFztujAcTvT6rkfBLajz6TCF9bAojy+zpk3+3ChdBfHgBdvDS5ID9epOZjymDNrE1+Rsu4n
vPHACzexHgCN9IvaOsJnVNJrLOvr6mPTgzwX6oiaJLXsRS6ZgwUEW+9+rpOaV5bWPMeVifx+6aST
86WDi+WSL65SJTMVx6FoeZGHPnLxkkLgPNGW53fssoU8ylBRkI7npF8pewRZBDbd15Sej2qmXpyl
Iizyg24qUnG04mPC0zCc85T5/lgxE9egEVAAwKqMH72byxAcFkYiUDeWZ/CVqIVytZHMBnw4Eysu
dRyyiY7U10bMzwPrJNO4Ev9ftSpwy8uJ9A6r/P7BYi2XvMrkbFivIUOpeoKSchNrx+hmXfYlTvT5
oecE42eXZGRxsGxQ+XPoNDUx09HHZ2n9gXVNLhS8kJVG8i8Tdbun9X+shPxgg0xyIZVw70r6Imkk
MegLUBc8NQw033Ca56/5xv8bp35WzputHktasxwDOaMU2pwuiQVMOO7zb0pLW6rcMgA0DL2YDnDY
3kFjp7NVV6x66RUWxdN4t09UK5j7IW7cnr37n5Rkpdasb+PCqtCAS2ZRFlZuNKrWhNHKOU4DkWms
GRDUTwnB2SbVO7NQ2Y7GNZSNdpK0BmDCoi5KFGXFdzf8q1dth8tbjpwTgvlOScXZZlB7aA9ASWzp
GBOqPWZo2cdrl57bmFHP+VE53S0etejJ4B6l+oVCmlpNKtuC65vo4qltVTaLlG29Suj4Ng3RNOk0
/631qELiGtKK7/5rcjCP9805CN0Im9pjZtu510wGo1nWnDvGMN1WqJKRyMyyEPOo60lcOQomCo90
0hFwujguAORud2nR0ACtccZVadHPfP/SjzTAabzzguEVyluSR9YGXmMjRj7vIREW7mCUbAJT8+1+
Zj9dqD3WUNcnKwPxrTElxfW3O+1g2bO//CwsQ4r4OCqlEaHPUyRnQrOiseBjbFkHwM8jbEaL2P42
ypzqbNmqy3vf34ytnZrPYYosmqzM8XRJjV1pjREEL9GiYbS3vEbIveBBeasG8WLVGklGnh5IzacG
4pBMH/TqKX0uV2CDOWM68BfrjiFsARpd9I8TU19/VKS87mm3UuiFr6NSSErr906hAqzk35xQzwNe
SqGtIgSQrr2Ai31XyQnMTgywX54YJsLYAlWSZmx0ojgATa5ceRc3gjASm+jCyq4bzDSwexJiOBHV
V5TZg0wINOBLmCCgeAOIw3bQ8/kTJU2mILQi8RKOpR5afBGLXSX2PBZhKM+1ImujXmkySKQa+btp
LLR11VQd3j1smzOl5nV+2tb/suGObnfboGFJrV2/Ai8L5l1hOIlA75J5G+RFtAa1GSDqZ1DzYKaC
Ysw4obn8+t/SbO2eu5zzkMgsHkvbih5qbEy25juvTBUXeqy7qvKUazMJMtIE1kqed1oaHVg72xzZ
Gl+b/coEtnAZ62VkaHwBc0OvnxINKkkIgfgtZmoIYlr1cL1qtHneI9d50RwJMG9G+m4l1bsr4q2h
0skpyhJlwMHhPC9BQLluEXqranbd8k/ga4jypVR1ODk4ZcGgXCzRNyHnTaBaKF0LVWsX+aGev187
ZlqgV+cvPF/f9ucFLOUmB1NAvpANgvU3TRoXXMuA6YwXYS96YX9HJpf1FFxoyqcQVnH7tJ5emLg1
9y7gsC0UUe6G+yB/lQ9b8swjvF2aurl9qkdxB7rMVhl8kybxDUMK6jnwRYv2jXjBcGmdzyrfcSwm
Aanxu24mL3CVUJ7w/KG/2EOFTJ6CuVbceJFILadW4a5sPtmfgJpPwQjgkIyu5K0MBgLLbS3Tg333
Na58iA0LE0fG0jJbiE3j4B3VC5zXFOLaEJWi8UjjKt+D134+MkVAwvBykxtycQ9C3obeKR3J6T+8
EnKDlza9g+CLDSu72xFYGAp22MFFcDhnUeGxDSaJWpIaDD6BPpRy07qB+NVmxSaJx59gW5m1Cm72
vRqyAxkykEvyenxC15zPt0U143YNuvWztqNp1LxH1HmlqXnru0aVnyaJ192z+GiNCCo1ZLQonweW
BJx4weu5LHj2XiPV7YQqzGfOkv3kN/UPvkBsSMo5qq0EBFBh+/BUcf8kM1ZDKRbSrEy7ae69MY/3
g96kiGaGPZPDRUNY/32KgEXfSyBo8HMMlT6++fxxjS32KL5gN2H5MDUJOQ9EAs1hcnZt3GmAUJnl
s8PkCY4apXTwxRRhlT075whUWWawdAy9czt+8sXppxb9Uu8fNnQm4NzppRvvrECz8RismhBOJ6ni
B5JxJmgHFWzjuVbwStuTgpTnLjaGTLy6c75C7wXUJU+tIUDvP5pDsa9ntibTMmO7XVo7S+B/x/Uj
NbTpo5ObKV8C+B8QULp5hAwTpCFZ42R4vQPKpuOIDziZiaGQyhjYIortiWO2D9uarC9Bpc901eSf
ACa+UEU1U6aJ0bjY8du6URKaTzm3U8XBd2lDLgnI2V95T3kgj/23RMFrugcKMIYSAO9pZ4srdV2P
A4xGm4Z7GU1y8/LuhFtVoqYY7sdOIYgej3FwQH02Izs8LyndFYQYW9W0/CeNKm6pYHLygRNK5Acs
bx80aXyEqL5KAGVuveBRV+9ACa5TUBc3C94Pp5R2TjsF6m0okL6DQqWueflRhNSQW27z9ZAKLTwJ
wV65jbcDiqPsvDzynPLHkmNU16b53n9hSgQo7nr6EUKdhV5LzbbV2DSnhK0hTdeRYXOUGMQ6X0Gi
PdddakPiG9I+SpJffRI3t/V6csY+M+qKhXHydNMcZj0gQRDLj/2O9t7nJeJdxNg9GTw+vSv23rlL
K3Jw35KK4ekuUvrDyKRMlLEMv+ehRBbAvI27j8z+csYbYEX9s9FWjl7K3VMyXfaKiGhB782aCHHG
ZF/VszprtfoDB5w8RJqGAbFgBrFy2reyXCOOsUb7U9sTaauuooe5Wfuzu0cnrxHAixSakMW2T6pC
ASXDLLo+KppC/wQieYMQzJd2B/2Qr2Af3ow1LOYF/bKOMfSQCJ7aL6UpIFgr0iwKDTWz2AYK89+6
0zPOc5xnsiNlumyKvFBTGAvDpDdOI9ToHH57hMm3g2uRCb255IAssjKwqUlqHhGXSY6k7p2h6fA/
AuF9I6aM0cn6qBVMkpSdO9EAJM+SxnFn+B2I/vNcE56Xd6+oav+saeS9inszRvqfUSsWAzW6wMRC
PgboZEKdie+F468MaN8v61uIzNzjJKWSMF3LL/gY6BNCAY6ZiNjLjaXiuN6YnlHcvc4+nacYrQgO
akTzStobV8SJQiMwbRyYnOZu8yh0u7BWqhfNRvUF2Jz/jj+CXYt2lHjRXIu1OmUn1XHbtdjQYRRi
G87gAcX5A097Vunm3uNhOyw7tTZ1Ryt3Z52eB0qMVyklspJTU57i9T0rzKNveXKXwnpvH4SrVT9H
yCYx5DTf5B4HzJTp0NGccvU4GFsYEgcKpUbgpjCORObJE7Netf7XYYiclbJ2f5XDkc9esHC9eC5y
uTDYvb4KtRxxPVoKgttDSB4CKUoAhjLfukXKLM0IU2bygnaSEFQ5CGOddkNx0Lo/7VIMGSwY6Fj2
hLpkAeDXlhAem/Dh/RkrN+HYq45UeiHFHHSIRABgRXgKgrSu0IqxJ+DuyPZYpUp/BcnITuq+HaPR
WtC9nSiAezPpy5K7156RJlRZrZCg8NjiwkHSUivjdPiUzRbQgxmqWE8dKcI9z2hJWq0HPDqCLNms
3IBwOx5FW/jK+0HTnaeoxBwM9r/4kazR1EuAZEz4ICjUBFdFD1/qrNZw7o8CiMWl+HGKpkCXJJpb
gBUGyi4GoPSwco7AvfjazP2IUnOQm1e28XOpQ1HeLVuFF0VuMValCWV7Y30umznMoKgGMpn96IFL
UDFZ+hODx4o4ZpelKxjvfle43zznxn5bD+FAe6gRNpFhEgzmFSJ/dIP+i6pTMl33dyLRFNjMU1Ap
l0bVQlBNXTdj9uT9DNil5HLBo1bs9A/NYMhXREVHrPEn7x0lONU66e50BN6xkeLOCv/WbcQJ9Wn6
3bbaBfwRfYJjhVnt8sOKfH3lXo6GnS156TjeAMQjE63B28RO+6G9sNQovp9siXUD+rhBr+rJCIx5
ShZIgjl5yr1Lj2xKvXv1OCRIphYvxxHCv67DShqGogpTKXrtSRODS0RB278ISeNos2GiKW66BTH1
AVHbdKkQbihsFuLsoRPDhJuhdXoGiZjteXraGbeoGiv1+OU9KehC81OyLpoHAJFpUfBCtRC7IWoz
RPv4EaJ7IX2XnPTWRVmiCROGXPvALPdfcF5YaDhrNTuAqNy82AavOwVqVhsE/M1Q06AE3IN5EYUJ
0LauR5Ss4KlkMYK7X/YB0mIiCO0TFgSHdypwv0GQNC+l5qezc4wPpeTKs86shIB2Rn0BIFTyWkoJ
dCuj8hgKzOpRF8bmRtUoDKAZxFnl09BjgZcimk/eSLxDEx8EFufvSmamVXw8unJ1+V/RKsKQ1K2d
50kpGMkXWL0t4391ormdiJhAoo2rHseJmqm1WbPHD36fx9OoJkhGVvFYC5K0I4ZwX7ArC2MuZAaE
kzIQ3JFL0cxnWS7ZjnzZYyBAD7J+VbGTYNxlAJxaa6OwUWxqfGwgGHFG3FY0xv0lawZ1I42MyM2q
tLgC90rrI/Lm9fzapRqniSqxEI8Mw5fuHVfSp+28rP+jIGQqUoS4E4Dj3Jq65jXKWz4RQszTxd5N
NuPyowC40s2bOK/WPLo1FyUumGgQ2KTRd5jpm990uwovwBupWQ9yT/9w+KZ0fAv1MPfs+qMIUoDL
g5lIsH2kYG9/bzvLyHFXc+F5q4JLb4+kWACK0x78HhMPUiswvDNhvHwHtJd6xa1sgkV4vlq1tC7w
8tRWM01cwLV99S4LlcR6WqWHk/UPXArFpdZvz4aQM0pp7ZlOCNYbxp2CFYo7BiPjziT8gEtARLqH
ikP5nGH2rd8pKnEugwXl9PSfjv5z5ePQozxkNRyYl2Zd8mKZsl9zhUbqz/iLoesCy1MIGAKDQtts
vsyFP2dkznNKA0QVwbtAQJbWCVBzXfKE4bsl/mm+S06UfVP/i8TieyjX0yIFJLaHwEbo/A7DGjns
FnChD80qgajvcf32AZ3QSkFav/8vL9+di/hHfMPDHV+ae9k6rM0N6k9n98E6YzPnAxYYrzqxkzoV
zXuM35iq6qa97z9wiltOMOba36J0E2GvYXlb3PFfUFi8pw36T9jmwhD7q6tc4FDYBP0ItPD41qrz
cUXfrq2f6zeZJdxSDtL0tnuHi3pVRPTnSAGp6hzUVNicCJKdIbI6FhFXOeRAuaFAA0A0gZGjuylC
4bcpk6c3AmqrEdTNcaf4/HZxTTsEb5N9QRNz1i9q4t/0isRFeOh0o4EuW4jOsrxhBo3MReTjn9t6
PMWfakAARA0stJmdbw+9wXkihXp9W6hn9mzLbo5jUKHLjx++ZoqhiSBEZ2u9/AlJEk1oPo+Gfyiv
tAjhf0z9RIefhSojdToiJV02dKWkCSOTbK1raKH73UdsCOhI/dDKUlZAnK4AJfL4G4/KxPDJKX3E
6somXveB4Kjyz0WE3dLWkzFcXMWAZFg0P38K/gUeTmOmdpHcs3acUhSCeB5nNga8z/8o5gDd4dNr
JFhGk7LgjxGpQtk4TAPXbLnJ/BYESkyR2+KnmEPdcYmz25e/EBTmJHeqBoh6VmYrKWB5Lm5z8o6O
ORWUuPDr9MtrBzPgxJdln5Fuuygy6GJMIlkbHTCflzhUorgXxlY/XCRzYtg/SilEw/EWJtsaYOqB
czYUE/O00guTe3wgEaa9mQxi5TodCr2JMsa4py30MpX7cdGzR4UC3z7DMKad0D3dofmfpMmLOcYe
74djvkpYGJfWqiql0dq7r/bIlHDkmCzMBS1yoMOtgvTW2P+kLw4Ep3nxSjIi4r2fnWnbbuH6izbz
IMNUHQO+lC9gnNAh9+h9RGYRrngn1kpoE2tln7UKRx/orrubRDBlj4GvA8sZfQuC18CdEiY9vurK
r020yJcHjXZ7ExK01s5G6OJR/bzhdU2KgJMXmU8Jm+Bw+X4g+TJWz0n4zNcAR9cLRZxULVW07xtt
dGbWaLd6kpcx0OXDucW5VT1XuTyHGSsLietS8+k3ec8jsUNYVxsmCM1qKwioN7inkdQ8VXvj07ak
hRNFqKkq7DNS8F5b807tmqvRFiX8lZlPqe68QGoh05tUoVZ5+yg0go8Je8ssSFCz/18IwSqASTze
2QbKl7nkPVUwBf1L8GW6jdwqHjL5BIsQ2zKM/wpYt0p+PFFyf7RsitIIjifDCcrTdc7MiNnx29lQ
SKRPw1T6nDLG+fsNwrma3pJ1LxcfTzlkh0gNPvbaHyA+KSb31RYdRmcahHrh0kenQj3YTJoqTzP/
Re7rjIcyqu3FckVpWPlYdP8+w/vZnksj2OIeP/+MTFGy+F86mb7lVOIv3F2Oq/FKXqCEccRXnoq+
n6qCHxG6XhpNxv2F1RTNLLCiF5fm9uKA3+EHVyUaO24tFqiqIBDnwciZwFmC7++DSxPDg3L1hJ5H
3cEDYa5aKFz5DQMh5zA12OEHZX1SSLkvqgN/j2SQdqwcoGyLdN8ptH+2KFBxgD/aCBlRFW2FIR9g
jZl9xXfK4zY2tildlxywurK/Kr9EgrUn2Q+miPQSWM+pQU5J+cVeubzFTErV4G0ZAsL93MqmlAQj
OeDN37AfQsWfejx++Y3wman459O2FTWeHLkY2Fl0QewQWvAvsohP4jrzW7VIy7jTcIYKqUcFO5Zx
TlzSBalHWcqUKStaL8mkZAHBlV7H/bgCxWEWsJeaQufv8ZyY+aJPKnxsxUHbY41Cv4VODj0Ke4dK
DGAmMgS7DeU8xNtSCOTDggFQeEzYwbV4PsqIh04ypnWmDHPLGM8e9wYZmykXAXUD1DBFFNdvL/pu
sMI8F7hTmd9dRUd4G1UG+TZY1aiTopRp/uj1bRdWekEcib1LCqHt4Rnx5Ydf9kbJh4HvmXoFJ/ED
aT4zPqS9gby9GDc4/yPfanrY3W8rX+evklnKFE9HRM9ciYDN7ax4zm+FZ/RfUiiab5Iv3EMAXe8+
XTE5ghOL838JAxwI9NC9IlQ97XUOJ2JKmXGOsULCJUQ2HmD08x23W91YboBgOcaX/ql2aD07FpOV
6QlaP2GalKGbevRDVW8rYMDNDKafuBDQosS7RzoP/nWVTn4+bNcdpkB+5msH2D5zbm2RY5BmV8hP
kOeVzUVXGrvjWPdC7kzKDDlJiKQvB4vVnV7FKlx3WUjfu508e+JAXx+idPLF3oVVGZ/5oUUNDFB0
ogXR280k5HcymTY+grGe8MYUAoLz7CMP+FHYIyKGc+TwyOuSsTuAL8KPDzDVKj13Zxd2ROvFaWOO
vnxKoTnN4MrkYg+WlfmjxDsSdjzC+87+ZD+YfkLhqLRTd8KMEPMANNDu2G0vcly/vihnW9fxIQw2
9YElAJ5DGXB48mt2SaU4Il497yeBSRLRRbuS6n2E0Q56L9SkoF/sc94qLRJ/aGhhV6Wz1UaxVoxq
yqq0p3pzKcs7DO4XC1WeqGntniFQ9pkUjB71/lb6zebvduxsqGKF75NUnK1LT+qYTI7SPWznokKl
uq8YPOPwyVevfj4Fg2BTdH/EY6l4XJTMQLN9PBYGEbouZdjv/H1Z6rMvQtsdtDj0Zfm2tar7BCZR
q+CiJhM7EmN5jSQWgcOoEjHnXtPoTMUX03fg5Z7JwOIa+B9g4N4wrqh7uSwPsGhZiFDLmgYxpsUF
cTjOg6BKHmFJQlsDMVJwhZjPpVmdSUfrW+ov2+XrU01ZZY3FkxyS2vfGxvzj7vLpDU2OAx6aWCLG
2Ks5YTzjkSEHpBtwPpOhlp79qwCpjjMkA+JN9k4zBk5X/+MpJKMyAtHQCn7qc//xcFEP7tYFoE6b
4DQ56iYGC/AoI7Zhosw/LC47UAsxDXTTBrROs7kPEEz4ZtbmFCfGqkdcA/2SRrzLe9p+KIHw7I1A
RruZyiA8C6lwYFynfCMXD9TTgUWVdaiDlTLLH+jvEghw5J45m6Nz5WvDsReivjUgZ5mOzyBprOal
GY1iPMzsOm9Ez9QxG5T67TBpzfWhYkNRQWK7pcMIeIc3NAvIboX76tS9SqT8ookhGG5ciObr0/fC
0KNCuVbu79a+PCo8nxP6SMBPnpNaIZHEO6IX68XyE/hF3R+5QVDAKzaeFvhH4x56wiPLGXnMbkSs
ObrcHNQBBV65JIc1atjGcV0gvrrG6CN6BJxl5VQpXSCQkzDB0k64tzVfxWE0U0GRTX+asa3nwWPw
IOAHOa5RNioHnK1yR5ddHUTRvYNpns5tCNkfkx1FnJeV+505j12AOWizEYeCA4wY7AggZMk0nK4s
rdmieTew7wh8rYJwx8GWEQOPej+C2g2h/AouwH6pPiAj1m674ujFTTyLUj84+eH+QhlG7OiCmbMA
h8U13bLcsukgT6HwhtsjNSExarpCldiR4r7Qw4f8z+/JYFy4vuvsAONfvrV8aMePwl87NxAml9xM
RIH5Ix9JDfpm5HU3y8htc6xq5cN8FW41KGtoOGRq8N1tFYS5XktWOx6JSGzvskuBEb9kY6BFAcVV
R1whIaTTRoNpA84y40B7TW50T+cSKVknCaLmTbQg+DG2YLRBC/w8ra5dq4kbxFHoXirqwWjkWkxl
oUkHcg9BixCMkpWoin1wUX9Hu2Eowql2DenKnzu9oJqYuWs2CXIAVw+X1GOhFMqG6LsLQY1S1FDY
EdXvO33uYR5Hx2UK5R+uHgQGtHUmnqSpkj3MkTta4MlcK1/dq0Fwdny4y2NAUScBofdW3Uyx/32x
sJ2FFXhebIUFHVOyRkjzb2JIIIb2eGyZiy1yKcj8UIHykOyoL73BEKDT03SV/p+4ucngWHPpaPLH
LhI0duFdQLpQJRQqwRlPrMYI1BH68Fs9aTWMmUYcr3wxEkFhs8w/Vn0gHUHUX11VwiXIQXBMkm3W
jpb6r0uN3uh3hYtLisq4UGKsd613PYhWHNy2pBUlTGs9SpUQeNvzs1i4U6oJEFalqbsnbWrrNJZZ
RQhe24IE+W5wRaDb1yXBL4t7Tb0uybipq5mIc9l91G3hHNOVR23xcDXiEX6t+o3DMuDf+++UFS4v
PmQn4kyej0MnDkuzCmbF4f5429FDAh5iHEtKelKe5Mn+FBnv6ZbXPJlFrrh9fOr13KxS29o5YGzt
2P/5+y9M0lNhZrR43G/eCzhjxTxg/roulh9K8Utlu3oOh7c/cWDy3PTg2iy4xuN9bqcvqfh1UwJy
odb0o22E/hozUna9Tk54NlsaBnoXSObD2kpykYei2gzOj8KC2F4z30JZkuo9KvhHxa0CUuyx/Sn5
2w5Pp/hbl5m8ExZ1G71reePtY4VxQ61hJmpVB5ciPDmsEky+/NEAOO0UdRd5aJH9mF0OMcwYfr+g
09Sf8DhktmMZMbmoPs1aZJgz4Dd7V1ZhQNzrfzklejsYWtMQ/jC49a9hP9RDcbl16P0gNDPEsIYS
X4+9kHlebkY16T7pRrTvWJFVwsobbKu8jzpy2pGKdu93RQPfhYKMds+p6kt3N0SZIhz10/aXpBdK
HSUgGjynkcKc18Q+/yci80bO0FfJV1fDWa+uEt5JStDWFqrnH+1J37hgmIT208i2Xc/peebLpTGA
qQEqq3CQDjcZDP8QHecieWuEpUo08/1qjqWaRvfvTX2B2HJ+pC6DVCb8TAUZVvxAl36HMeC9KXuS
xOE5mgDRW2RFCzTIhsG0EAgmWqcmW3sapYFAUs/mLv/D9lxcP18gO1rb6uNRF0jw5VkVeurU2+lG
C043hp6SRDzY7N4Dx8B7H4OeUHJC3tfSx8myoqaEowJvDLozanLOQFTEKtXZnuNbKL8Bi34pmB3E
3tPmBONztROLW96GAeBbxMv9c4Iws5xjqo+TgU5mCX32hfWyFNlqDTvRhbbIePHK8i9BP/umM75O
WSlS5Ynd12p6eqKiTZT0pr5mbWfVOVQ89R2TVtQgYmV8XSKpuC13tMXruZa85mIngNiefYGNuISQ
10PYCfvh7i4YqtlPmo7+3CrVbQnEWRey1g4rluRWVfYc7WU03dkZ5NbxnCZBypJ14UImWJcO8lr0
IxZxr8SIIL82L3vmnQJg/hZunZuzxThJ/AV8FjMvQhZrV7m97GUx3RUiGlGA29Ewl277K40/GP+M
9OFpZsjbmBT/btzggoj3KzqGsjaEfCCflaZ4wkI7pzi/tQcMn+kpkePiHVf7qYX7DCIWY9DZ2BJi
PbtzoRbdCyNDZoY9L2sGPz6kfoKHIwTuKx7LdZM01doIxH/Hk5w6kFwnU3VCyfBh6VBf9TlxtGV/
qFjos9IC2FjSLqxv6M9rjmAdwgvzaiPP14SN41ouUJx9a1ZekhxhJUeWsJk5ArD7AdINtG75HeSB
PgfQcPsggdDAGAkEcZThceEoUhzElupHw3RHoyg4QJw9XQaObHgiVUeKRyqNXEpbeWB+2Mb0zRs5
bcGnCVjkdMEJMr0IyaQdteQPKWYwTmg3bypdSeAF9JTNhf+3ueV1Uc8Dtd1ISL4i/pEq9ewjYQSa
hkxQX97Xee3qrGdN4d7yEJXID6Kbjf0kdSYfVfqISRp/NsnFB4I9XarI04eMI4UlzYbNlwabNHQr
EgFZT4mguHPFo29Ty5cMMhZfH0ho2j9RgdJDYcTWCe31iQXp049XIS5g2Fymz/i0gGdouJ3ZfeKg
JXoDXZX7femnXVCQmj7yXddcqCmfxTZXgWZbX9R4hjMx5M8svJWt2RvhVF6H17xkDwhxkr5SF5j6
AtzoqpTmVHv5vgZJEY1fUncjoXxCtZTG6YN+c2FzKB16XICmXjdKaUdH+GGsWuqBthtCe4JLLgx1
pgx+Y91TRDVLN7InzUGqh0iNyqSsmEiPwAaGALQ+YWHfpnMuu3QFpIrI7wvGbMDMppelP/KtDDJm
YBSm2bPhk//0Hv4uS0s6k7YHLoOaMN4h4Y0r+hxNflNVgbh03jdKUS1/6rurOyyG9NqO46iezSwa
yfRwqwsALbwGachL3rNy+0bt1wc3/L5+Td5Td5YFCaITWzK1hmthyY2vp+z4NRToCedWX5ps+ZqE
7WEGPEazMN1JG/1LR7Dhq6//SoHXRZFo1v6X09CvKYpYbX4LaHdw1LyCTdakZlVwaZlGZpuQQ8Du
lnjDPDqLudhA/TtFf65W14/LlNxElR1mDqGLUSFV6Y9khPzRn9ou+d6pBnfzMSEn/7T40C0ShExc
MqvhJ4o7W8OVRZIaoJjMKpGkPlvKIEyAqk+fxH9mz55JwmkIx0yJWgkkAn7S1gmNYiBqdqFgsFcL
OMKbpHHQ+8/W6irGb942snniPgtwJgSAexULd3kBAq2Vj/zpGHZC/ayN7rp8KVYYpIULwl0Z1diS
JC/R///0fGSpgFMxsFgHJtx+Flc+KChHK3icNe8u0obycIWHryW685M5MgvLissO9Jmt8p/EtmM9
UPKKkLP7hbppZ/v+Qga9kalO/0J8FXioZyjnVWqCs3+JblHJShgNhgtRw0QySaugHTDg7AQrXO0U
xwZG/2gYvL76WFjDPZyyjFfTuO8lKnWSV3w5iWefZGhJIcqLBj7bC/cYyOPELNKqSqYunyvVZDRc
K540ZDpRLVkIuog9Z3zuZQkwFyJCxwDgLu1M1l0WgX9s+9Lr8oS7NALKcREDSNzMpnmFMKfEHsmV
sNbpXfapLhsIGVT0qJHuh9DV0+FHL6QRrRlOs4dOojVpdGefWy/Y+hFf9eh55Eu5sjNgMp07FPGx
TSRlRq6HV/ByhWOdNoghgxdYSKr/ldRxnukFQxGtTXFGeycQ80D6I6UbBTnW0KNjVxKGx3wG5LzG
Mtk5AVLFVjUdhVfR4zbSR/7y4WtTN/Xt4SaAXMQ2mS3cRWmvSvIiqZSFnG3KUiiOcDnmYcgueO3g
0ZDKURdyK/bA+16Pvpso0JLLCzjs25nSVNiZxjYOypvSq46ZTCfWGQ9Ly1e9llPJjCnBspXWTrg+
3xgs9ZRA5ZbHxtPfgH07wjoQA4oh6NHb0pDUfR1jLLkyIy6Y5KXyY1J+fJdnajcx13w/LlAQuS7X
DR/FvcFjzjoOwb+fD9DeHpW12m4DlwTPtuGuZu1zjJmt9/NGK5YmSxhc+ImwUH72XVwGI7bLQavb
JQl6U7giyl5nRVbkskkDb1OZxCh06rDpAIQkRe5ORaX9YkU3bOmV8uFyiFLlig4lmfic/qTw2osP
+QwqVLnA7JSp2XmFhEsZvjdzcVPA3p6UIYagY46eOHvewqJ7Ek3UAFZprdiOeITrqcxkv0g4Bc/L
8bYt1L8DQcZD4KNuNNpw52CQG7b8x7d4eE3sZgjyIasAM5ZurFE3DAL27REKSyPdhZEW5HM/NLFl
x+cx5MKikxeVIMGzE5fb5ZkPO5Ir8Ttbpz7WD8vhZOeCzmsFev9Gz6u7YdeVsBwzh87HZwcd0YYU
k6oORwGMfaqGliDFimogpTqTSRVxlQqtyo4A4UZogDIIx3cm4EItnArttNRIpU1/oY68Ley7d7en
2OwsDUajLquY7i20VlYO4dFiUhnupdBGl2HqN0gxRT7LlS7hifHDtT50M6XxjYg8mNpCjOCfSRj1
LBJXyRP2e//7UooQE1jkLqxfCo4Am2PIGrJa9PSjVdXbdwBmSUyHY4vi37h1EUQ7tZONX0OPc1ir
w0VwnK2u6/83peS3+OTw1Z5ZIuKCAf2e64KrO5fZ3lDWXlcK1RNJydCJO9F8/AUSb1KrEdLAbHYv
cwHkAD+cMl4D+Qfgdf1zkCofnalRwY0WXFDYtTBWhxKewqPC6E/UUojnUSJMTTlMqnwx3PbnLXWA
5dQQeXCVmwdFscn35uDCFz8OK0uOPSkmgqeBAOAeQf+QE+WTkso71LzEMisIUCz48+zt6DYb1xGy
JfW5PwAh1KnXJXXQE3eJGLPtyAnU1FHgv6OoWPL7qaJhIbwvOgFnJSOhU8A1vl/mWikePYGHpgeg
1sb/I3qOb3fnOkWTaGaHUKwBQqKcWutTAz+uQ8lwRxP1vG9z6/0g9Q8Z/OmqO9vpHHY0pGBPcGoc
lqUSyW2MDu4ZR/Wq2Ktm4k2bmzI07KcuYoquuGOl2p3tkXrZOwGrdp7uZueGZKNO38lU/Bq5Dn10
3ZnT7jSi54hAsu6rF8rSHFWJ63nhMKwTiZ+2ol8eNzvb9AAF/pyuX37ag/YaMVn7BE2gYIWNurln
gpDbx49cD2wM8piYc31UyuTydB8yOO47nON1grKBqToUd1vjROgfi/uGQQQ5+3uvIcmkP/HulTzc
4Dp5+WRSk1t9LB22tY9wiBTdB6ogN4CZzTzvEP81JTHarEDR0k694ElDSBhO6AvUTR0pYMFQSvgW
qr95NLEPV3bSzsAHEqXIs5FARUD9tg1htZTsGVcZS/MM4SZvO7DPcvZ5XKQZuwG9nXq0RxIIj6Ie
g3lPpqVsohOXEDQPwKSb/COSCMxsy44kJo/nFUA2XuHX7d4J161psa2DgPnXQMtRAdA0gJPa/PoB
LiO6MXpVjrGNy+JXEk/tPQmuWiZMqtCRq/1QhEUhVRtWKPtaAYmDpUyETEFp1iZGx9priItXMf/B
qY+FUtRGJOSm7yM1h7u3wCwkUpwGNEnGMAu5liD84kGT5lUlwVnwlf0n/BOD4F5H2JVjFPX0ZuVc
6b2qV43jzeF1119ik8WFF4BUb3P4TSLPSVRDjoYcLDprV5c/wUmkh30Nb8notVl1oTWzMd52ebq6
AObFae0zQTM0oz0Kaw5Ue1QONaWB4Dtl1pgKbScNvem1LrZvZntgZNw+7I+lqgtrveY1HX2NCThj
EUTwOHSfe3DgH6axQWPQyvafcE88JwyPr405NpMy6H6OB+nB5VfQ61WtO5u9wfwmR8DIi7H4v+KF
nWKRVjhbk3C4ntQnVQTbvcqy/Q26Td5xDNKqGAmOV06AK+YFiV7SYTrCsvzg+gWz/VoUviCYeN8v
F/6fjYulppfAOyPLZfm/l5u37/ecERDcbBJDM/Xcu6eXjjKpuuwlzcmNGdat7hQg/KhssCD8gjCV
UJWku+/3Cg6+PJtSbW5zzYn/4IK7tf1X6PxoZV41WzieL4CkA6AWQfQNXAEaT9djyU6Yiwc7JYES
FsuNRD2rUw81o1D4ysB374gnzv5f7TShgxV/FbZRZpNw27YilyVOjKMmQ3qKj3YcHyRNpsEQEdbY
P+XHrmoOjlfsXzd7f7MQKSjwZiQcW4prmVUXyFG3Msn3Hmcu7m0Bm2/slIyv+AJ1B4rhJLWKBgZO
WH6TYTOJCovS2a9qoIl/ZpBWidVe+MwvvnfeTVt9jxCf/RKrGfjG+kIhX76YjBAgQ/ID1xhK08tK
5ftTWJdboPDb2yETyK+9MOcPO8oFoWojOpq2eFZnaqzUme/k9AjPAtOWorqXrxsXPa2D04I3MOOv
eXfVXMLz9HjkSSF3RiyaH5HSSt6EUhywytspuBTRZ4KNi6XG+yKJY0AVPEl52ArVAGRz/giGY/kO
3FOMZNXaz5BL9pZSRNqVoaV7SQ6SIngJrta9PNSFdyzz583adjTCCxQEPrmSIzeP/TfV4EOBQ+oS
FY+18mbJ25Ji1hBYYD4kQOX1InfFFYR7NZycOxcOdI/OdJpKMOIXnbszdtEZMijrz4v3ziHNXDaT
5KoWq+Pd2WdotRSNw+dCIBaQ/jBbhQ8mEltr1OdKUBfmwmR8r55IRtm/PZFFq7HKSpAlv/egOKHO
+SaTDvFBYCY3J32CcNaxSRinynoUOyfqkIBrkatGBPH8GOwurgaj3kSWKyKRQSoemtKm/dOBrHPb
lK5XtwB9iGZda8QvnX4lg1h6mupTiigZzilglEZBuZvG46PF4jiriGE1FBLTYVUmcheI+6dcQU+O
I0d4zoFvWPsJOVQDk8U36Us1dO6TH9pNAjyxe9vhZ/HKS5N1Wq0fNaPOrAGWA916VtqunBr+IbRQ
5dp6LPnO8pwyYuYOt5I3/UaFbe7cxKKiYjXN6LiFJRw7Xd2BENVzRl3Cghfo+ZenjBuqqq1GhO6C
TU+DJAJ9QtML4ZQxsYiR2fvsibRIe92A7Y3SwO7TAhlMq6kgCh+Tj6b9k8uxWj7BGHVtpttM7QUM
T7vlzsztjs6xPKBCnZ6brSsFN3c2Sem8X07I2J544Trv+V0/5X0eqQC1GimkCzQh73hvcvSjs47i
0gAih8on5GXBNwc8RfTUtKTRlgiins97L+Pi8kaYe9qX/wAcaWTaAzSO6tPiUC3HElSJK74wpuUA
ZGG0hwmFFC7fW7TzSJGQC1gm8F9ZCDSJ5JLA8n3AXBfTUqCSXzeNBIx/Z+WCB3RMQMuRheuOMg+w
a2jybT9/K8u6nZ7TTpbT4MKjZY/QhojH/oCB7LyzrkQYjQNY7jRtDimfi+LffCHPnZUlVZQ3GzvP
4Z7NU+mWaosvI5a6MJt9ST10W2Otw3Wd5Q2EIDHCNazVzzgQLFCGlxGZfHVrlYYY3inQp6fmmFjn
VNv3O1mDmNSgsJwzi2XXXOnW9n4rzt4FISVroXUbTCV/Ypg58f7ex4CNxz1stOnkFvCimaRnQHoJ
EJTNlu0BwGLPoar4XAxKY+h3UbrmcLefZYvb3D8HAX6dMuzavQTXOzx/1i8rRcbgNeeMF8YSOb2a
XNOzkh+ToYct8/vKSuOxv9rVq+E6LvAvxRf7HNwMNDLLRtPWtcGmIX8uJfBNVdn5KvkxKhp1Lpj9
j+Skow4J3RMeX885wVInnFF/e7DfDVzHg0KXWiOw2WSeRwpapTYrfcp9E28EEKfZ5VYR7S14cs9W
1s3su15/q+YeFqTXFNaGk8c1dhy5wzIjBMeon/EDXs5GWwZ9avyJC+aCyopV2ehierl9OYYBn5S6
0v5oMLYpoCvyP0Sdb2xRayT9N74MWFGX2RbC1p43ZMOK1PAtdBowf85SEbAx3W4S6HoE0232mdpp
2Au8eGq7JUIaOm9sMAPleOKyNTrJSZXg+lpTZpEg1V/8q3kpN8tlX0I62PXZMglpbhbdWBF4AfxO
53vWCCYGWOE9xW0eC/ySFG5rKBYlWzCjY5ta66jcCn0AFRC4ybVGDSMYvfF5F8bZedXff9dO9PYC
EPqrD6y0obW5KYBBk0EmXpOcAFgpKTtDRMT3XB/SYvWcKDDlJCDU4lwKU9T5OuRyEmW21gxhueSN
IJXt92fdtJ4yTIpRqYZ/j9IDw1LUwk7pIBXJwF6A4UY9p9bHtZVv3wx21Ws6TqahLsRTmJxmBJeR
T4xuSuOePa7LHuJbZMLuxZ1TlXs7Bf70dc+rf+ddo1L20SrxT3qJtzIn9eVJfFTX5eKx897WodaY
gTxipJa2ee2LqNY8JPGoOIAZH7f+2kxVthWDEMJt/WgOLuimV+yGlC+ECmRv9VYev03XEcwAF06+
/yRKA7nevuAt8m/V9gSjtvabe6P45FhTN9ODD+Yi45jB6YDtXroWrs0Flcsx9l7Are4FG/2YvESA
JrQpjCe/YC4d5n4i3ln4yBXoWNlvpYRTM2PyPMIRd0+bFMocnlqFuWrq734fS3pwfkszSDJ05MIh
AGigF4E9EalX9t1U/+CUg2KYT10xUw/5wTVaM54O6DHkYW0qmgnssln4EgeqPaWhOGuu4HcFg1QK
BfM4fP/hSWKFfrXzOxhoC4P/IluZ3y7XlFJTQifz7Q24Qn1IrPVG2wu/2jJbhjd2VupLPJzaTuf0
B63aKxiuD63WGO7UXyhAjfc2hrIrdUTwJ6cEhCgk+apwrxqXVrOXeJnzOBHP9GnECpNs9w24lYDj
KnT19L8lME9vk3By3enCL8XgyED9Ns3MOdi81iKd5dmB5cfWNOXCkqBdLbF8dbiJVRHX7knVD9+y
L5Jh00+hxns11XpvvbXdwkqowT4MzqwxsKoi/A9kRfX85ejQYoPSlt0xr+h8Q1C4RnltcoKKxGtd
TJ+xX3HOuhmlb7tZnGmGQFdgbER6DvwY8yYSrPgSeMacET/iXIqAfmdFBihytUR7y3yAWI9pTuYv
egb13PkeVUQxVycQw338+Vw0o20fHy70zcfsqsyJHNZeRsVKPJpUqfr1Ch66KKBbvW3j9K4n3xMi
sYQB3bkDSqnF6MjavNxpfHnFgpe4t4lYZt716wc/qMNjvAv7qwTm0rtYzuTvE5XtUewBqtvofVzl
Bn2MlVpo3EdNafIdsyZ7zh8TDEv7BSvR9DCq6WFE+467SkAgpLqQUwxCEyDA7fZtkhqLXQj5L4UU
UiaiVpXGInd29Pc3y89SOeyqWrn6EZpV/IYeMKwKWw0Yu90oHdUd0vO8hxKG5TdZN4XfKX04liMW
HL1cS1TDNC8oMvub43rsylaPhPcWY4285KQH6T+w4rgUZ6k/lj/zLsugFJdMIRdZXjTSipXKEM/h
Ksrl+ooJliSJaHyNRTgFcWMkt7yBqbgd8l/w3Yhpq6C+fnIoDcgZvvgzIHVFchnYx5MGWasmzYwY
1+hkpy7hqN7iDV+HMjR1VJfUdgM3NXds8vU+kj79M7lWXsdptqTt2kKTQA2H8pY+BQIrDcTG+tI5
gBUJlK3sENZEB9bAqyjJXuIIWgjTZVbs7f3rBelMe/iOcHg+u9lKZPho2FAliCsX+o74QTFaJQYI
R4GyBFdUwiStqmaizdmoF1cE5ZAThrDPDsbFKECKQ/dIXm5uK3hUA99dOUqjrK4i3WcKNPjsidqo
L1kFv2cnsly5oWFUc1CCEDG0oUQ6IAzdPDrqxp2+Ja2Lu8TtqYz8fgd3gdlahVjAn/AtM0RsVvcX
IMjBEJPOnn31eAdgxrTMpC68WRAj1Eu3UNnOFpPt5VgB7VViOjKiVOlZozSSMPU+DWBYP8yrxL2T
Y3zPp8Q71ItJ37BwhiD++hSAjXC1A4n3rUdo7nRPieiSaod6cqaLdMJFSSYHvvjCVvKaMHOZvaXO
Wb9CLQRQxLh7mg5oCv0devKx0LSZ5t9LTBTMl0zynD9cS0mAUkUufRgZ583k27QsK9LFxobqf3+S
urSm1URYnzA/UBrvT2IQgUIFYhFzyYJsnXnHg3jUmiEhb+IVjsurfevym9qaQI12dus35bDTa8RI
dTbGsjNcuvppDRXeyCc++djWLvt7tIEde9BiKSiV7pBYu5C4gx+2H5awCpZAThBL4hBrdQkyFFht
ein0f5LXVqNM1jRERlmmJxIXSQd4tS9daKKHTxIJm3FgpNIxjCuulECbNXX0Urr3frZ0DZWmpOxM
fTixAW0nue92cHFsbmuQ9Jn4Y2sIfXG2kiVc48TOQo7aKSnkTQAEPQKx8hVJAL65n6iLgKHrcLTV
0UeE0BgAXjgGUsk4GsIfoLvq07bXv2Ub4A5kwiBZsm0MUIbqlIKcf7FF1ZcUziigSGNIrPBqHDGQ
dzO9+S6ksogCyczh9duSYrLaFpu1qwCTi0Acx6bOcw8NkP/PvVCRcRdkJ/mcFGMJoRKzkeqZbzZe
/INcR99bekellgwYJXaQRh+Ufq8FMrseJqVakuuBbCytVvoQaWvz+aFhyyuGUOcADzSCWwYEFqX5
7P2je2O4i88dfSOC+00yLl8qZYmFmkfyvFsHLxKBLuW+YNKc32KdQ3CXOHS/LMUariOVYp41irPf
Cr0Wwdx6bbOypcex82ov1VwB64XIBYJdHNk9ybsYu1CDwshO7MTu8pQf1RisFMl7RI5i9A8Yx4Ca
GYhVJ+jcBKiCX26HuPI6rwpbBWETy24Fnvl+SEaDJeSSMPIvCT5Hd2kOPxjIaN08Zumi7ryFDaJO
yn5iXH+noT+HxMnZ5VXcLs4cRaec/7T3/cqdBF3isf9rZOL8317kQkxVgU6cURdYDx1uTi6fEZcr
0bA7Urn4k2g+d4kHU17P630ObUWvabJ0vmi5wEXKn680meRiN77uTA/vLiWEsrEwhvvjrweIDY99
pL7ajVK7h2q2dJRpWqNpdYeiClP4JWTMOGplSdN2xCXOHf06K2l1GvGmDlR29Y3Uo0z2Xs+Dt7HY
fZtFEFIpxwc++1ZEou2I03HBhTgVDlyfq6WUi0K95o1+TvwRbY1NH/REiAhy0CnKr4CTCGzN7P6U
x4GDIV0fcPE+buAiL7PTpKwA86au72EPoYOu+sMhZDUUetJiXRnjdMeC4wsVdaVSKuXWapzTTxfP
L5Jrl84fTMw4OYc0aLXXBOWlBlzMZ/9eIMWzMAc9eTcFax2wV2kBv8mfSy1Q7jHEwO5tkUVIc7KQ
y8UJCUCin+Go9350d2rjTufFbNgDVEH1sSz2ZqL7J6BdvqC+4EmgNmTDv7dQRZBWSBbzEs9429dN
RP9YuR+b8becURAkrjfUT37IsDUf4HLoRYY394JecNgLHiONEPL8iQcifGDlJ7VUurLR7FHTbPeN
rAghqgqPWnTVJsxiGdcYQyYGMScV3TE7KUlbbuxdLg/io7oEO1xDzPOP9Bf/fG69mJf6689RJGWQ
r3o+p7q1vHu171OI/oYzUCFXAriTJJz7HAiQBCCInIuCjIiapPJtYBGrn/MtccwDvnmvNph4Uqy2
1K1c3KVU1aSxmZqB9ciiPxAFbkHfgNE5x0CgTT0HDI3D+03abKhsm9eGNz3y1oeYnu+WwfTHVTXx
Oz/Tp19w7oEy/5+mM7JymCKfs1LVXOymdVD165TcrOI6nP6nXfCq7sU7onlk/q5dHfeYHiB6RqE/
nJyKlYnHcxDFQMSLTAAoWn2VtZJBYo9YZwor3zyP+CwPhcFesxJHo9OST0TmUp+o1Mlcu1qAQWLB
TayapyZvCJiMJ2p+++8u4CBOonWMNfEj7lPfdjbDmfmbCttos7wWh21ez7d3ytUm9IjVAlra8D3T
aftorCFxlEYJx4J4XL6SdzjEAnU/XcHLTt7HFVQdG5UCkgt831RmyTZlM1ix1VFXPqnKxBpK6SzD
r6TdZFAcllBxMgvfYBstx+tHBuejddnLR83KgfZP20ompOtOsSpgqg3HWIdSR1QbhyR33AvX+nCh
8MFs12bK4GEdiBbTg4ILFo2CAnsowrDAxuK5IiP7JP3kDP+Q/f1e8EJdLLk09wPEKR1sSCPYwjoA
vGt7O2CHNBKwQ7lrzOTuUeUM2MgFYvQJ+FXsAToIv2BNjoXfmVI3EqInPqOoSq7T6/BybfKWGW0Q
/5SHW+xC80D5suVniFHF4VXl6hq6yVabG/+4uKG/PqafG6Vy5ZnXLllFVEGVVU5TiibPcADE169f
QseEvJHK+lDCRfcB1+SQHAkvYuCu45C8iUJKz9GIjgAJtEJ5OTZQ1A5dJdQYDncTHnlGDnUiKvzo
wjTzxPAaxHG44opEBmK1q/GDRciYhBb11MR5clF0suJEyDdpgqqoZe44AEYGuiCxFEuxra6V9bUM
1GVwPbQGtQZcOuPwyRyXuETVMwm/XkDk2Rk52VxDtX7YdneeVbR6rdcZSAvsH6C+Vzghw7Y8mYo5
fHEdSpiXIvkd6AqkEtcWiw+xWYSjknFzsY+GqRk0pQU/yu3gpLlrNzBQEBS4EMSPh/IoDkb6IzXl
tFzABBsqgZLoK/QuEjwaHI8XrrLYDS8czuA91o3i1aRYmGsgGqN4z657bQPeEwEvJZa39zvlXJ84
wASOfMyS7QoI2SYkAL9KO/qbbWs5cHj+HNyuH9NzSGxmrWv3O5rbk5/N22S8XXCIgR1T7dhDaFjy
j+CaAcRec/VvNnyFG+O5vqFIpYmvnUsDoMi9L0Z38ppGlDW7SBC5/4bQEV3UMlVQ9+kVVIbv9ewY
M8ydBcPAdYVw1G0B+U30N5tsUPpgNchjwivcIBo6MzMxmWV8FeKCI1v+r1s5jJT9sOpRju6LAAyd
YMYrRSIq7xUMT7sX1KlQpm8QYaewN+jbhdd/BtKqKXJ8WnDVLJOKo4HBiEWL0uPJZ3FKxQLaTWIb
9Aw/pCDqKZcYxwW5UNT/ie9MLQG0GukuhnGGFeP5ylRl9ujVdyaSWYhS1s/34exZ9xpfcpuUJ3Xx
vItrtAXCoI8+GEZNhM9+FfM/Rc4gRNZ4hIBFUi3zUg8y9SxjbOLqDxoOP/CP7wskD6TKeHDIyMr3
vOpWjWUts/oMBWMtD/SaxODRINE8O6RakY6QerV7Z+Ns1XHn6pthdQM7H97U5lzbRphYfREB3oRc
SiVsz9KICdP2aD9z+obpHpjzOPRJAFb/IEH6dKDtVkIFRvL8993VlFwAgHHvGkOTfQFJ0oJI0Rjh
XjQPLo15kuN99gzLwXOCfXFYoPAspu5nZR6rR5VEEq2MUL6lFlT66ZUXCYEtQhRDGpCpEWekNUUO
QhvotQ5KgzfClfOt1d6dGxPPmpy3B4Zqjg8VoeJ3C9uxkl5tfILxLyjMJqL1pdgkxbDajXQvgGCN
51T6qJE+PjUPI8QSUVU/yJJcGBy4ZWmrtNhNi3Iy2HXmprxL1HpnbdE9CFyktyBGDKt2qkyMFwyR
/iDcnwyVn0uEccS6E2QxuKjuiWN8VxKIgSoSYZxCwl5Mxebe3tlFGaz2DWHgXgOtW32ME/Mc849h
JR8YXhcMV6x1/cKO8UbISd1xQKgVXprEP5eNqfZGgITX0jm9nfdH+bw0UfeIl5Zb8BBlAcpuDy2W
f/NQMzXeeWQCHiL2AvC7ossHVX35rbGRIEuPDjw/UPKWhWGsca0oZuPhrcJcb442HASPPLzFpwoZ
HLbIJEVAd3dX3JoZCe4tZAh2bQHRCgbKi1yzv4uxL5T2hnLJisYPG1byCCKjeJo97SBn56T0xcsL
eyTQnbOhtIL9H+dq+/SztzAWQhWuNl7fmp8rvJaCFkEa65/pTnvT3d08TmsOBU5Y9SSZFb3yuv+q
lbDrLpdmj0HaWFQv9UNb3XJ/y2UfskGst+iWMr7GqGhnuNaHcEObwi26+1u/fiU6juyXN01Tih6P
0pJLhsf0i0krogywJtTUt3t934QN3l8tt0w+/jLQvDuS7Whb90oqOHqeZaK3j4QUswocszF5uVqr
eAXKd7dwLTUSxi3Ar2H3ZvGDQ5baBXI/zBbM/U87NTcc05ke/JLCJwk0w9iyPP4Eg4b0AShUqX8X
s/M6GnkV7+yWTpxFDqd4vp3pBSQfRlHmHv6MQUiqaGNvYST4M0JbUJIbsunuM43GcoaN+qlLukdm
zH3AJH2MVjiV20a8G6URReFRqhiYpOYXmI9PD3681h/scx0wqUjH/3qdCk5DvPWZ8bPpJ53a7gcj
+lUraJVbYGNbxqSXzWo75jG1ZOuY15L/R5vdIbvWEsKyDT4jh9/4Mo/u1UZ7xqLs5XDctbCY7PKQ
eHMBqtm54h+dtmvWjCAcpYrxd+2wjboQS46+3qkvvu5vcA24W3q1dFKi6kuOqK5LWRYHYd63sEc+
Bmit7kZrVXfT3j3AVE4KxF53PhybZHB2abYkFYafdXv3yoETsVHprTxFQ99TI1/snAOqDO+M8eGr
dBQY60sCo3A981uIu+U1B8kUXtoLopMsmgJxnuncUXX2lR2VvYQoJKNV53zVyDz/Ba7NotfrAkq9
nf2lODufkUHg8FUawZMUC4zpRbQRfbmV7LwX0wlDyvbEctgZpMDBh56VLjztXxzYbCgOoY8odz54
BU5w9HbCtsiYXlMNPM6j5CdTxsk4CBJzDbFXfDELJ3hGlJ46Nbpex1Ebh5SfsbtgD/XT39gijE9R
tA2FejQeXlIGb7oR1C2SwdvEjVF7iQLvfmHlj8eKm71ylfKZAiDMJpKpxumTo2jpJCcOCN0//NoO
P/WLPRoBLNR0F2AalLZehD8m27rfMAKC5RZtTxXYx0gf9afSEv2fGZOWf+BBYsrlw1JnsMv8phnN
Mqr7bwXqFXnbXiOP7J89W1uh3G4qofQLXnVH/aU5ujOttwEwtP1ayh2R0WEL5P3tk4y219bYZ2pf
5c52rp8IUKVLfuSI6OHJisTmXM6US+26TtHJGtS4Ufimkgv09lnFPLUR6l722S2viQpiUBmtZ1Al
/qDP28frOKufsSwxgquM2FEXWUNX/+4wrAPi7Maj5A0E7gFhwJhGLFieEzkwrPGnrOp5vQEs9L37
LdAUfxrLVa2ftEPv5CBhhgx/PeCM/AYnLQnBwdeYYYN6DsmHQ5N4keOVDExAhn3IvfDiLBRtkw/z
A4OfedD5qlVDnbfA485ulYIhvJLiJJuLFQD/iNk0s6e/EZb6tiMRBlIF6xEJ4YzovHYN1HKUD0m6
xBh2YZ7B7g/wguXdkuAS3G3ic5FEPIOwPdkqKnrIwN7Hw9ASx9q1FqttCZeZ14C+8XePZACMxXVC
lPIkayq0DqX2lMBXh8xX7tZXeOguab5OrFlGY3qfUfkyU/PSrJwE9l6c26uc4yV5BIEN3U+7ko6L
irwq4x0eE9Y7g7eRpurclLRWFCArnalOmODDEaXH157tEL+nTALZr7abNn1u8F2fcGWiq5mp2VRF
oJMargLrxSx5u4Oq0nkt0xsWeRLLDJi2sQn0ryC78W2xR9Zr9do1cuinecCUQ52NWjKuFcmf/ccJ
sXM6u0ou1Zkcv32m0CLh1xap6uKLoiWIa8UNcT3/JaDIMh+HdcN1QUY0mHQHMxA3ij3TVaHau+yZ
ttPQ7M9H1LwpgW10Ga74kpJEJodJoD/R/79HFAf50w3fTQPCs8Xhvhdy+yF4eo7WbaKXktBrqfz/
eIwd+8aLfIZUu2b7w1CI8pSQrQlvCoUCzXUi3KHhp2FAr8msF9Bo0CWfIKPuJYAOJ1fWLu6olvNJ
3atgdkJdQETab9j+Qh0ogbD4NAT5RbJW/ge4KhSx70jnO3inHPhOTO0p3AkYhCSMeewHWDYAh31j
7Y+GdVer7RODKFMJtzOlOyoKVFbhsrjy7k9AlQFytooWPYn+Ebcn4Iv2Egw4BVMTEZDP5/oueyA5
8Gy9bS5Y8eB8mLgofUPUqepJEbDeK4komvPZyDm5mmTXm4V4N+kCRU2hO0gVGn6BlbQy4NioXG91
qENLawvH47nI+PE+Dx2ygv67mC5DUvo9QMtfRhBj1ywoKScv/MjyHltIRaUxLsHl3cWvGPMzUGSh
Nae3OOWXRxbd5SEJry7iuPWMskToQAXMQD7jSxWXVrdJE2/k2clm3GJbRkgllf5J+OYvyskNfsdj
GIErYhSC6f9Zskmd3MHFeWLsVfGqL3n8xY60SyRnPx1e9mwCnnOQ9/VooOaxeLwEyyH6lnJT6s0j
+MaGv/KvDmmpSzGszq4d28474kCJH/S9n04IxkB1+9ZX6osAr7L3rL40ZPdUoG8LWWgE73bOBQhr
rh85BSGW2/qPi0FmLDAR+dP3gr8F5uuwr1A5tRRXeTbxY3ylHiHUaWmdpykd/ri8QdmKud3cTpxS
BcsjR3WPX+lcTAozDi3W+n282Ts+4bFqgUCnINvWd+olCFROCN4Tl/As38vjWKqyPYIcLWqqvBF1
b7FxR6lE5XtUe7aCv2a4W5zwQQrdciX/8unvbxMVmM+iJ/dKjDaUpGFW/ZwXKubFAjn7L0eBawrD
2ulVSFQ2AAr+yZVYIUgGKO4dqeQaMx5WJVGKy5ayR6CSjVBfhAleE9e4b7tpxhr0Hjys/TAFx10G
m6tqTlSHvw1WHf607hLWvJHI/oY7mbkGjDRsBDYlyy/U0kMPyVXC0SpvFB4I8K9STxW/OWe0sVYk
kY6oOxopujhGG9YQTlEAeW296sVDJj69pW1Ari4QC10YE0vkaNS3mdu8uQZNygM26FbMWUy6V520
zZAoQX7eMF6ZQP1F3bcBmVUTS/HNzCu7SrhPMpF+52J2RLC6QT0ERZxN15P/++95LHVQHtANUSXt
LydSvDVcf9GA4lwz09gQXx6pK9KHa5Dcdt6Br8hLsqZK/54ljAcGjMmKZw+c/3kuy5sQ359+iBjt
rjwuE6zWJ8Bls8+K/NohwxjkEePR8kugV/65vLl+VuCg4Q5WuCM0gL6k3qv+AvQ7lWk9/DVQ4ffD
u6OqB1skMsOWisRBCKu7G9s7yM+iiJpTji3rv9/PAijP3mpYjU8dBEmGAOq27f3ZnXIQXgtoPkFN
CWACiQMcc7peLavQr6vqTeOvrPu8R8u9jcLgW9a4rv9S+EkS0boPXO3l8GAUBjNTVSIeISYcu3SE
zE/y5i/gbdhk2IB8D1NNLK/8XvcMBLxQbCmbaIC/HdV5pYMsHnbyF2hbXCet7uuX4oXAgONAaJQZ
2pJlsFyRTNPih+dsIYlKUcUnIn0VDRTq0tz+tiaTRksd3uZEMprbRI4cEckUnEL184ArYiNwpmXK
jaYdnM1lIxUe3U/rJws83/biHAuf9ftANTEGhPc9z13hLx5rfdfmMu/xtv2+wMk8ItCZ2ZWozQDx
kVdpNbJfLZENuW+Vx46E6q9aCUPtyhI/Oiyhi1oRBaywqIuOi6srH6a6gF9YVib2Q6fEPBJIYT5E
1XVyeFVi4QWIP4M4/gLritiUZj/JXcTiSq3P0k8NKY0Xxld9mHkCnJjrsr3TEiiyKxrwjYHkPCYC
9sPNBYUx2WvBKMaCODXZlkFNwOEK3BobbEgldbydBoJ3ZKxsThquSe+/SBOEMvTgHc9h8fX5tjD9
wzDtSIGlS6u/SqKMiJ4+ykPaCYFSLY/fx3GqXsGptmWG7xYYiqDIgOqIbU97Nf3+0ucb7jhLFdAA
v39SLhRzDiMyAo7jF/Wvm/zOyZUOGDdKetX9uZ0xh/f9XUEzpn7nHUZkppmpOacISRo7UJDOyBfX
bG3GTDJbNnGscyKGgKC6Ux5uTus8X01CPt45xrzAXJ4u0BXJ7960SFie266BDy3zGYdBVkCqvSF1
L29qBGc0qRDzSP6YAuLGcYuxPhowUNYmBqY9qYOpIojPI0XcjyFcmXKKieV3GbmOLkIb33/V1Hg3
AqToh+wiJyPegFS1yR75n7IUw0dkPAAGlcPOnvR+WZdVbwIVTlEwE6XN/OpXU7ZxJH9SJar6BLtg
I2GDhNONMBJAoLTr79h4wySexYdeoOmReHVxf7UTSQgKTXB8NyFG0Rb2Io6BjWIPvfIE62K5dEIB
HLo5x8WV4CbQGSkLSMS5YNVux8+SX6RH9UCo6SoOUBbak1augcl4HKim66SBFf5eqXEri3mL0dvQ
v09rzd+5rZy0b68N2EYq8mW7ZkMKv8UlaNo2A7RUCjfO9XNwSOYTSxhQQBt/itdI6/fVn2yeQ6p7
BGdkj3u+SAZiYWQUCb8npDakjvgEQj6ixZJQsqm0Drd4agGNGdtV3anFme2BgPFEi3TsUllCsll6
i/edYNMZiVJ3uD+3Jzknpa70yMfbo1C1B/Htd8WHo+OkSY3YDizKAOb4QphUWun4IMuhL07Jt5Ky
sfOu2XZV8F7tkhSL/3z6Qm5WKlGyFPut4ZJwH87ZGJ9zGvu3Qobr39MFqp0ba7Z01toyLPOCIf1z
3hvv5MDKxTmCUx3prF+Hj1I97gGMtKzrNpTlOSRI1dpncajmtGFiL3gOSvU1vQar3C9RNg/tfq/w
QkhCwHlMsWxY8uM4mOIaM1iYTKRnh7ZlCosREmxuskbI0c0cjZkzZEIZ61vBVJ/eClYDO+bqLhPq
SI7yp7fJKWTbOR9WpL615P0ZZxvgSuRcwwkICqbiBGgerBrvFbMEoWT0ptsNTLjXJq8Qcq2Ps8S9
KhRlt9+IDbAyTi6cIEfXgeQX0cv/sSEoXKKyHKhpL93Q8aYGRYgqAvG2/JaY/n3NXU+VoyRzmJXZ
Zb3+ImY+1daZ23JE5MTy/12qch7uoDhbv8THzMoVhhV5Ff8l1sbZHbHTmnxkJnRXYK/Dr16uNaxq
n9kl/1Ahm2lLauuuZ5ac2CwPSiXO8ZSYxp0QNvP5wPpH9tY0Dt/0RjDIq56cf1MQddVMIqwP7JzR
khC5uEMYwbCpspQx0AMgZT276YpGmZegb4hfTib954kt9/34HOhkwEju9KxwNACSaKWn+RiV5rFG
GgETEVIyusvDE7m+5Jv+MrF9+moupq2Kz+TK5wMTkAHl/roZgQkguq7O4im/NT44p7xfHpfZAlYL
y95xKE72tt23IqRii5kDUoEmJE+waDbQxLnpDKKZeiNJKkJQj3aCRWKaOjaDYdHpExkwUTBTBmGR
vYDmilZeIWLXQo5i/cRTFUAi3pRAw2+wn5DD4cuePUaWrxNNQbSOT3JW3YBr7oXf8FP393kEPBAH
LLDLWx29U7v2/N6R5yvHqrnBugvHTYOYPTlyz0Yw1gj0zL50MwyFOXJqofNV3W/ryNwm5oMmzrB/
5oMopuiaiq8vHyJUm5APijIdQeiU9k/FLGUoNQcwomuMaOrGH/0HjjoEReXf3IHiCfnzSCtT/nzc
DzsrqdKz0KFnwgYsQ5HGXSYV7+StonUzwuGqsQGRyfdmwsmSoWb905iARPOvt3/xt4AIOPkcJhB7
9XtvVm/NlE450K8sBfRCAdpKgD+IADqmj2OQvUOul0uEpHy2EfyCp9lmhfRcvYDCV3cJjL5kjlom
BNt7E+hKlFDlgGI/gascZB9wRHBVxJ9x+MiXjzG1ooJFkbqcTbV1p9S0jVDDAFqKf9Co/wo6s78w
+Z0FGZrUVxYMX9x/kBEqwTZkXXey+Hw+kFjaMFs87+nNIkcZ47zRqJV2jCP5ackI8MwZmQ/mPLW8
HP9p9ZuOPZRrpNz2vJYpcaQVn8snsPBgz82He37Yci/b7snERy9/vYKw7wm1SweA0qgiab5URw+x
OIt/YOPCjD5XA3yOBGli8JXGDdvmSmGbitjS0EnJKup6NRIJ/Z56d27Mvj0gLRTXVRMMpABgogGL
LGJVdapXQXPtPU1BFhiJxrIXUvaNS2qEGVYWuW8yIg55F6IKKL9d3ESUIjz1W1/tcdhvYbozaiBy
4d+bVCMEszI/4sIDp6NqZPzN3HJSUE9lbXnwWXCPC2bXnydVtWMUx4vpoaoWbA7/c0n9o32ByFzy
z/oTqVxgFcQ3a/gr5Hg9e5J0X53dCJebqBsQ/GYpql0fs3zTtE03mVMaQV9H/P7S4TogiHKHlnSF
OT951BdolRf/8Tz6cMNR5Q0H2PdC6eRCJXZCGDay7QaitLoc1Sp6EMAunsJkGLVRsAW2M+jJZERz
vnwFH5wZnYZ28eFm8QBj/jccCif06dC2Tfjo9mdSvsWIVlXco0QO2LbODLLliuniQbLwxDqLQuGW
QBa/0UKWeMNWLUNtooACvrA0gJkqrlZ7TGzd5Zs9b1nTjK1ljg1icHGswkJCPUJxHbKF+Nft5QBi
RnAOmpSRyIwWxsNcKny0KmGcxCKM5zQjZmyO4ppzX43KrK1g1ZOIT9Rw1YOUjzbbdLKkKChmgjz6
4cPg8FKV3SsBZpXOoJU6lpAdwNlAVcbQyyE81e+e8PvIvIFaOOazbJ0Dsw/UAwzqbEDrcAjAwCq8
kNnSUE9SGHM2OHFsu5ZU+w0QsqSKs2YHGvgk6H2j3poBAfwqAY62KE8ebaj60fDIrmrOHiVZe85J
54g8GFtSM5iKyRMNA7tP3LfPJszkYtCDqGx52bZq3f2fzKiA2rbA/tfghqG+e62kFWYmD3Eqg1tw
iKibOI3+o0M3t3w6SOipm81JJV6S55c8urGs6MXL3Sl2Xs+nFQGkjrcMQlYNkJJbwIqQ4Wi1rdIw
Fk2UfVtOofhN11rFw4bZOYd3DEAypga1SgiCBMji+hv0K/v3K9+N2FH9GI4KCakTqmNVqKewPYEg
UciSXrf2PK9s7cvW+St95gbYN3AZZUV4DaSdiNU1fBi8mWDnbuWyMcsirvn7zXD6Gw36ICHrohQ0
2Ll7pSa2L/QNWBgS2K/UBza+Nv02WBRnw6GL5dIGyJaLWha2Me8sv9owmUTcDVgcvcSljzuAQ/5c
O206NXnThD9nrwfoN8RHv4g5jEDM/O6MQV05GMl1bYhyb5BdL369D6tWFVKuLQcvxoJUZhshpn7K
J79tOxkYJ20ePJ7HeTnY6ZHLym3/RkNNGxkIrg1qYEQwPqR6ptXgErG5bJ/oegECaudeTmwMRrop
HMbu12TEPEMyORxWFkYt/WLDrVn/ApAmk3cFEJcePcKeW7dBL8euWTJy+Q6HDDF7MVNMJ7E91PQb
kkw5z/u3BthDB5JGsJ2gjptDLP6Ur2Z0CDngk/mIJgn9tuYarVY7rSz+98ZJYHrYGSo2jTw/vqP8
29wdLCr9rY51OG29w6s8MrLtvQnkAUONjjacqRHZQlUU7HIUebFc49cBC4J0D6gg23W3OEW/phsm
jBybRRsT0ZQ+tPDLk/vd+UQWuRJy/Byn3Xxh11YimtSx1tbD1wbk26ar1Es2dgKJ/ga9bJCsblWI
lJkk2V5yQPckNfVQzPgA3McpAryT97GjfwQ9KUScBAdkuNX1kmIFC+f+NczEutU7Ihb0F1AHcCiO
EkXS2rc5nKis0EbqiVPrbdnUAw/aDxwi5bboKN5OTmjLlczPLHH5vvF1rLNcqaXDuwP8EBQZhXkh
4c5Jqyw0lLICc5cgGIWQllLlgWINmD1hvnSS7bgVCwBBptNdK7HjyEXTiwmKdAna7NqoCPeedkkZ
/zZsDBtO0x+mcEJeLedOwXcq3fdRzc7BI+Diq7+VyhbQkuAFdWbcpXVPnEz7VAGcjVzWXNPUZqlE
bTTMzzYhgvNlmElFv4mb4TFbo6mx5twcQnYv43z6ojRs16ovNvncvf2FFI95dxedbEppg1h6oIT3
zSuUqN6zrlnNEZ14qrjm6kA6whPpvAvgh22GaJxXltWlDy5ZfLYmV6mur6p57KQG46mpUO1V0uEd
H+GFEu3qIhGhIPIQVB+53xwPJwLbEbNADSRsCCch+UgKdIDHAYzOL9gfZW8O24XP+NZX4Xn7kZa2
1PfLsqXxYWuRTZb2DTneEzK3xqPG8oU4BUMWHNLE7kkUaBL2pLCH163Ooa7zRNJsrjGsZbJZWxXn
p2Zt1Jw2PK0AWXK2QvyMJmqW2tVOiNNsbKrgZUTqctjaB624Xr86vzl0vqAAm/Wf6jAHC0nBI6Uz
hvs6K69FM+YBezzaxR6uQ0VCdgnsdYVYg3Z14/84mXLHSVhlPPzi9XONPKvrTHfhCi4QLaiQ3OIs
/41eEXw0U6xnZFvNMLYpZ7lleo44Z53QPl9wmIprNzUdXRBPvwSS4g6PMwU+7NyFoSrSlKQQmK5r
Vq915slquzfHtyp908INTdPE1msxUBP/cLrZcZDj93II/37M5/PWeY2hK6juE6LmBB/TyLoNRtVD
Mog/gdmOA8ab9XIEYNrEikjo66TjpsXsMUgeIxiBbey43J2UJyIh4gqBG35qjmzwF4VZqTicwH1F
1VNnjfNO6PMRO2tEk1i/Mbo8H30g8pSi0hzmgAXH+Br1WW4IcigFsfx3i8bES8GMuomk3BTtTzKx
M7cjpXH0ZzRdsdGP7YToX5JPCtF8DHA9G+6rYViJ8ED3YO1IFvmh3857O7A9l14JruCt/Cg12qUi
12glFtPMAkValtJKc2XjzVmmGi1IY2w0pa7yNpLG7WiFUvK32/9VJ9Ba0vwprHHNmA8Uj80K7QtM
qLUndANUsp04cqDoLHh68n1ZomCGNbcCehjk7Mk50IbHyGuajyUc1H/JAPKfLmrUcR0GGx540GLb
TOrKK/WPk2WytXx06c/7QZBHyQ8LjwiuhSDo+HLS5YnKFuOVurnpjoricR1QzsgeXNBUOjhLeAw8
p1/aynxqe2nPDTde4N1RG7fzt/SrTj9OLZUNxIvXIl92WUYJ1DqLzOWySvMdJqaYdS/PG/y7bZFF
7afnn/w5ops58/CrOT659MRhYSiUM8FrEzR/Z+90LpM1WUBJaqNILDzHjS+2dTZLTCz4+clJPjkZ
SIJcV3wa0UtcSPI+ZxmXeGOS2lPGc+EK6scrQuwpAnlzHvymuDufbE11McCvU8EFLBUHzq9K014p
oky4ip9aJ6INecRreOSeiT6ZS7Gn0syDvIxcdqSFGQbiBxUEQoYe05VwlvmNqNOWQHof3kn48GCx
20jIXsZN/N0uy+WbDLQIRdYFlRHDbkCQZ+eXf9LFaQg7gO+FT52gEIOq+qHRKzSTyCrD/Nz5UgLL
SSHVdvhCBXwm9lyeB3MKdYmdpX5rBj+I+R+hMe9cgkIOK9oI2wxUSA1lqCKF6lHO6rtHbFWmVlCh
sbw27iE2i+tKEHdoIQCNUO3LeHw8Gp87BuOnohcgWUlozP0M7eRPTHkzXy2BI1SS+vTK2uMDFVsB
myjfFoYY9Uz7BgOZLqs5VcxZ/g76aXzQJVJGQ6TU4LIbv1n9QmyuKLyI2Inh10fvWgNy0B8NgaMV
7kK8T9lbgy7t73qYbNf90y55CC7pjMx+wJESnQ1TYuIlgdXCeDWM1hUe7QO12mI5G4vBlJdRmPo3
+JHYMBO+z24zY81Fil+NiOZSTlYeziWdB1YDS6rPvtmCSswE/7mn5GgLzV5OPoqUFG230MLKss+i
4CAlF334b4ZPH2/+wRW050EgYic877qsbSpPhHlimkXXj5r2HHZhO9y8fLKm5LhICap8aVQhf5vP
ibEN293YFcw29l/gwK8auUcmYDQMeTAv48cx1DAE+CQG/kQMfeV92kxOt8TX+ZAg0WJZRKOJKB2F
73BmlKd8l+8U9VKjZ6+gzkPPl7nsCEmPHaw9bNPSZCPw2nNvPAnfIoqzyHlLVnc87emNufw4mE8+
SBpIYUNiEdwBdfsWPBulOFXfoFnimhbehlQLtijHuJI5jSpLpt9veYIuixYw2HEBecf7aMnA9e9B
rN9Btsxz2t86Boj1ZSFWg4qVwPh2LGmfeHfmZKmRqoEWyBFHxQgHB3X986WMDFm5Lo99Sq90E+pj
tAUWaCddtBDPNqVNSWDLdsUifZofrYkDQn+4ExfNmIvvTpx8+Khgfj9141/mwmUjs5x07ncoL5rJ
zSD8wA6OKGwPKj4OgC8YN6PXWt4mP4RxMYcxMv90rZoeVBdPhc3ghTQ+JAdrthuiTq+6C+i3uwQq
yEeLMsfw1DSwZV+ITaFv2rdgWtj/giP60VKebBMQWnElA7ZzNDIOPE6rUSd65gLTxjSz4ivSZMbi
jp1hQW7/832nKxZDz6qZxzmDpVTlhzOtz9Iz6H3kij6y5NYgjN9EFuJ3NOU00AtTrWHbzv7Bq0yU
ps9oRktGpPyMMVl6yJ2ws4L93uKzE3Q2sVYvkpzp77hjZrxqyaQK++Onpeia9ESsYOOYRkA/rRqH
duZu7coMtYfPZj3gok1Nk0LgrZ3c4q1Sw/DoHTJnZ/S6WX/gB9ej86sMkYXNrrDt1LEqFEHdKaKl
ZlfIekyw3vB4nV7DpgAMXXvMe5Q9XKpW58pPkc1ZCxZ5s9vNRoI6q83dhfZQcunzIlzZQKv/k1Dn
Z6oRCbH45oEgE8fpr0xO8LiijbW2B38GX0rwAB55T64JbNjlpU6QkW48ac3wjXiHqGhk3IRO+Rpw
PJUw7f37bCqgRW0CfmIMrDuIAk1VsXvnGvHlcep5u+6An33UXLJSjjbSvqpLZkM0fj0M5fP12j2x
WWnYqXo8YGKphgod7Bwo96Q/CIoF/waDLmm2008WC0lVRCwiqfqJRzD3MIg+i6FK6sCyh1JgsjYW
fAKkt0HO2ee8GU8ft6s/eDtsq53hiLbWndc/xkLvZu4I6xv4QpkOGbpt5QR/Du4ww/WXSWzyndwx
wnqVgvpDKlLJUOfuqkJgrRJVz8OpnkUfFi8KbNilpe/bmk7B0MuTgvtuhAjQX67Qrb8ACNECryLS
BYMVNyFwjgZXMunCWEOErB78IcMKBSOP6BMVA9jdJ4hX+B6an1hdFx4fIGRwfW6D13XQsRll754G
yboWUBNLeHJuXuxHA1abVFs5B2y1CPV/Zf8HwHAU1avm+KRAA+BhpFhanx+SPdqyspt5YQO5anEy
/b7dOtlgKN03w3f0uitnj/ncc2f5s5Wq6nl4Y0HKtlZ8tPjKFF38sLdtejYFBBpqhTPksdddHOnz
vh9R9Jn6NwWOQCy20lKXjLY04CnJFv66UAsJLQoXajvEwlR7TQs6p97RvPNwKRtnYDonKRxYJoao
SmXtnDSgNeux0oAmpdUZ0RuLKzMIFz312COrk8qXL+odveq3wnci2KzH5xhH6qS6yKsKiDqCgQEi
wO+n04jEDz2LK6VuFGWu/rZI6CclycXQuoaJ1Aej6b58k8QNijpVvKblWCBJ4XLBHumQMQGkGita
E2J0krsfU/a6zPVg2dzXFruk40n3Bmey2OwFT/9od3w+lXKKT3K41j9bxZ63xMHazHubGqMGxLkO
uFZ/x2n0ECXYVlz1rppxDFIOUTbBNkrZ3aC9QUOVKVKRiYxAyZUqVkOjZXNTeNWAOpBuWyA/ZwjO
CO15NE/Mno63zd97x6UnocCD5Tisg/03KpzaPItHvx75QQFQBpEZAa9so+FJv8Ouj+YnTVZ8rzJk
pXzlA1AGr4lxCGBMHzApB2X2stpekt83o++eAmqC6hxcRVFFgOsvm1J4XNi8BeRcg80RqffyW2Q8
ua2jmKv0n6B+ItDeRKR8ytEdSKijiffohYU5W331QOXvikUHL76RqdzpaFV6uo8XFXI8EY1QrXDU
i0r+jSeQ3Cogfbr3zXc1tXP6CIIfZz4oGcn2tHQ2IrZnOZc0cUdonluzdJdSTQAFsIL+fCHFeyqU
X0272i5U0nZ6027xFuSZTArz9/knL3AxgwtedKXE7l2OFf5hf4x9Bv8P5CwLktjyqwvOG5IenooM
iGYrALUv3UdmNqLnhqaOh5AmISzLXoFAnllFzj4f8TsjlG4Q3H+put6gSqnZbaOPrgInzk3htm7U
9BdZSQyB1vuc/XF3U+5U60iavcUTKwSoM4X5m37qvyn86T1c6Y6njA3SJWnnzsHX/lGunzEJXz15
yDD+d/Q25/gjDmxjNKLMsboVKucUoIgqB4qVcKF5SZTIaYgmxFx4mhwLAb3NEd7ln32OmDDixcoc
zBHGYj6/cCMt1vSec9a66FZdgs9W57EGDEMJ40b/UR9jJex+1XYsbcz15iFf3QTXbz0lQ6Qxv1G7
Zj3DDOadc8CGopd3+bFy/UGB6DVrZPbLPw+VK48U3brn9vxATM0jNVDDdQTQWLLNKSgEMPzLlgiU
gJbCgflyfmR52HpIfchpk1UvDdDO9k1ZcdotxRsV5pO1YHbsdh8fn01V9AcGY0opPovM/UR8Gd8G
uu865WGg5/lIDZJ84CKq8VtDDt4yQeEflb5+zO3oWN+UCenA90g+1zgO24U1cYiU3eWpx33WmY5P
DGaVg+b5UFBKKx9IKVouvA9TcxZmFRGNFb0kf8IMKTcUW/2sBrqEiAE71yHXiyPswJD1F29iieYy
MyhYzM0ZONeV3WYF/Ve8G2skkfyKKcSQUkQy2D1KJbB6wnc3OnE68hMMcjfuZ7gQw2rLit/P3Xbl
Wy0z+IHPS2KrJJpB2YaODV82I9Pr4568fxAypMrBF4rv/DrxW0+johw0MZg8bK62Xa8LDiG6H21B
su2s/98G4DWzglvstovjEapHWWyv4NgxThoQDYAgXurFmxu5FCuJ9MSm8XxmG+xlEXA6eNnzdhXJ
nY7IYdYYxKB0fym00UG7y6mOOgTZJBx7695ApROX1JCXUhml1QJ4n09RhFV9lEhOXcsSGbVWD3D8
wzemUA5A8P269dY0G+pR3soOPjG+CLogSYrq1eNSqLr8cUbTy9llh7EwKLP37YaS3uxaJoUB2Yuq
R5TZckIMKR1SSyae9MU29DR/wVl6L07Ku/explv9+L+sYdNL0vXOENg+irua3YcpKUC1UlxS/PMS
HWpPW3PZ+nXzcO4HwrN3PzFjuR7BVjeJ8kaVHuIEQsrzzimvcS2DEtIXRNy/RdZtdSFTfFK/Sx6x
SppIPUa+n47W09OR4PWMAR58HHd/pTHnYcG2J33e52wJqMuYYDjDCzS9GTFdG7rFoUh3EMOsqHjW
ou3ag+WmjjK63Q0KInW83zdqmaCoHnsMla7AJPwRYblxBeqC2r+0GHd3G9/Let3je5vm/y2evt0N
uRecCPdUZN7e+mQECWyCHTjFiPXi2SEpCAN0cBjp/ReRO6QMqWAdrBw5746lbdcDCHWqvgBWRDEb
XZIxe4p1k3qU5Q+FHWan+fF/EraktyfxW6RnDF/A64B3Z3VsPD5/UQrKWw+e5jtjR2oRkR73dJfZ
TJj8Zdm0/vFiu7vJnMW45cc/0XH3X0T49nKvgT0nHc0XaNKTw0waHZadFHn0PGiBKYtKsxM9zzL+
BnP5+y3f/8K8oxoyw+sEXhJCNaNRdZdO4Pz4SMjf3GR/NDxWBZfSDUHgWGq3E4Vx6458sxvOgJoX
KXLtSypCeHUYVznIZ6u/tMZxgVhqzJ7z3fdpzR1oWiZS0itQOAt2TgI91S7aJSoYc/WwG3ldIK/A
BphIldgl01Fl2bz/bJoqNxTjT8hSGG8LkbhQcNILS5F6KFSxgJYSGihvaaysE5QWE0uSNcf76/kD
fjSzJUKHRCjpJlHfqOGhm7scycTycB7+jH5Z8iJgCNC21YUytfyv7eMNAYkbZ6YF2iQEyQZZ02mL
Ln2eGSOutNWy4GNGW5MSuEvQBsjEr0ZnvweCC4Q/MsTLm/vPigCADpi17ja0Td6hAgfto6C49vaE
v22lE9MYr1wCRPLf9QqEn67veJGYjJxH/d3fJiTKXgujOLhbpy0YwY3EYWclSDTtb7cl8N448bsB
EjBC7qrK/m2YEF+oqD18wOPcDWTrL8Mt7wStDhOsXYyir+fubSVk04YScvPqjT1Gm+wfoveKVjrn
RHWY8cgCHsCRspXrftSEInprg9KbFMb0DdBsmJjfZY8HrK6nStK8HCHT7ry/ig8CVcXjfEA3H9Rm
7v0GW2VGRVSytNQGtRBdJA/Q0uaEz8h5Dde4tLGl8X2n1RqNOYmAgDzx/4czXjSLLbKG96QjalSk
bElDGAf/SY11MDSDogFs+Bx24iI4ChMi5k4MBViwUPXtS7QxoHhBrOgLStmfvyBcOQXHlFLJccH4
qm8K6iQgHsfRRHaClb/V3ixgSjlH0QXegGeuh0YZBEGUDqDRN9oTVKdAbwJUIfp4iF04xk5bHA5m
sdgTn6Som0gvMXJt/b2a264kZWXU9JUZ7G//PNwntSrj9U2TqUb/2YLNVxsMQy+vVzlAZYCAvr2/
HzPrPFle3EDxbKHcbqgJ//2c+58mRKtwJ/KKMIHRI/D+eBNGI1VYIEKUDeGU2W97F2MjFPtSZZ/H
XXV7Ry0+GH43DyV5QdrV96upwUNUTNgF3yxCYs8lu1JD+POzYxviDVHgdF2POtwIdb1ZltKdJEJG
EO1VGZ+Fa/HNHnLBTemwMWSR03HLKUWzWm2Gdn3e+BQTcmBBYmNarzfZacGH2PWHAGIgXnGGp2hH
9UqotMAQqs1ELw+P+imN2Ruez5d3uGTJ8g4/+2iLbJj/uLWOVnk/7jgAX/byaVAJWgHbYs+WNWw5
0C3tW9SgJ/wZb6dlQkqF1XX0SJxjdBw2G5U1IL5ywGr4fYioF7U6estXGVAe7qHsYGJayZFurVqQ
IpqHTHVltbM15SlOYEe/RxDuUc33nFwCvZkoYox7tE96DZ86xPlyn5OCndrpFPo86p4FzpqGghVX
qJHd3H/w6lTU9kMgUOvpW+JOVTSpEj9Lc1PhcvacOZ9kDpJRTAG72fNQYqWDq7BHlrUpRic75Qlv
53QrgSlkgCbtLLSpHZCVE1uPeP003UDpluYjswls+7/BdUcEbqa3fblaq3bdP1fZc1GQWfuc5XnQ
IV2IvPtwrVNPldttS3z/gHsijVbMzd0ZzyaYNLNRpiZreTFXhuUb4A3ys7p0RoNcx9+wPwXlNBvF
Ita6zsJKFxVG71ZQEVTFJdkYWwe1t/EncnDPyCtmPrtKdXsZd1yTf7oTRz3CWBXlB81Vgn6qhNH7
NTWkQomVsd6668+F9t9bWQUEsW2FTzsUT+MNJlA5Rag7+HIq5zBodjwxCYLOAPF0Ifhh5sNFr8xS
Fa5IsqW8N8R4lbsZ90nNfLYt65aabXuHBTfH2y63YUzmzHZaeY6YGJ3cytk8NMkcrw8bqkkm+7WW
geWx9Oqmov0Q4RuBLLnRkTGCQ1wO+2aabRHjwr8DHfwVYzCO7o6DtnIqo0wEJzNlsu4Lcl1pJlMh
U6BtWqsCbQ8i4hygUAAv6Wrq/D5s3+tYlNSHcDqVUbPU/NEAE9s5PFqI7XzBLnGGB4qqVNsmRhC1
m3zsiWh7z3Rx/E/kRAG658bSyjqPaEDEgAVXxJV0BSLAjrdhFzUQ4Y5/yp1vtN3XDVIPc9zRn+S7
1OofhUziQxFKjsCybAw9t0ADP/bMwRoejqdCOZwagNSVcpbLL3LK0FUR0VI/DcekVNG9y4NHXz/m
baGS/pr82OI0XfTidoD/CGgFpLE3CqvvMhy5QKYLo8SQz1IfL/Ik/NZL3dYC4vY9d6uoAJMWUIlI
iO51DVCKYvGlSYMAkMslnhGSkO/cGEdUR31zlUZFIGDG7i5AzYZ1DAlC/k+KqTBYgDptmnkAEC1z
t0aI3F2ZnX9cmdXNwVW6rk/PSzJte5yyovhy3jjGDof/pkWNkcOFWhiPuxqKJN6v+hobyYvbSKdT
QGq6c2W1x0fi7t5qMxqjACbHM6ljkbVM2vzPQwuBPjxghGMMq4BUePbgmUHpt7f93YFeXd+XSLUz
v8Ci5Ckc0WvHsJKug6iXLHI4bvF5BbPOw7WonOgore1XXa3CrYIux2/Fq+gVwTv5uL4EcBdzfWig
pp8AS6NWUrNbTq1QYqQ/0wxTdmVnHBS2x8fqokFXqUQ5w8exqO4Qt75I4XS9bTQmpb04hOn203ul
dsEhZZP96MW2hkAaA4qJb9LnhurAjn1DQ4IkbezOtmuO6SKIWfhC0kJoxe1W0XnKft+kdPAv1zOD
E3JHjSurnPz7ZXrC//uK2p6C3qcJ2G6FBF0ah5pYLfj2asBCa8MssCfv/SYHFWKCggh4jXwIp8d4
4nz4UCchl4ff+IOnbqxM62UXUiyml/sal1xkmXdfBc8FfTieFbibbhAge5uAkl4yjFQKbyccveXp
PE3sPnf3L+BayyCCS4mfZks50dWKY+PFgPywoJDPKOEIjRSgcrDu8YfY8PeAvMrDoIT4SjMM8Ufz
ov9o+qqV2uZzN/PF/31a4Z2THm6i8kv9loXdM0OrEXX5XaK5CuMeiOfg5msrTO7SvzHvZ59ZYXMd
PtulgceIyzba6sHRjX4Rg8XctK6p5lpQ/TCEJcLGYtDuKDj5dskIQn4gB0TPvAGr7LRFtjoUSk1N
5O2filUqr3JDzgTA4UMU9tImx3iiLZQVwZDh4TKYjvGchKL7Aa2aAm4LOjnEi6N8sphCDczJEfHi
HHxKHyDtF717d/n+9ytzA7yyEqG7/jzO949H3ZCaT8o3YxmR6T76EmmAXV3JFEZ6h9KcG1QCzk7+
xCBBR//F31P8pGVp5g6uUZHXdFjWs+s7DjRvs9iE1KMee/EPbq18AjhRk/KQvt/6GSVhf7JnMpiJ
3QsxnO1Hh7B0ezuv7Ns68iCk8z5cKUhQmgZhJSGG/pQdRPMFK6ZyGQrX5npSL2EhtpvGmPlnHM/U
Ns46ZOV7kxM8U7JM2pcN7b/XtI2Kcj/wHqvIgdy9PDOtctKzSp8jMo3M5Up/D81Cj3k0Dd0eVRfJ
1N/4Y4BtruH8Xb1XGdGyTcG/qtjFTgbrka9Z6OQOTy2wQGIlewTqsFcquB+iGGmErR9Lqbu9DuW4
/mBnD9nlGsVpVAAA0+hz5/IBWuY0p5Nqkk+vL7vWYNUPTREu78X55HhqwMdjn/7VRbW15/uIsZ/M
YQELz6QXwVDIKPotLkNLAfTxjUhb2Z7bendffdKbqxYeuwAWCBwxxlMY44iOPYtmJaBYp0PVwRo5
GE54Llv5p7mGpcHKPQTt3BD8e8qVu+dEBYVTIDldUOg8ITwZ92RXWzkXwpqdLE10JsZDQgNWODJ7
GjEO/+KNELy+WQ5EZsd04CLxWxwyYCpeLfgpINqrAcva9fRsM0cSfg2yZy5Yy2fwaCNzYPV3k5A8
r8bNP2eBbOo3yjPG6NkGjBvGGBqlNVzGUHjR2+U6W9jDcCKlpcLeB9JLMjtkyMC7dTR+FWWPJNI+
G+inMoDRguZwmHyhTt8MwZ+ST971lBkXBC1uQWfYb1Q4DvDRQ2IqesfAcZw5zpoN8gvbjDO3WMxC
spqLwOa12bVqbWyQoJry/jmZ/dogeiHUdI2ThTckX+qNhZyDeMd6M5OaFt7xdzJT9os5Gs8VlA6H
LW8G5DmXyxGTZTVNpGXUNlKYwhWl/cqDVKf+6fuf3aSiZNIM1MJ6SMHdL1CmVILnWQ+kTOJCGsw9
Lc4e2nu06EQsqDhoujuaat6DtQZfljF4RBLtL1VvNE8UBoSSJmC8huvvitGUWdLkbR7f3MVYBWYb
1EPe0cRxWmUKJSvNOy0U+jjAv4L3OHzG8Ivu8Of8gik4EYuAM2ufxTKaWPbx1LAk0tW4ARLbVyfC
DB+sL8T13Au3ZJEWhLPAJyjkH8bg57DiiHoQK2u6j7g6GuoMbBD7PW/w6dokaEv/9NiC9ycK5RJn
RTLG0+TZxAOgVQpMdIhi2wv+dk7EpF8vRjSKO128XDnzmm5sDkd1Mjffhcle2jgFe6l9WEJpPgII
GuX/Rt4NOBHCXujDQNKbA6G/CEvznIAiQeYykXcSZ1frgt0nzfIvPtN8UiKfOFILC6XYNdgk5eFm
22SOMKN0LACwVLavv7jWYUrn8Xp8PBTeHyeezHGfE1RhQE11NbUDnClZJuVH+biJhzwb+ZvqNi1a
0qrYWOzPYC0aAcxiDosUrfDhnDgKc8P217A3gfBOnzUL8hpFoA3FNJgZK76gkfq7PAZ+3WMlpKMh
3gHQ9Zjot3RTlFsdRUquGzXRHwP2B+I74sjMdL7J6bdoLx5dX+iSL/Ld9BAcJTuHBXYz/a8rPf0L
ZZO2bOAeEcvm8JQ9pU94cdAE7srGB0Xt3KRNpZ+4TAifEcfUkX4loUMqYqddSW31GP7YNU5GuD3u
bLlRBPH2tjh5afY2YB5hfjG0S8wQ0ehYuvV/WvR19CocFQD/uvB0PaG8v0V+ICQlx89HTwOxlF4O
quyU6mSHPZa+wJuapDCCO3BCldmH70C7bLfR8TmpsrT8O058p/Jp+z0B5hFYjk/iNSXdNd0nv1pR
vigyjhMqU4Y3sfnDlYdidobcKfWfDPLGNcApcKF1zPQGxt40r+ruoG38/op3yWWiOY5w3Iuhmt2h
uZ/cSrjNYb37ldxEccjxEMB3vZVspBfME7afzlcNyLNFxt4rnkYRoHu6POGqfHI4Qx884QmwvILz
JI7tBFrr4VoL3vKcOHRXduATlJTsqXobTpYgj9akocRzXWC/hS86W983b709ysytRwYanR3kPNs+
zvqU1oWG9A1tT7NFiB82mt32AN5mICtgu+R5axLEFLC6/DcV5dqpynk8csh1qo9FQ2iZShn6OItv
Jk67mBI/QcI+A/I0x+/iSy1ZTV16JL0ZYqXPK6ZIwxclF8BMpoF0XOYaq+rPwp6Af9aUipmbEa9x
7OyNiImFN0uD0o0BaqI2fKeUMt44GiisKr7GqvK+q1kCI2WpYo5W0SwjYL21kM1s26Q8tqIOh44L
wbZzkN3g4VzTqty4kKWlO4DIY/TFfb5nSsK00Fw0AJKehBKKUZDdrJurffeisuuqW0arn85Q5R41
F6+EZnPw3aB0npEpXY+JZ4DUA3HG7d6r02KR1iKan6Trct6NCF3EABrb8w189dWWH9hDvc5unzPE
vRGZ9SxSgHXYAvwcKR4gI4+Wy0kEuDNDE0ewzW/7dKVEAH3aUn4m3IAPmAlDpysx/ALYnCQZpKeD
0rUalAmHiP56OcGr1/cBCNZRqAPfFSdd68yl/YQ7Aj+xjESMR9gOGBmDl9nWjEPbuX+8bnEh1kh/
pfKBGRFncStPxxAuS3pf4GQIFFMkmCtdaPUVvRhscWGFic/maOY49NHVoNAKva6ULS6CX8Lgq8Ey
X0U/MzHOGd+qjzMJLzwfM+6+NjH3EQZP0OaS10TwdacYsTxKtbmSfNRSztg05xhC0szyHucMij7s
D5TLHggZ8SqC37OLQgTq3ro42VPtV1AmE0RQ+oDBUlIgHhU5fbUsxg2pToxvsDncsoE5MPbxaTOs
XE09j9+rGHCgFCAVzgDqU5/nDUAT4SlDoBMqmYxQA8rF9WXKFYW+H1S9MIv77sTH/uskOQIqExup
v1Q7FXOtT476dd7vLTyMKHgRV/BIfpmxn3arVQ3NhxT91sgcJMBN+hK1sJk0faKtQKpGPtYFunJq
KyewYrGA4x8hhB1nS+cPIMDwK3LFCc50KjwXY2k3jVi19QXTeHX/f3jla7+EsVOC5azsY2i7iczZ
NNIhIf6naTt3IqA8TwgIHNDuUpeOAPzwuedOS3T+rFGvIOk0l2/WKBpmJM2ljjN8/fkNcjkIV6K4
e563d2WfVqujOQNhxUnfAzF267ZbThE78dIYN2shF+cW9RM162gj42bUr8rmWDo3msxZDLLtv3Y8
bW6PLUnccJndU4spVlKdjl7Umste4Vd0Frisz/2y7gYlfIY1s394OL67L53llTLRLMP8vrUlOpsI
rOv/ZEfFBlXdv2K7r/QqBiohtjb2QsQY1bxHMCrPTFfaQBnM4I2/mk7MWoo1aHcADqXhCULHxBdp
QCRaMQuzOsrRUzYc90fJbh5UdAqwaWyKVPQVvwl2JaaGEowZEe5GSpyoTMRgZQjpta9TeHDMPm3Y
z1SW5Cd+pofuW/TIgC7ZdESpPPcq6V9Kj9N2eV86AqP3GPAF4RCQqiZ18mS8gFX/JAL8XbNM990X
vuQjcbi5F0k5tnocsb8r8SNnqs2xz6OblA0Pcsm0UXPsi4ZAyRzflalTL7TnA2uo9yYhahL2VuHB
vlQJ/LExPiO+WgrSQOphXEOE4nUNo9qQ/od9S5L/jVQGJV4jNx9bpwGc0I6vM2nSRF4Orb2J/X5Q
V5tcu7ck+zmeEN5fXpVduz2/pJdWif8iDB0wmhU1nkmfukxUr6mZraO3xyUeR0smYGZwIGyIjx8C
ec7AG3XGgEBCEJVYxMy1Odj2HKNUdbGaiz3qgvynC/dO28uM7zMO/u1LtYAariRolP1f/HxQ8LKt
Q6usb9RRdWqpjFr75AzQ0hxDsJczLVuQ7SgST5Rkj2qowd3k4bffoLBHiBEMzPdQFgQXWPj3f0LA
x6p6aJoRzgloLxG8v6YHtAfAfhp5GjwiEp6h4WCxpiFeM+fYqbRgMGHQGmZ9YgyuVPacV0924u7N
VuqOrACMIi8/cS21ghEvCoKGLqeWkBwdU6c62j0NgejP+q0iCEyn4bW2xtR63KibbCNdaz6MVsqC
PgdiKTm8V/h+7ATQ+RxpEBLOloD0t04SisiJS0FHHaGoXZRDck+VbdME7CsXVqZ2gFa4tlrPUuAt
fV9sGVuJLN1884hBeFlf4edV+HKL3/FjBOmyWKECqLhCk4Z9R+z82dcgMe77sq9o2BJcWY6oiU4P
/FroMDCglYnkXBYmoxG3B+schFSB4Itffk3gH9uWZCg/l/qvJReO+nFzTXWl7ceeDs2rOI49LdJL
3BuC9ZEWGZM3Y6CaolgYWfiND2roZytunBb1Pqm4kznIDmtLCZDp1MA4FQfJy1JeWgPntPhvg3eW
J1TmJcz52kRQQ5SLty8yEuq0xqFr18uoQXAHfkzfJDQslbL1jjgFKAVElyMzC3C6+fm1oJyZnrbc
UJ1vOySeRl3YhKimBRHXSaMFn8IRidQ2CtDrsAIpcMKY5ifnl3SWZM9MmGo5Yt22rIUExFQtIiDS
H59WW39Ast+4231gp7f4rPgyUDdIzp34UWWKhXJGzRXU/9BUI+tTqJ8a6XgEBsV33/XFtUcDE9Eh
1I914y3XpJgxuCtqM8/FP+J3dY089kWalIoHOUUmXMX2tSnE/bceGU+FSY/HZeDUCkjt4KeFrFJb
gB5vBsWSYmPpU1EzVU1VlXowlic6+oyJ50ALgOBf/1IOCAItfl+muxqaLPNhdz/kjrm4t13vI9FM
CDnWuM2kzWhEq+kE9mbOWRjblp149qwGExxFnj9Re55zesjnmcZ0L/WPjnEiJt8wJ3XkvdPRMBwP
Z2hf1NdWZHu0LqXutNsqn8fiadrzyTp4vijrMbUJiRXuEerwneGAGWqg7CoV5V+r9cvQxxudva6+
B1Cq1qN28wh1JpJzuIoeXyWlXMQ8f4h6Ezs4fNARkbgy2PVNyYtqpea1FB28niTXiP3Uhq5NQXOz
dIiN0203ZH+Fc5uec56nYL+dTg4PdMtcOCdcIivLB2adIbssgvudpxvyjzKWDjm5mMzjoN7GrySY
YFWbihC5RLppi7h9xp11r2TlGKx8QA7lR86qcjwT5hWIX7enULjZi95PYCVNyjl0eCZ55fJxGvRB
cRRHiZJNL/Rlbb1AZj5RCzZSFtbGsDwe/msIaokfM2L47q1mOKtylpmPBoe8weepNmIwLO1GzHfE
HDundgdSLrBg1AqcyAUhymcm9dVOQ/rscN7oWbEgUI+aeRIhuPbLYB3t/sUZXxVJHDeO1UapZq8U
AcdbhzjFkIdeQaxTmIXPQdpQRvUJkIFszSRd9CnStLWv/P2t5mHGVcLf62ivM3CzymeDd/FkqHsv
yIEEbpOM/5mhUBKxukcQrzIxVL+KTEB6VaVOo8dMUVXKGtyswOKd4ZBBnt4WkrOwB73K+bUB3jTu
4rRl6bASburzq3xvUU8gmdcE85y870F/IDXiRO5wB464CXkiuTnxH1c6nDzwN7u1mjzpZMi9qUcJ
Q1Aa/K3BAt277Z38ak+5wk+6Y1I7f5x2ny6TIHyBwhfEq0kYPmAGzi2HVFRGKFwZ+kyVnXjUKZjf
DRC7dbCdWo5L1d9Y7MO7B3FWQGUgnN1oSbmophQaxnt82RNR1wL4Ybpfau9dZqcsXhGRDapCPwdp
f+gzu0u0uzJFLnwacLix5AP0bjIkJ5s6GA5aXIF8WnWckReeKOtzp8FLpPpOXM5piUir46+/FQjz
Gn70ICcCFcnklKyt9+WHZzkzurw5V7B5nzLHK8/wI0SY+ZAwjvWRcGOO6kAQTTxckF015hWcnvjT
XuE+mYMDqr0Z+ig1WV7u6Mg8OtdpOdwd4oUbEuS6wbU9ZnuYb5TtMbBMPDCW6h0VHUS9MmSzSC5E
5tFh8mmk35gm3vxw5hh7QeDdK0AZVxp+HXyZzKslo23edECyJB59Pihb8QFRsZr/jCaUYOzj7k7G
u34xDBqD+zEo/iu1H9YBF308KWk/M5ltELSJQ/yFdbfJh5nzes6b7GHCibcQZaxHp2hMo5JsnxOh
u+R0AHMy5hF0yKDq3c8Z6BEY8sutL5e+prQoqzCB8Y6LHSmCeLDx9czvwc5mfTeavxlxfCo4PGL8
vmEgUqx8WNNHPEKkMpB5v5mWTC25cDFwLtflyXjQEUps9riFzTs4PaaqLAT6vfeU8aeKx3y635qS
7df4PHwK+cRgIsENAdMl1vz/HUiSov9BCB6gyEqCw66CTTnnzOaJBAJeUpAQiLfk2RxKnUPUJKCT
ag75dmbSVhAO0JctvDdu6cgb6LOlDjzUAtpqx5SC13GTtAKls5EQ7BSsceDsIBrMHXXU+4egg63y
tlUDWIg/GGdS2IwGcIU296oxYW0nK1nzidqf2RkQAlUJoNfB1DW+IGojVyq2I7mE8UfGTIYizQ1B
7DbvN09Y4WlusFwbk7efdIBm2mNlF3JQFXrCXysYqrp0DDmdAdOCYUbkp1NXOvk5rfsWXEsocn4o
BgLFe9k+reCG+8/ufj5LrbhVglAlC75ML0ymC6tIa89jVh2my71FC2izMEVGKWwgzAUE2HpWc/Nc
t0CppjJ1EMkBFRNx2XFAXGgjOgAO+z0ZT6c2Vkw7mk1yQkE4krg4eGI05YOUakdgLDhEr3QqowBp
UMljEpd14dghjXJ6sCVpzZlaBotKyBmqmlHHyFVYDEcXV4Q/JMiBD2uSdT7S/oaxSekiu7hf6mQ/
Ez7ULTg6+i58do9gv+XO6d9qe98mcOyBeCPcRCyG2kKOvPSosIJX+lzkWdcKtM3WyAZ6wJ6FTTGc
NsoKAJAc9gRSxUizmDEFfEeMKCjn/0z8B5Fgy2ZWnC8B7NcExwW0P6Wqk079ahIrIObWyg7QoVJa
EyppZQGIMvD+4WXoyX2TizOyNp2Hj/Gi4g2ED7S/ejY5R+YaUlwg/AL1ktITIF2xzV9cQU99o6yb
2jEnE0dh3LCd2OMRAuh1h/ulSudzMIKBDrk6pjC9yX3QPS1lnlVLyi38Y+7fgFy2vF4dKrvGEd9b
qxNONh5MtQKPnVYW0ZLvI0b+vhR48hbcUSjurXXnLD5q/f4g869r7ax+P9NDsrjokH+qLhiyok98
oMNbkP8hOEEbBlHam+mqs0lYteDjazVMzFTxedUlQZfMGUbjZHppKpBOhBU+A6GQU6c+gn9L44Xx
Jl2pVe+wDQD/7Nsog0CgKyidvRFShXL5rNBhg9NVSCvW0DlJ/oz2eZPhs9xNN4rNTGXagZChfjO9
nFWmIp6s0tApfuch/uTFiB2nQ9KiRjCzhSmeZXAPoZBordsCDg4VnL5u8lW0e15vLG+8oPCsmHzv
/MlGtLOmjzWNwpnuHYruAmNQQ8zw6txyfhpop5yijMPO5iU6nGmWzdSRlH0iRYx29O45cK5J04iD
9D6Jsm3o99zwog86epKZwSaST7p5BJCmrpIZRkzTD/smYw5yneypw6pnoPmPO3JyxVwCNyA4V2Rn
fk2036ckc0KGIqHhN/xruxK5m1yVjqD6sE5sSnLrrDa9AQEi6XgFh6SeOHM34cV3J03zQydPjQ87
JiT2wgDQ5Gl/xszy+Jj8rTqy7nqRyVyh/9mFJkiywoC1O3WsCK0IxXpl6EGpnULyfk8OUEUNQi7D
8QXNNMIjFJ6+wUlj+MsqfivSL6zBdxc8Tfxi+xEDBgB7HpUNh+AN+S2p+sVSHw3XRzE8i4IrQD/K
Bgxzx7phhzj4fEJUPZG8IRPW06iucaZAtkn05L61EFx0+1GDKekI7thJXTHy/ufKSTfA8aqPxUBm
m0q7Usxe9joRrNseQ4x19btpH82WtKM7v22GJyjVIpINhQqTpJPi9dpfibZEl39cLREZ/DwkzS/L
U23ISwBHf07bAnHttlPQyv4uozdK66XZKGqDCjkQSS5lic/CEmON9COLigeCPOvVsb6bNzr76R1h
AkjHAZyUGIhp54yH7uQiV+ZJGnSo77uk3S02KycAJ6U2c39i7d6HqVggUSYx3rsExlzJKB+dr35v
rmQy+Xoz5lOdoZGmGo3KiRySvcE9K1edr0hvrP7wEmr32FLTMd0fiMHrRXS4Xdh6hnPe2qF5vfVo
Umti/oD0ixCzym26ELtbtJsWWz8A9bbj+BjCQvMTdKTcKuwklWoMXPfNe7B4PDIsf9SylSGvJMKi
T0da09PHVChSNCNZO7CCsgWb3K6JGi2EMAgEwmVy/4g3/BwldEUi45fMUv4Tnjq5K/aYPOPFs8nn
Zp74fkzyE4q7PsBGnwacSBi61AlYb8Rvu1aqgUrNj7eALd8l46HHuD79kyRrGy2E8598DljGrk5G
LfzmczPaAW75MkEKQxVdy5ZRCzoIT1CxvfZcXwtBbw/j+3fc2E7wZBMLSwLZuCRG63YyKLwqE8sq
x3auwxPGlxoWyPtGyNcgN68T5Lw0pdj6joQd0VDX6LJ7du2t4zL6Yq6bUH6yYpWxLJsGEkyY/Msv
LKOx6vVcQ2ANyCdT9NtgSvR0cLt3fEzx6eTJltU4XpwckBiUqQq/XQnTeKAD7heONkzJr1f8r7ZF
EY5d6+dnG92F63yNzaEVeLJxrcnYXAIfSUsaT+3LczH3LrTIGj8MygbhhI9k78QE4/V5lFkVt2sI
Jo8S5HmefwBU3ghjDJE7quK5i9WRq9KrurrW0vqAs5u2GixoYfS8IhHRMDocP50MECjb/Nq/QdbT
gFJ7w727ccv6wgCbj2mYl0DHrgJmvftpSg+cg2+YZUiH8Q3PxHbrKs4HEpGzGf8f8msKOOxcpjxr
ESra2rGT5Wj6V3iKDmYqoxYpFcfKbJwAH82FumtwE9v0NhDmbdOuFfqSH8evigyErouUWoa1NWNH
jknWF8swpL0DVcX6ZRRRZ/xXHTJGxdk/Cw6eq1qUPWNCRpt4bZTwBqBc3oxNGg6jDwZQLnnZRYsw
BxXCgxOwAzyvMMC+NInHEBWORpTtLEfDSujVeYV2r0To01AfCqAiA0Yc2q+5cyLT5C6NW6FDiZlf
w7ppRY3ZS/BBVWnP9go9GTGGhginHdj8+KLYd+yXbtL94ssuTSkPSfsW5EGDu2JEuIEafsaOBiS1
j5/lOYoYWT0bobTZFfZeZ/d+XcwTJJAeJnh/QRXmpsWJ9gexGTgLctSKlxwhv6ZRPu2Yp9iW8YsN
NIW4NQTNcBBosLfcmXU+10eJisz9rTadcf+ouXyaCP0JUPpkHAjPFM3RAczMgka0yHWXMniftnqU
WsC+Hlw7MLar48P4KsSJujKOreSw9jsvTyuBfySbFqfjKpSxV8IjSiQW1AU+Attb3H/lMEqDQjUk
+JmhUAbNUES4s7uB7WxGCjR/OMFCDPrkkmjbcyd9k6bkLhjSji0arArCHJ/gGvz4PWUxBrIYxxF3
kSTCex2etwVjwutDRsmnLEqbP7WX7zXoyVhTHXnYXm89uIDGOv0QRlqobWNln5vymhEGfYiNGt+6
CoKOJSpDp8PG1786M6IfoLVd8H3THbPcuWAEKt93ejy/YPlzUslABIxQX1titabiKkPLomFBBsiV
c6qI4vxPQPfb6T3aDOm1575H+4t9bzUQcF5xVgggI3J+LAfrKN72dPBkFqWJ6j6Zipc66F6UqXcV
mAGaCc7vmGC3UKms2UmVhscHQBZcIt3ZcWXR47NyMiLLKWx3ys2s3PoJsztxwLR1RrSKUp3iRn83
tVgxAO6xY2qDVe+41A4ooz0ClaXhn0bVOHXFagkXVjIgvUx+NSKsUYFDdtuSFyvZtTpeb5ng2pyI
Aal32iZ7/W0b/mYbLVgwFqnfI8YHUyAOMzrVelsZS16wuVSPe3yecdtjQHEcUhs+91Dfcq352jr+
WTV6ckY0u8caXKZhOB0nj5+yKEZZI13vtlA9bM4wOBxyzSU+bHBLE3x/GhZC5XbiPQI1OCddtmw+
KSw5u4duh5yawx65WJ51RxFxK3QbQI2OFLgHzqhjfJD0foDjxLsgzf9n7Qeu/+PA8/FRtLbEFCbr
hXFNVcA+P90rdX2dEBoEEhedaJNCKu+IKCNhbOWT12FFfkbmhhry1JW1a2M0Pc02Yw/mZ/BAkl7y
qm7ZAwLMHfvCfxegQDuhDmD1KnR67fXXsQ5uVDrV0WyLbMU0IUIvCMxRHG0sHDaE5DiR7RzQYqF0
e3eWITWJS+xzQdlHGjus9ybG7mEGHAgGR+ZQF1GthC6ntUcmNKAcx0FVlemOOI9QVFY3VW7ZI2jk
mJPx7FDzhQ2ScuAbCo5sLIL0ZRVz6mSPXzufU1tqa32h23zNnVczKv+0kk/gZZLunB2ZHDQIokBO
149P+asJBpYwf3KxOaeIxDdB+f1e9nY/W1rVL1p9xh+/+9LMq1ilycLGBDP9wBp5H64QLeNALI0o
MzAj7Jbqij7R7KCW4+epQmxFu9hdk/BapIayNKS8EpJXh6gpIE1+X/A3Q7ykY1yeLY/2LzcknwvF
CCFSRrmErwcUcC5s/OfByyQh6IODvfGV4d/JMbZxxRc/rdJT8yZTsXgcFZMbVS+BfCu6GV2xgLt8
khyhf7Ml2+Aem8PilWXoX9b3+hQvvzZedW+7PeuwH8AJ+RJf2utNip/sK/zmYY+6T9bybRrH+qIl
p09HSEsvesSgCVs1ftaeAMZkYSGqPJbsuOcK9fNPtVnREeZAjcf/9v+u7eMbJXO1z6ZuRUZgvuuY
iBm0qR4iXdhMZHw8mj9ZAHpdESrYS5x/DNdkZnKx0pLdMK5X1KzT8NTpXav4CNVs682imS7l6v5u
UL5QxqbuOmOqyH6A8Xric9NKsLF8q1zMcH1uVupyKfycjrYv9qj5a7dllpVbrWIB92VpRJGAtNkN
gUuiXY+z5AiFbyK+F/Daon/k8UM0KFhv0KNgpLjQtF+zrv5BI3W45JyB884dr7IDk/HjzcNd2v9L
UJ+biJ1e84XAf8NTaQgdGVFIZj3xWEX8Zk5s2sxIdwqf5u97YRU8+SzS0y1rLuLNLWQbtr688+sp
LVi4aKhQGoxURjw7+logHc+umCCKoHZqGp0fQz8mwCZ4fq6n0iP9b9PePQuXmeQRKzjxfybZfNqD
y1DqLWiLsRCdULhe04v6BkJ5W8BI3V9xvlPOlOWuw09t5n0EzOw98X9XP1hLj473J8csrX/0v5r6
Xv1HqsRuz/I/cdhfQ2cdx682Nz2gCXtMsaFOsN3cEaTw9yCTaVNM63yg7Fe1qgjLcbjWUDg8TSEX
4I4Uei7aLNCCIE70VouwsbcOm89S/SQJHpipq9Rtd8a5hXBnfCSfWcWuIbwd688ZuWqen0iN1cO/
rcL4ijSGMCYQZExyp0GIkgybZLRxa2/yuaiuudHDBLCmk6HZ/Nq2Bw0hxyAV5NxDQiLpp4plP17Z
jE/8d+I51KCUYYUcxTFL+oBFXJsWDgyG/ZaKR0eVBeIiXuE6Wo5YS7Wzf+82F8FQlcNgJenk5XZK
JMY8cFPCL72m+6wPUz5ykF/WDG7KdJHIaC8hL32DotNRWSS6OTM6zmOiL3mUzIum7ZvowxR2ho9h
X+FzJN0/CohtxHR3ZTdZAi4npaNBQofR7n4hbRhmomFppaDIlxGC5O0Pg1eB64bpDj6HRFNjBlj1
WW5aAeLzggg2W4Qkv7oGQWlx02pRjZSqku4J9+22R2Cj2PKxuV181pEoPrMGse0G4hotkM0mcPvR
3E7vAU85RVwB8+2m+EEUe4VxyavIOxhDGe2J5QZ+sMLYFiVN5KZbAWri1m4QDtNZX7E2zQaPl2nc
5jk/7YDQVZTWAPy0MEBUiXVOkbIA6Yn6+ZdYfXftLozj6O/qXKwJCcoqeG+Y2ZGAtwxBpxUK1ESt
1mi1LeonOR1eJ1/hEAUrLW9GJv4ctHAhabOd/vgtBQtx/EGyKNNkRL53Sn10B/O9oXPF4wt3WX9b
TDLYgXqQitpw++ugdSBrM9gA+zY5tI0ZmXLgbxP6Hv146N8PxKVZbWtq/OVnFmV6Bzj1cyI1t7UL
JEco7M1ccMCZp5Rm5S4MoHitkm14wv71Nu1S8VTkPxyGBZNcLTnnt4P/6jCbe/X6LGG29zCYl7nI
5HxZ/ND8sEeQhJUKbezxKhAvWp7AdpcmG8DfQ/CpwwxNPGxJBymvcUcQIhL9l4KM6UpWNvwujdK3
VW+qrfdk+LmAhf9hUMlj7Xrs04PUHZQsnec9ss4ZyuWuHNU/YWo+jGK0T5jryguGMrbhn7srIxlZ
qrPa7iABkPd0XVvfdRBKPFDYvnZrratsY5XxasWNVARx4+rOWAeAH51rjxWPFK8BChZhl5YUhA5f
bqc66pQFKghKRGOgFpS4aFYBMKJyDzniWUAjJnjYHzeSyt78378GhlHVc2ri7/FNFWuUWaJiek1Y
k03izDdMVxKIAFxF0RQ+ousdN6JgYArBy70+PMcsrYAUBdt0ZxtIWNeB9JpYK1lmuhZchGsOrqqw
Hvnzbl3eo03vysLH0yYPaBMggXYpDobauAQct1UpSUDn0nv8VJTvhBaMMTYIWuNZbDPmlu+8gMOb
dLSUXSk9Y64bBChofzvHcbJy1JWP73KDthosQf6IHM3W+43RoKIinFzZ26Nn729JueS7pQaKTBF+
VLVh1xeKch2hfmgryW/USnTRzDzjqEiBHPufy17oSig45PM5CSsG493Sbq39aE19aYa59EsK2dik
vOL78M4wZ8tzyR5VNdn4GDJ1PA4mR4HcaDfEzJVWcoIKVeCdQ6LBSJtUISMl6Of2mhbqDXjAJo0a
AO1wipQDJ+f0CsnCpIMT8R09upJlRvsyZUt+xLn8HkfGkm+DVorZ7LkRlgRXIGEcGqW69GOcfV2I
yPKlaI7THauTvhEXnlKpYFIGVbuHCYOVd14dG7/nbBJU4K9SilGg1kotJr8dklEBZWiXS2RPBTV8
pZsKgRAStigL094fZ9/wGe6zmCSrWA4JmIQ4As6uF8egBUfCiKtDqDl54g2W21QSoch4Y71nHrGm
DZopNFz9IZQvLd6rEv7IaWTQZFUoCXCQ8yaqpKqqO+Z/f4ulA5h65rIF5DeEunLWp19fg34AYWHU
id/5QkNkgJvpmnMkJ8WKkVt7eiUTb91QkhFxI4eipv68guHzkUsRSKbrwJIoqcR1K08Wv7HizJCt
OAPHvasWT9TdaIQXAv3PFA04a+VTbGhinf21M3e7TJtJtZkLwKMS9fk6fAzLf4RYAyP82b8GfjqV
td8r5OVkEZvTb5cA2frNi3Q7HPWV4avenwRdSCS6PCGljoAGge5RHd3wBGfHX644/dOIohr+1Sok
/qSnYbv3rdQ8/WqdObqoyhdmrTF/OZiQ0EZujY/skbqORg5UVSu/6T3v5ycR6V9Bzz4FgzbIX/dj
Tv1ZbD3h7khLBCpfPXdJem7hMqfnwypSc0FSvLkUsiJtl0r79Cqk3r1CaXl/QfmkvXZVVDvjCp/+
NJwF8KOeXgXhJWmXlnlK6v7DFwKuURaaCMEuGqi9t9e88z6FuQ3kacEVm3F5GBzb7G+q4yr2QA1r
jIEOSPpHS9s0xbkfqaVKZJ9JD1QYr9FuiOgdM/kA/rqb2JcLfgZfgB4KK3BYjS7xrZkwJ/BkBuRP
YxhJGCyz4NrkAZ5Jj6BAyaNblYc1V03r9+3KBsxu36pC8SfPeFcMiyFVGX3v66XfznE+nufsDGnH
wT/Ej/R7u12y6/3TS8fB77Pqrf6Bat/JYjxUWUHAWxIdk00dP6MMBpvHBYExgOcQO4Aiv066SgK5
mHHYpfCbPBhwHBMnT5f29e7y9U3j+8ccSHHiEavb+D2vQaco/f6nFf/Ocq7+23ACyrnC2+ukvIjj
vYFHd3P93PGsPwqRvBG3ZBs12yUtvO+4N7vpmyhbuM7zqsmehbz3e+GpeqeSSzlBVB3k4ei2NlV3
B1bJaieG/PSVPgxHX57SfFNiahCyI5nxXu6YI6R9SuVgIYSNIZiHBMSGdpTITvBtd+i+c4p67w5H
V8duxr7dQVoVcYVxQVDcTKSj0RiAxTr/TAvvShcexKrZ7e/el1UuHLllTBwr7AzqDkvlO44L2K73
D8FVdhTU05mZqbG4qU2qxQqlHdV0FUKBeN2bBSJppWVNZ/P8DdqfMEoEg7Rp8W3jlZjh3nb4F0cJ
mXBD8qP3F6yuW6Gso2KHS+kcfFZcHJUo00ojjiARZafUTBCpMPvdKh3aa/LyUgclC6O7b/ig48CY
rh4p+Ctq1HU6JeRUVleB6VZDfQerylJY9TAehAnv3f87lKtneV6FyC1flTIyqzl3PCGXedTh5YDS
4noMCxKZ9QaotVuCtr2dOBVzRQDfAS7mxFHlxhQWni8HXtXdGIfaUqIwjlXNaTdQsYf9QkWzrl94
unQrl1uN5zjkn5ovOZfQihHmFyK2KOYc3FtzTN0kYnA0KhIS9sTRcS5zpmB03cDrLlP/1gg1+3gl
OVSZE1cPFNJru51v8kDy7uGHJ9pMDwzt6eU/ASivmg3HntwFuZF6ZptUvR27GaU6+vS+LDfH1OFo
8jq0/GN7gf67xMfaKu8tAxuyLFZHPO4vTB/0EWaHsHkmeGJtiJkurHbYahssg/EG6AqpMT8GT1SY
1Ep7BdvErgV+jma2qh1eaTpzivSUtc05+UCVd/+qdkoP2QmCnOMNGUS3aKQG198nlcUJpAX+YA6m
REYlW4rg/wzt2w8S7wBFb/FmFZN8vOBEweQ9Q9ee0fLSFMdbsfzdDy8dzqp2VSEKYRKjmnz8RxDF
fZ3ltl0XZNd4NsFQfSled2/uCgNJny5i8aWKgBcnsrZafvZsHqjFSRiRfZi30GaGUyYnxxn33k15
ixTOwDrc5x91tTY9CjfFPREwt6oOIekGHZptJZQDMIIVcCKJBBbVM9Vq/784wzgkm/SJzSyLH/wa
TRXjspFf/G5iZHJsh1Rf1xAB96xHdPx5LFYA7UejEM9DXJxU9dZGtgWiOdvgW8M7SIIHvY+f+TlY
oSRDpDNYFoyR5trDozcyoGSebN5l3RO+JrjwXuPPFGGid6sukas02Me295J5XE2hvsg89WtVQJzM
vfjXJQ1ww2K00u9dAzsElkXuzQTDJyQZtaKoUa/hBo2Gn7BobcVC5L1u7dY9mxlIakQQDPBXAmRZ
eUye+kLftWSUyoelcFuEWUsR3iJw1sHNqfxORmyOYtO+IaYnaDlVkBcZDs9RQVq47vZDJGYaeg4l
moP3EwXiN/JBdWyA6Yr0UkVDRsd7gCM0dI3gM9Tz7EJ6YlhO8JkMjuHFXV9PxHTa96pYzyZhqged
2OyfHNITuHF8o3zbbPUlWF8lIH54D+HxoJDJXV/azbeo+rMUwCmf7vL4a3H/QmBKtODKFNa6Q71t
tHG2TD9d+3EWaZCljrlUh6Cp2SKqCEYw5NjC74cJyNRKYQ4o2rutWa8JF5SKvgdpoeBfvysvMmVZ
qzI5JlR95SG/hsTHrolO6J67c03iULOv4gMDV5NkqCDuWwfkZmlhHzvmWHsFGfHqj72O/CqB6Dcc
HV+cy/bXXaNIboAbIOdc7YDzdgLM9UkS65TzLiYXapBB75RJNC3IdO1CKibpGZf1vdd52nbt9kSv
6UxDpenq5PunQzkfrBX1friyOrGSu1sZTYJX4fFpoquCbHAP2lh0c4G0fpDqgVYMBVAGrY9vylNu
5rXOkcHBVfoTmBJyVJkTcHPmCal11pQMVZL8ARuDU+4uqlwX6y+4LVTWmSRKw/1ftQ4kyoSCidvr
ej7w29YzeiNtk5mHXbFbSjfBMS2Ss66j4t6nHoR564X/+tHWJzQeoHp8+0BQVlR+sLSnNA20+KXQ
OuIMnRYAhnCFc24vE4nVa+C/96zR6LvcitzbBn9sHjyWyjUMoGCGIaZJ9BIuZgCGxKPP5xAZfBqH
DNABlEcCgzTvK+Ekqj/4TBAmXlloKU/pePMMZQIw7Aq7N+ISj2Jl01RpzeW4keHqtQjyeNAsYJJ8
7mEPqEpGA0ySKLvPQSU8j1xTwFUEsHK/w97/Z0aB+CNCf3IWVCFpfrC1naV0QacAxzWBfxzP8GiO
r3ldaOqB8sBxaOC5WVWeqqg8z8tb6n7heqv8+p3abHQv/FGkGuiyaF48jtq6gm/JjGMENg1uaoxT
ZwLoEZlitFzXBqhlmhvAibyU4SkmkFbkUn9PUpdAcWYCnUucXUptAZ3Tx/OiuSKeclD7Oadl/hGr
1vdT8gme2zSGwsuGU65fQw8FJRcfxTvyKH1lnP/gBBdRBNxBKdYmbsD/Nv33n2TDmwQrPVzr9hhA
C5K06M/i56aD8z2naY0FY1Ll8/wkkgAiWg+nNAgooj4dsPn8ipGeawa2XW/2iMwQ9c3UxMLNCmUD
pZ4dw665DLzBspeJUp5wJk3rXUxjQ4aSmKEDuCxHUgKMmxRzhrjnXbqFccEQJzTTATaVFjrZsxHO
uJTt+1uf9RvoBR6W2Ih6Z8fZZ6dW1lqjtTxcmh/528izXiQm4zos+3UAD7kIgV+E1GORoi8SFkBX
a+YZH7lKxScd7X02gioaIOL+j7VXW+Vt70xSgEmR8y4ocwc2JbkBjnCGPpDn5Sm3EvJRhIL5rdZ+
tuFBubPYXbyiw7ve/qjuy4x7L806TNaPnYW4CQiqOfO2zx5BIXdCpyDujU3UJW0z5zNsMmGgxtER
DXoIvpZMDnRbuINTuIwtImGrgxz2IfJsOGc47IBM7/7OcWGI60lREiXuvEOGJtSY+SCUTc6uNp08
OhNtcoHJB48whU1vLB2Q6gtMLOhXjQrhQRV+3/Gus9ymKT361yRAGkfEeGl5mUWhUuOY1wSXA8V6
jHsyFalXttcyReszSMoWoC3kRmqlzauBKLXQ5EVF8qwsz5HC0+S6OUglhLon5+T/esGmze2nHlgG
QA5jGfSwrSK+ve5Pjtg0Ok7THGFcjzjQOyZnDsEbmcKEJd1nZZ3uMjUPTQD7sb8b0VkQ5yelbD28
P76YFEx71lflLOzPFkV71jfDyyQOvm7ckCK8hDXfwaOyTFmg5YqD0/hVfGAMAJloIVyy9TdkoCxL
pbDNjbs75CyWUBlGB0Y9WZRGPdoAexHIi/GhXfQf+zwzk+y0jqkJ8GJ8rHGJo/UXr8Hn66g3oXUz
NJWvTz88+47ir9LcMnzUmE4OauPdEWY7nVy4Cu/8ebewgxoUIzp1+DDuzfOcOv2GmhwrT4LC5s/4
XRC1HRlEfo1uwJEFw6Kl5A+PA5J9b3GLG0xZ3cgyY3RbaAczI/FM1cgVRVpONt+ZNbTORLFnPDPx
knyBRsV3GE5mYYuqYD5hbxS4e3gwQHzDuAzygh31tODfbDkFOOMjYRTJdV3mrFUhIlDCO5T+TbzV
bGvYQmHZU5Lx+qgwTlu2kpyOSKa95z41nzbVTUiHEN9M/K05fciMUh8S8cgAfK6h0KyMdnd8OUvC
9eAA7AR0OXGSGhi+27uLciHr8vpzc0MHSbhM92+c5HfzjTfw45nWc5s/d/wy/rg/Cn9wbbaYIUCH
4/04/DMTtBI1U8FtumvD/rjjPUVDFxHjV81I0Dr24/WR4tUMitiHOgknI7yE2dJL8VDinCJRtKd6
L6jJ7MOPjws2HXPsYV/I0RigCfGwBYeV2/lCeThLyqfl4q1E+U+8rN3mdAmQh5wL5hqsCh7NGee1
w8huf2s9N0tiOqiXEQlO7rhWQ+9mmt0XGs+IA7SmPuhrTlELY8UxCLW1IeqZwNEaTjLQxIzsIj+h
BoVAr1xCJO0NJpWWQChaG+4xz46MJIbs6b4bMo7eaNloNvdnJRozmB/vFBDsGoM1D8MuHNGNqHes
Z6dyN6ZXmtzA7fLO42IcJonhVaU7xxMATYJaqKoRYdBoP+4Z1XafayaTgZ8GaSNFDW2hoDO24Ln+
jSuqV5PYsPiI4zolxtGS9hO2iGYbkeevp8tz5Av5Y1U/9XNmL5VAekzcytL9pFRGGHQPWU7/Ti5E
XMCzV9pxKgkrLf+0UBwB5pO70xG04/tNem14pjIVgATlzmXaUS+2W88prA2VlJSsLZbQJVlQ8Bsf
NDdyfHhKxXqhPtQuoMZtDeROS73pCWtmhMiElzZ7RNwm2Rt1OfJYzTk9YPbVOt5OglEN1QzkLmpQ
dV4I3PIcSXjkODNesTqz7VOoHTGB8UhCWzNUr5057JqzgROlCaBuYhhj6CDEhDgjaVfkho5WqjL0
zgnIitMCvFSUD/9xaFJzshsnewQ58pjMSLT+Q93RNLqoeU0lggSrPA==
`protect end_protected

