

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dk2lbe0Kq4fQU9wJxTwM7nrkKf0wGLR5vjo5hNB/iBdEEx7lQLSDQZQQjl7yoSnl2U9k2tNT8PI3
yLjF1Xb0pw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TBC1mrVezvr2GlJZKChgZflcOacg8z4G751EQIGLwtp3MmMN3Y0N1o60lw63Qd8x41tPcFv4653w
1DMznx/mkGzWcxNBivOG72Y1yrqI2/pxzXYLtIN3oSs4xMARa0CGXVKNM3JDUuy0t17O1+RzoM6+
k+NgxvvI7Ts93e4Q+GE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W65o26/G1ZQM6XpDwkHmjJ64CaYJAzVLM8ELZKZC5RvC2AorgSzz6M9PBN9UU9g09E6q0xkqn7rQ
hgyLAhE9KvoEUToBxNNHdI/tFJ+Mmrx2pZl9XEmTHl2VllusjMc3YIbbgEsweryV2gRe/DpSeTCv
8FjXn/T+J2o5My7qpjn9P6OIyZC+/+Cl7R6OybpZugyT3Bh3KJKi9QNsKYHb7c1XsOXsxgyrX70J
Vebd5CJCr2gp8RsC1k8vX+dnIe6ZS4TaXqm5M2JkUU7gG+y4SGihlWeRC7bTwSPg/ZDfu0qzbh/B
swzazvc7/3BLe18XbHKJJ3gM37mgmqL9yLmMzA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yk3Vp44FfiFRF2d9Sep3Je/0HHeOKV3R8wFvnsSd3+e1HZIGii9SHbkP9Xbabub2KOv30Q3Ju8lo
NTssBIZg8RykvF6X30XDZ9P3cpa/5C3Jw7mSwF/zD6KClFjNtKEeksI8ZaO0ZoZP6R+yEIKKfbNL
6Z8VI7Rm5EX0tN3poak=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mibbE6Jw6GWMgRlNutuVQgb54hm4/6E5jb9awh0xn8xsIHtf80uo38b6GhbI+BzY1OKD+xdxPOcL
AGfMQMsR13EEAbePmQDYvV0gSt6gUMCbuwx9LYJEjrtbrxLXZpveebmwQukLDZPQagKokh1phmHh
WFWEV5wQ8NKnAL3SKzABPobWtT46FDr/qYFUuz4CV4eU9omMOUi+yfbFBKpJl2HZBxs9kA8TggyS
56IHg95/Xs1S1z4h7yBHFAeP9QCOcG3iGRLukF/U4+gBbtCH/MyCmcXkBngwJaEouoE3Pk23qg5G
/C39sP8cJhUW+ZJzUcuEY5QlK2BZTSoXFgl4Fw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6144)
`protect data_block
xtz3goAoqav58ey7eg8tou0Pn/ec32cSTbr9JH/GOK/0Gkfjqy9i1ObijObS+9bdb5/00/+l6U5T
uFyLdHf1adrnbcPmnfSHYwC250jKAARGZvGpfckt4nLsiAUbLs9SSu38xkpsoZ6a7k7uYgTjSfUQ
cWBcX44Hy12RxVZT04yuGyNKkzI9QRW33hgNmKdGoV3Uf52RwQwCErqEznHK9Z0TwlRIiSVRHtbE
swyL59DGzDSEtkauvEnBqPqiYTT9v6wOYDt+srO5kosvYAJ2CFd9duGnDEsoCmCufYj75RHg8+Md
KQbBhxBea7EnX4dsHROxUWi9sO5R0qxnTdfe9StX86Hx9rZpNucoImjrIMbHCgjtBbvtptXc8ABQ
zqzw6gmGB7SigdmILaOCjVwaff72MVF3xo0OcrfQ+Cv0U3GLeUUIEPMtT5nRNrzn5oLyBouzzTJo
aZN6NITufjT4HxbZ6rLP3XnQiXUHK/kDuDpIHwgbHQoP5GJsCwI6SxaK2VxioEWLCXbdpXKGNMpo
kPhUO3NdPR/+jkccRzBw92BfioPdxNe+Q3i/JT3NIuvoybLy1gahwQYJ4mfZDzLg7PRkiOOn178s
it+sSAP3Po0Y+gABhln4Ope5FZqhhYU0ifKfTjHTuD3+23ET8y7B1yabM1+pt+/7X/oui7iDtMlz
1CO2rle38LPDGd6VaKHfIaYeDbLnevvc9C3JAgOtD2mixbgiI0Ddoe5sBHQxRAWFDxfEmeqKMrOp
rwQHtJf7R6a4CAPFu22C38UXmZll3FoJdps3IoT/YUBOmc0yIH/V2sDPT9E6ZoQ+sRci64zOVpFt
Rj5j8VCQreRlxoh+b8DzFhmySpATzs+je89BWYSjXI84X8Lg9Cd3UuPYCMSuLxh+tWHTJa/FRq1x
FsNwaKHJVtpoCBcfxzVwIJFLQNHzz6hJ3V/kU4pdgWSY0a5Txr6jzPjHlp5XzlOgPK5jAYgdCUEG
o6TFC2+4UgdctD6rCBhBIZh7QxHlFwTjJt7Z6sls9aa2cZI/YGO+IYUvVxPDjdJt2lYGr4tddNVn
YdHI9D1xY28sRphP79IoMeVl/xUCkRQHwC6HT4ClMFtmdq12vmhSZN+bLOGlKMygKd2t4SVBXj3C
9NFw/GdWuDjWHY9qs5ZOaD8u/pmb+KGQXY9mieQGIX3fXN+rKqH/2JmRHngTZ922TGFCwuQSv5FX
DM8+Jpx67paZ6gdOvb7SPPEvgEe5hOHrppJ+V65aEFocI6FzoF9mKymg8vSPsNGzEFuzqREUzqp4
KiRwpO6u4vB/bwYPUKbRFYqYRCY/heL5caGEryNvM1ptr9OZPu1yZdVINi/BjPuWWWJyGO1vR+tP
OA1OksWNPg092fo2rA4zblzaZpoQ5z9yQJ7nkvua2y+Us2SUn2FRclK5UJKHxAponqESOJKeY19s
mEslg+w5c51JwpUrW2zWkVMjsBzCRKEBZC0wY4ggSIwXnUs0ne2bIYEDQInnn6QS1Xzc3+d34XZe
uKPJVFHME492JfUw+Exr2OPF920Ic3ysdCLPhGe2k8yWc8Ioea0OiBdBcewggKBj+8xqS9UkTEg7
UaFmQKvXdtqPp36y2Sp1T3OHWwnzfLL+B6rWRVAPKj2YLTRFC2z1mDtNQTk5q8Z4w0OwzLJ8Gzbu
2Yb3W91hbEfx5RibxPiKRJrVnkUjwn6ITV2ZshNVLuzgdymh7PFK7cvN4GxJ/ljL2KKkLOTJN+JC
T2fzEgpnTZwj5h1c5+RCrBD5mvgnTjQ5hxaPUmj7x/RPXlqXn/iHx6Sou9xCU6fV7v9+xXQzoUoJ
Q6f9w/9aWR4Lb4wfdm65W2C1p1MeR7FUYxqRYbqEi3vmLqiQ+0sFOcRnlDUjLgRq67IDdJ5xDT6O
PHlLOXOjsBnPynGNdk01NrZPxyVPATRY12Lu4uihRzpPYvS2q0KAqOb6lTMXJ5fCJ4wBVONJkpyc
DK2vnhVcEO7TW7wiSMebyu0dXb3Xc14tn8hLR/9TUrMqltOqnnAnNn1Ro//7LWerHXEUMKOoA01t
Qe38LMZ44bQT48NN4IAtIekHHzgQkpYMLIi0h1kXUQn+k4ej+n4wRQD5i7dods5i8qUehtiZEeEf
+mtCfquZCeVcTcgztCrmgKtJPMvih4tCPfb97Ej+EGBlRFhnBoTg7UwH2Q76x5Pt9BwDsL9w/oDl
45EqYEnBzcWhwpkoHDPB9Qvj7FyrIz+q07sRNuhpwAkqF6zhFC/PkNKfn7iuYdJVTWO0z7gEAtRP
IsiSX0+FCd1v8r3XNp6B2SRjKifg8/z1XvA+uG2qbG+fWijfDw0QnPVwfWwFVQgOcgkd/Tzg167L
XE7pt9X/j767NrHO5ViKc2Mj3Y/3FpHgwa1IBYi/uH67tO22TfCXZcipF/s+iAxJtFR4thpQHiGq
2Bo58yYosqOEReyGFnNOazy5HcIMpiqRJed+4TH8eOlBO3lO7D8rF05whpy77lh5SIcpgeUb0Jdg
FaMHxtLSHJeywvUuK/U+upMteoHnOGxxCDlaX2VWUQH+PtwKyCsTXN8GMZo00ktBP38QJTOPOzWb
uBGcIz9tZAEpmvCA1CAhgxWiLxm7a6543htYk9njY2Lc8XOw5ElvVSaOSyqyhMJWpwqwMBkxeiqY
tDFEUigRqEvNTZQmX1QPhVxp0/YRCCZUV3LYX6bMEBele8RZUW2FgZ0HOzTHKr16Yx2MdcB7nxbd
OOVAL3uq0UFS4aTeZawlvPNqJQsl0poAUlgysT9LMQsgBdV39jGWKegwvTHZ/+gqPJkvLAuiUoV0
K6OgCHK1o0JQTNLvGiMa1iL8DEOa5lZjnFQ4G7bbAAvlEI4+QQu9+n+MERFK2vmLec34WzHK7ikV
7Os6buyydmEpkYunModRogIBx00P8XA4cNewSEtIWzcQzFu3Cgme1IEMgJoxvzBgQQxyhimbQpEz
EIaZ217qAfr9kK+0ZzEwWZl6QP97vBRfFgBkODr5tRekU/GZPabUGVbzSZ7tVqQY30rOhTwAweaZ
9HU3OBsSh3oSsXzd0X7ciLVE3tD2EANN1bV2d3jbQIEOYgwXG0GKIYM/69D7Qfo1n3RNBNpUkGYe
HC50x3aIb2AIHCJUrBimDvKmfW84B1NwxgVFtekidGcVJ3xAWY6AnE2dDgO+JJYgIozkvAbZANdx
PL02s9QJlrWcpjyTRbtSC43OQUJ5UD6EVoDpCaJK6LPDYlkadKs5IrjyhiakdEdZbpgh8fEknxte
ONuu7JQGB836YYBkUa1RYWaIbNlWVPoy0L5lUm5X9OueGNsihaaFyl1xfy8u/gJpRxf+gJQXTIML
K1O9hvz78RCOzxkH1Nc4lg/8/mWLtLE4JcMqlahV8MZei8fZ7eRAE1E0qJIGXQYtluhhT9w43Q4u
lnjIhKxD5U+1lzDIk/7jbZQYo+oelu2f2Bvqzj9+YbjLXfjbsnpubYbX/oS/EkITxg0pBmmQAb1l
Jg7jVD+yb6hv7v6dQa5Lz85IhDKuiKxwwTaPGvJh/A/wmcnjeRZjZFmP/gelcbqg8rvUQgX6srlC
Q1lDDEOnKnJ7zOseYNsAat69MmK1N/CuOieC/TXUfCf3M9E4VaE8iQQ7+27tes9xn5bB2ABw5trN
peio4dKVHY/OG3sVZJDDKnY9G3xCtz/hyq5P0C7p8zh+pO1CXwWdonRPBdSao+eM7bl6fGmSrGYN
HiaraIGAkWrlCwcGhKVDJVnBDulSTAPaE/84ZW/aL4tlVj26tl5zkMqwbz3tsV9F2McZaC2WffI4
9+1IGcao8GdbsdwtvzgtYT0yEALZz6lgQZhaB41Fs7e+DZuWBdBdJEfF4jU/0achAQAb09YjEAKU
DtF40sq02ikmWt6+IojeVjSCf8oMSdnySD9bHn1cPhZ42XxsjLltonJUykCDGk17QKaVqVQh7W5u
+ucdVj93luVrEKpyL7Xbad+DA47GfQFnhu3D3ojyZ7RfmWfuet0akvVKrY8xXvybmgrwe3qdVbrM
BI8mDPU15wl5iRvRA+O+3hSKJhyH7znlFrzgabAhGqWnlV4fLz0neHR0A7GNaulvd0jcDpohp6ny
EVblTSDch6JQnJwJBe9arefzTpt0HZemEhfRmq6xXI/zs9v4/GnRcl0u+EbBjn2etBCqPg9tNRl/
7mOj5nqRhRuhLBAoWjkAuvgtwWPcT1jbwA22gE5ZaDfQA0hwfgx8Liqb5arAJZrOvPXi//gZq895
9iJ8g61oKr4ks/pVoFDYOanKYOW5Ihe0zae01XutgjPJjvluo7u0wGaOcJAmV2PWR4DU26JJPold
GtG+qm/p00WfWgZN9GdEruryBz4tKRSrlTyc9gntVngrfwSXozsrIZYyOq4ou6r0ujByFVP0i6dL
+NQ2yfWRFBWhB7vB4msvZDLhnr4e3RYYonxe4I/KDSyj/SiibKgXdDUSEzUMmDoy7QVcYtSfQuul
qquRqCgDSyWR9x5qMpva96i+f1ehhuvFsUTLeuOX6GXSLJC+Z7XtNBcJ9bv/Su5+JqW0qpnEYvFH
1E0F0Tf4mKxFycbjShU23jGIZ+xCssdEkpKqiEubYmC4vR/xXHu1qgjejcfcYZPyGytngoDaH8Xl
DXJWupyivNXH0N9OfB8h+0QWMuDk9cGFXqQB4p6NTqX9BWkFslg1hYw9ijfc4uotah70y2DaXHZY
xjTiiYGQgJXRAQBg5MhsXBlL5U62McuF854CTEyCWpMBapRMBGkQtnEEQ8QVDESUk4N/TeF0oKn9
wmWXGiJDx0s9IRbLkDp3IVQwWBTD4IdMIH2ZVQhjQhUHOELwuK43gUWCCGgaJm6DFVwbNvrPMMPW
+A+xBZ952JF1woj2fuq8yo/XxrlzcYrtNWFM65Z7wWlwRfgOzCqDWFCOzhrV47tQ/POvg9E1NcpC
6CotfcMoFRjTEvDr75wZ1o+L0qnnMMC0wdK4vQHoc9aMOqq23gq6jtg1eTRz5y7Wz3HJQLml25q3
Gxtl5r9vtdsKexVPZ8D9HCwP2OCMPPqV0omi03D+zVod1wcjRhXFUNbrqI5c+AauqoIjNspPD0hb
jOe/Fjf3bWG65Dz4g5RwVRcInuVliZwHbxI8I67UNJOSjSXrebUsVgU7PIBIDZ7wb+eRJKvvLwgI
ktCmwm8yqQHWM29VKgy/UDfyeXNwZ4E6WtnchDPOMaOKaVt3PzKwVziXMZSClWKGcETg2mOxsS1I
ZJ/QW/1b8HduZxdGvO1qsrJJWJsz3acVJkHzTIrPvwsFErysZNzCvQ0iZBf771PyF/ucCjBpBH8V
tVJZ3v99R6mhDE2d+BWGBqzkSA0v1NBhtYbGd1PugvI+ZWhpVHGccqcrqVYfxiZ+Jc0ULcpXjx3S
He4D6wjZ7hTYyb6rcboQ8E/ehU0oFu+gxXLiO8rpZWmYU+wWzQcMw0DtTduL4GFhKBCIq/GIE1IW
R+MLAQb4CKH9KuiGp0ZUtnvXaboJHpD00zDt+Bgu3pbVGf7L9Kkc5ktRT7POFS7f/RILvj7mRQz+
5sQHcn+r9nRfMUmywN/3YshbLCACNwCJSjeqp8Mtx7NgC86U1Dhj6e9b2HD/ciMDVoF7Vq7c0Re0
6CYE6s7aFBbjkzLYktM9cHHjDTgABhyMGYAlvOAPIzC9DeFMLbNuyAcSL5ypKZRBbFeUDYWr69cr
1QqYDgcf4CnJEIyl8ggYq0ro2ibguC6sNgwsb4FWXoYq/Edzoedn6QlD3hpndHiyWppLDHArPZy3
iKJKaTzCKdiNZkwvH4v7DN8XGT+fPeyJocUCHu1eb0vJ+x7AmIiwqQ5i8LMyQd/ilJLbs03Dk63k
Kr3vhkX1RiLXe34n1CMjcw11VoYGMRZscWeGupA3V64eDk1xr/n2UusqbXbZ9Yh/nyXoGJY1EdNs
L86GT2jGvcGSbqV99q801tbV77mAYj607BGfnAq03pL+pSb+Tn0BKBBaDyc67I2Vaal2QyW9cMAq
DL6F9UqJ7VwFUlpDuTgB1RyB0w7YGuEcBJ64IxNpJIuyfZ7tCN5GyY8OzjeYEJbAvUjEt2nTtTHy
jRk5QRZpgsJ1Pq/rulxpUMSVWxkj9p4ykX0i89SUEo3CufMzrQWLnIUPfiAqii7ey9TK1rYwwgnx
rCZgNmPCCIn06WYwauYHck5sbTd+U7Xj6qzzPc/nGHhQPyP04SFEIZCAqQYoxnhr7li7IFyG8COy
8LaU8ZkEelX+bNxw7CmS8fn6iT5jte8OQbLPrlFEA1upzPC7cRV1Gs/DxWaJrLLkRAIWGP2hIDjv
0ujRS2ueJIu/jD3SDgpUsKMhlvBXqFYmzJDP+A9jzL7veJZ3XyblfLDsvnpYk2HAWlnYlqnjyRgB
bMKybrBtpESTjTKKkx9BPXAZbP0dhoUgTnjgX2KGTceEzaYQNKob695whXGyy3ZklLPLihBfDz+p
OoIgrsNAGKoKNFBSWEVGf2rbKxgytml3ZTSif8x/FBVbFgy0ztjDmUM5qHDde4ca9POs5L+DDwpU
ovMDqxP/okAhLh9SZSDV5RIhvFOkHhruCF62hB5IF0P5HNeXS0u4T35cP1xxpkn4SFEkSbOVd3dF
3GaN7/z9yE8quTLU9w0XzK91dIPkB6ZPd9eFU01dz2mpGoPMAV7r4qHV7r4Lge69fYcp+ECZXNuM
K+lpxPI8tnHTJib8/iapyHO3doFHT0CDdf7UxGxt7qt1aYvlvtHpBKg4iIrKiwMbqRAl76sWo+QS
M5rfW/ZO0YR1qKEdIRU03SGRk+Ja6qtr/HgAdO8jqlYVIUpGej8bgIF+eEsCUHo6wS9cqLBkuRaY
rhK8weGfMQ+egBtjaaooBqa9DAFk+9eQYcWcExJSgGQahZX2W2p6hElTbT8me8SF6cHcemxJ0ijc
XCrnaU6kdg6ikKbQTVw1J2F3MM4n8M9f1FVnq1nZnTOolAZYW2K74pMR87Nfu42EcuAFnrofdEZo
UJsYlVRTvID/wYudNd8bwqQRw/6I8+FXrEr1+NJ5Vhts2bSmbJjxI1tZhBwwor7KEPdim31I8toY
obBaY/RnR2tCJlm9y3O0HXoz4zhVZxEpm59WjzJGZOm58GBufLO4egXiISeNrCatwIw4HYmCDyrY
wUYynPiuZ5iChh3u5S5Qd3rZQllm8I6jzneuQKdntBhahggtddGcWO2s42KTbf0sh/n60jDNwAno
gLYEoodWQh+n+iOZctURnq4HS1nQ7uMXlw1VZNQUiyz4RqGZoKYY8BoIHNC5gJJSHliuOXek/n5T
KDYicpt3M/ryvFuMz45vdoO1oN1WJFqmN1MWLcyXtDBRK+jDZ3LEYMXzP8QSUbz6ZG4b+bYM2LCw
0t0C3YCYFYHnRueKSn4Sn2YLxjEkGY0OlErry/5/xLb5eOOlFPzmVDUL1DCnbiHl/Y+/3zNCuUXh
/R50BI21xdn+QNhn0wbSa97ANTV/gFYzqSBfj2SHSYvdKFTj2wL1scLaE0mT2kBmYU9GfQsK4EuZ
gGxy4rI+IKQQi4NQUcF6wj2iy1/bZM+hPfbonAGkTfiyt0pDErB1QjWkAwO2hZJGVhA1x0k+JCrF
zbG4Hx3Ym2LOAYokCZ9mHAV6hyN00MOtG2Ml8FRbHKqNU0oFn5+EX64qHlLpl01PI9HZwWXpArDj
e6v8CR5intxv6+95z/f2j3Az9vaz/vZ26Wa/5hCud5st16xo0Bfovu2vQRCLar1hbwlHZ/DZWz8P
LotY2ryzoUqTeMq5oUUZxwm7rlN7PS29R92UE+8HbGkT3h8+9dUieFwgzLavSFcchRXIKPnqOIiq
7dR7g2yalEa6gVgXo8ZRgMhFuY9XpkKzirV656ukl/fqkyYaoIqOlvdgM6zzjlr6V4fWfGPXsff1
gAWm1AO0Oguz0h6INaBBoom5QlMQgeC3V77PurubQZN8HSM8W/JZNjlw/ktsGl7qXLiUIp37J7tD
+EJFXvMiLKkf9xklACzc4xigBtJIKIL/pwSDPAWit3boo/k549ViL38GDN3ps24M8r67IkX/vcvJ
oe6QFNeSzNrSlpCIu9E9GJ9/HdJ/eu0rj1eiObetezLD/wx10nQhsmpFfTbQw3U2ZAe7qGPZTI22
74xyR5o/hsdFF7aqJa6YSlFyd4MB15gPyZA2UcsMzqHvcBYv24SMuDMVil+q
`protect end_protected

