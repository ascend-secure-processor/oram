

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MuNu1vhM5iHBR0V33YgeRMMRLNOTGvNsJKgG2q/c1QtZpdCyI6tmeE1Y8QBcA/OlQ5qbzKaAr2IX
cQOyz/9AZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HXfGfOcH213+quAPIWX/yNq1TzoLOF0lEJNAKSX5mYOS64DFesMTcd72/eRNPXef/QzUguTWMOAC
mD/xj6aJGHer5XrM7QLP4YrE00m/MBGQywT/z3vwZKS+PngI3SMlzevM2vT4+psSo2mwjFyH7S0z
av/S0uAIpSgReBGGLOM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u6MhzdMnY8By6h6lPLT6m4gCaiGMJj11dYCFRsbwJSMO6RsC0fIOaAtoNBn+u7eEeapGeZ8evvd2
VDY120l8oDdOitkPwik4nrm0QZ1LBhGgSxaQOA9zF9ljoWMXS+GqkQOQgZ3gVbmO/o3Naq2+Hr5i
mvjZOiroJyFeDagjQORn30BOkz7eS9OfpxbQ44Xp6PclDIdu/Jt0H8kkXkYAdQzK4k2XP6q14aX7
/QQJy2WRBy9PRotlD+4Wuu4PvBa+8hPaskEOJN0Do6Q/UqtnqjsRoVbBn4rbdAxdWegX5L4+mLEA
v/LEicmjsOwDrSc5EsPZolhpK5ezF2v2719aEA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rKFJyiR4oERgoje3TmCPew0SwFEV9Lp/Njbzw9qXIk1qkpa9ASIQ0Ua/qyM+xpLAcLAUnLnarczt
TJaqDiLQSC1SSyWNdLk4pxAiDB6TzOkmDe6tXL6/s+fcp59rseS17kqyY3XO4IgdDjFPgEgKq4Vq
4N8GGfGAvrJu9vLq/x4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ptspXwMpDNCngxXkTf7s1fs7ifynmA3PPElt+JG9iLVPkCBHJcifroVvf3RU1Af9WHKL3pPVpKuz
Ab2+XcZOzXFrpwRAUkZ3y0F4efrhERiftdw99wsiXDLOr+yJ+3Zz3Yl3A+jWh93yjidKgkwLL/i1
cWPM5gI/F8lKEc9FlV4xsdUgxhJBd9E5FwKBpY/Uz72wed/SWqkom8FFWK7VIvAxIRCti1n+AzLp
S4GythmuWyRS1BGwOsjm+/Iy3xrllgmOjv4NjS+ArwQLRjkSjvuVHhfpPDkwNB7o2XJhlg9PksxT
T82/NKtrcb6mmEYhkJFAdaG5ezMk/g8H08bffA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5008)
`protect data_block
leBtOP0yEk0ZFRmssGtK7dXD440fydJe8yAgjMDEvbnXxthAhp8otbyUPQjgRI9IfClSISgpv4Li
IDeYLRzq/5XLxNUqQ5jD+isGmN/LPaCgApEhDTWskf9riNJE0UG3rA47qjOEx9gvZyRP1ZTFDVv4
g7hoiFIIPhcnyM0o9+W59RPEXPzTJI3L85BHTr83x9i8y17acEeVorgdy2TikpfkVx5ddVOal2sb
3o+srXslrisuw5yL7urZ6gy99eRFRZEJzhXHG8oc2U/9UUwKggIfveu1fm6PNciqBBLISmwWIaze
9le66c3nNvHldXYZVXP//OAMGNs1S9jgFrIGRcdHKNwrpxY+WgkMBHZ3aSg1d2dyFQqep5p4gBgz
oxxXX91YfLX6FaKeh4J3yRYpv1ubcwyFs8DeWZdNoBDtvcFl9pykAY3R6GrOeZGAexcyqFDA16d4
vqubVQHXGXQPutoWy84zF1n4WwtWORaBSAaCtpjJjyzSIi6ovYrcr0f6AhDR8L+btra4tEh1qyXw
XpaioWoMlYRWX7h3wnCZQHaBTKBmCA2GHV6bTwVg70xYI9Xfnnjmux/ZxBpDOuzQso4wPaC77Ev5
b2c1Lgymd+OgTw08ASNSTzx26/+caKxClQ/GfKdh+F5Jur7pVBW7gk0Dt0LMGqTF0OeM4Sm+KWFY
3KTG3c4gPJnjVR9/guPxGVw5UGuwVQcFpE6NJA3Pzx8UZAB3qNoFsT1FIP7GWapGn/IgPWIxs1ex
f9AfJd/vXv5pWoA/AZrd9sIqPHGouqZVPbzPsW0KTa5WA5JlZaXh1E5pT2m8//AUW4EXw2aWWchS
+N0rDpw021Dia0MEN5hzAjxkY4rW0UOmd5/quqjlkkB6yOoW4JrG2fkgmmRurxLdXCIMFagCxm5r
OgP5ttKSuASPLc+R9THkb01Ek/NLT+zSgWiojIRut4+ZVOC7CZEAzi+JaE5/G6iaAc93NuVlc3cs
UgFYIbYz6m0aSLib59lBmotCfEFzi4XBdZ9pfOlxgdQQlq44xRs2SvjUyHiE795n/xG11/6QflUg
qW+5kTl8w3JaLEmZawrrNE093irw4YlUdMDwmFzn0GELph2/kPYm5CpqMH5q7in2Ci9uti9mB4kK
XdB7Bn8MIm1d3D9MbgN8EZT79qxC/StEgiQH1Bqhz/SmK44P86sKSxmVVxMcTTcPaEm3gGTHNDJM
eJBsI7othzGtSDLvRvSOPitYgikQUkpjseoYisSrU12ju1o1li+aArFXiyQBqAYx52habZc0tCd9
PmtYvGq4VcMMobxE4YNNtoh2Y/GJVBNd2atpNj6wOituGThwTZFT5Pljrs9f9pKV6mCzLz0XN3cZ
em58u6sJtT0m6AYGuyN0VHCECiZahYWGia4333uisjLWBRV3h7iOKbPCWFBbhqsBfxKyOodC3CJu
k2CM1hRU861xg51Hel3/bu8ipKhSVMZ3ohB2tG4uEtZQa/f1T77BbF4OJ7FmpxdpNu5tgElfYlC9
8aW7zdTyal1bL5IuS92LN8KhEgEqaFqoEP9O/jnzhZx5EEsRkZ3JzDN0Vjru0e2O0hLLnzobLEzf
MYLjhOXQyL42/tYRIU8fh49XYurpf5kiWKE9C8/yMwt9ppbmEV+n8nzgUG9qv9Xl+weMRN6XzCVr
QrUv6YWToRztO0IIFI1b/h6WJh6Ux6lW1jYTQRem/npJhoCxVDfbDeYmlJWDBVF4Pmk6PeEfRUpv
HS4T7QS+NeVWJo6BTgjsvxlndAl4lKeLI4GwOFfLTnFdikWsQYTwHjQhj8ULmlYcgGtPn8pRfOjr
SIH201MYaC0B/7qdjRBYDyxsvWfFsFr3nRBO1XlLgr4fBZFUM1A+OFecT5SXsAaZDYQ2fVAOcc7f
/s59QE1uaNDDGID1nnL2nfa+lkWHQ2oztnrMrjeG3i49PotOEskRKsxSSkv+x5Qp19w2jbMrU0Fc
s0sbGtcfGWfaaOgbWIpp5UDeq9ALVtxW9tIvkNh/sGBM+b98tak6hvu1BgefahAf1k87A755rRGM
28UwBz+GYr+1sj3kqXS/vJ9xbtXwoLJuiD+Bk7oXdtKUccFp8gE91IZ1twL5+L0o9DvttPUXtOcB
tcJEnbVVDfXOEcvSyHkJUqJkObflCHOOJRUInuGoICnKAFa52Ix9VooVS3wZKeaZ3fPyQIZO3XSH
Y39UeSY4PmnaCs6ifXePwFW+ntFpMdKbX6p7QXSEkpCRdYQqe9rzjESw2IEEehtngTIWAq0WAl5a
Fm/Mz3NOD5XR+VY7EF6YjwxOWx333X/s2KHJSxyIT7vdynbVyDHa5AdodB/C+Q5tnuoxxmtJ4KnK
x9T2EKnc8LQ7y8/dfDTHmtTaHeonjGrnwDQ9lkgfTkLIJYklY3CkDoN+iGrldwCA9Yj3yPt16Njf
dgsFhgXyqGFmGFwFgAk84iRct35FEAouJXzImcdsoUhrK5zhrBhGz9DrdE2PFuL0319HjXKDi161
HDagu6jR2benSVe/CekrW/f4I7hX4S0FLuiQHmq/pl2XUTRn2jJVWgHYtSuKeSmmUNl6mhP9lqy+
M+Z2ktE/9HfdL/liK9G/qPPqTueIFY+zq6SsE4tREPXpv8eCQ1e3T0PoAX2MaFTqD7c8MvIFxDLc
lzwVivHSLjUh0JLMPQW+zeDJqWLMzL3q8KO0kzSH3R7yJvBs+sttPiFKu7mqmYJsZVMYIMpppK47
mSALOHH+UDdhg48sxxDbUWK1+yeUocGhHekGU2d3NnPMiYx0cXnow3EUSkuO0C5VC5VA03ZODgbM
3by9BkbNFj9jeBkDmd7KHs7W5jGmxzigZl+v59YQafEi2cJm3KYq7dfX6O9hXpnCLZ6BWezRKNHi
xQVMVJxF38djX7rhV6HBjzXH0xi12ltbqzKB2j1ow/ZwPsAbPVAOCRPvLpXGrgZV+SJktl9ustHs
VNfzbY/yBLwAqwOpeYpbutVuXn7bi7ra8efENfdRISwD+eJixRrZ+VEFFCLCY9xfqcdUdpqR7UcY
nSf8nf8X+HKFrCy0m9yhoH4LVIqL/IpV84RIva4C/s4Fyc+fwVNwYJUB8nHHsI4h+SVg9NI5aoxi
7GHUaf9q6HBoHCAjycl3AcfA9fOeW1yjFuuoTVjZtUqoj/Xi8vg8lmlVw22qi6CAYkqNpndg+AF0
j8EAQxY41mldshQpwlOaoQxjvzTuZOn/IqjFC7vKe7oqAHJyf3p/tYCPT0EEROB9vTkHWQNBA6GO
v7H0VUywW4LFSsIY4oP7O2mw2euYKFQoMlHjfpA4I3cxYRQEwSyAawFCmFkxtj38ydO8A0/z078i
HKojf908k829ID16hAhXPmio9IKHw8nPFnHvs/DHKoB0/5Nza5l+nRiIU77540dIvCVZ9gdeCHaV
FvQni/R+1ZvYzhwbZXp3dKbL5w7sMAHD6b6Np8SaV/fAaLl8w7LQVs5tGbD+1erKto9J8dQ2oD67
LVz2R8mig2UTzMT2wnFJZkkU6YM7++XvxIJeDZ52YeVEgoXf7Xwu9Qct6Uxgm7LnamWoHHDNrG9S
5HZrjNTM6yRHubf7LyBi/iWkAqBQzhhDIxNJrm0rb+fsspE8ZT4NtW6GRnwiKvwEmbd6rkvPozgr
K9T4FN38FJXGeboDbTU529prBV6g4CKq4ZC4qy9ywXVcCOkr4azeB705/Q6ZwnbzlOH+7ohbQ0bV
hWMfkQiK4UagG2dIovkJr7qKUQUo7H9ZCOTqnz+zIB6NUd3M1oFaLl0GMyh5cQws9fqhqAdQsoEe
R1AOU6b9iD1xMrQtVcrkVimfexzhPaG5B0/c2J3b/nxZRI30wmYJr9rheGDXsggFF8OLsuCX8RAO
Kn6UqA3UMpdFkEsfBUe8WwZ8Pc2Mm3ur+lcoUEx4VP9Bdz7MIPNQFnyNs+IgndfAfI6FlWttISi3
TPsruOCbg04lM+AfTTTF9FsdE08jmyMSCpCKBtGJ2TSk7S0TKCHqNQyVP6CMjGy8dXdO00DbsSIJ
8bmGWkfq1r0wgc7wV/91CBL68+Nn5FZqTgmL/IcSil8+QjNT9wmTGVWniBO4qYYYbOTPwt3gFEgh
nru1VRDyVtuUj9LnlETwSjy5IKoDumvUsmye+RFHG432Rsg674iF+6Z+RbNHkAJxDNdj6JxtpOAR
2PA596TkAm6vbkoUtx0NvXU1iLK0LTJHF+1HYuCubLrDpyx9k9iOAs8oHOdPU7YutwqyQm+cMHGp
iNyDmJASbkQ+e/wIhT9co4KNrGkZEjRwGj3mxipv7eCKk7okZ5cY9NwUQJsWtLDurYDH9W6ae6PH
4yZLEjn/ntJPuYL0au9ofz5SzWHKumtl73IK6lSUuo/LVvdIAhsgSWwrvtNG4EBbNbI8wdKFENpy
78YKr9K8nWPV4YZOnhEItumHsjxyUBOPRm54ms1cFzmRm+Wtdk6QF2JtgloSuheEaJuTg514IBiy
xPzDUEqkLJDl90rYszZWdnSdnReMYcz9C1jXjYG3CSJe38Ohyk9NVCxtuhbexFzIUIycVCi6JIAb
VdmnKFwBGdHyE54XdD8VhX4TTNSgz8pK4ntUwUyznaa0dvBn8ZikC61k2CVYH1t7r/xQh2nrtDP7
wUQaIbl0rGbFSevarlMvrUkJjfi1kj7XEDlfojqnHmLEkS/Xahr5+g07HhQd/5mMN1PjvWugg2bY
6BuKCiOJ/3pgmi0LrctyhlHwpSDPX3v3Fc036LlqaCLJor8mVVC2Jcr64bZlur4K+QuoTiFB/bPH
D3mvq3PKaSa4xwH4b2V2NxngezVLsVyab4+BTR8kpFPnIlLP1ek+/Hga3pQ6fiClpZY489bypN+6
Y/+DL5muTuhI36BGhjvJTNPpNrij41b5/+2q3SLMi6amVlpfC7uWdho+TbAuZAtI8Clqozx/P2Hh
GzW5wJ6bdbgbfE8Ro/q+lZHJRetLl5gXHJNNAx0ICexOBfcbGbt8K7RTIxGF+kgqXwc1zpo2Z/1Z
jbqiKQx36yitPGekNJhWVxgITGpk8OGWbgJ7UinC3LlafBVYy4jR27s4t1oZeFK6uym0++vHR/nM
pE3/VsNPhjhJRCFfxtTwgoaM9Vr+B5dXEp0fZcPN5hIYuJNA3KJGC/oPZ58qxloqFSaqq5t8U4wu
+pnpG4MlZzn47El7g0HB5pw/uz5LxyZme9RLhv0Sz29PWTKVfGURHnt9Kj3J5rLVcrlVzLf4wEIg
UAFOvy4NMYOenYd5SKF8ZDvKfFkOEXod1hrPQPjAd/yp5XF9YhYObjckjzdoySk8nVNb8kwr9w2C
fK+JyPPRG/sL+9CrAekeX2acjPZptdOi7w4vpCuq4t339LLhU/Puc52DvyI/hUI8IRrgGA3GSivF
x869OLmGPw2qIJ3tOrBWBZOeZQY3gQRDrOgEv+rkYQf61zTCl8/qd480bneUH557tMvo31SerUT4
2rwoz2n619I5RBelVScLu0JzdfMB2tJjdJgq+UFAbAgEAORaU34CiE0ZXfvuj6ahIC75vycV6eFD
m4PIiw+wE6a9Mbw7IEmyGD96Kco96aCYB3+sKth7JReXSyEWdJ3EfnDsjkJVAPZBlonUeJflxMB9
8KbZa24QTMlJD+5JFGI5wFon+RpjgvSo1iQvf7Ro4x5/zPlJshia7yLwdnP/l5rxiPi7kir56ls4
2TsoPXtrfA8N0Bj/zTvTtUXBtz4ytTcUGxrocLLyi6SwpkwXzZJyGO65V0E7cb87h0uu7lmewNMI
rfyVx4IbB8iw5stCxJ5p06+bXTvPRw9sQ3hgb1wtJdF74FyxLZjrXWj3sZZKqPw1RUeu5/obn+d6
Ip5mfheKHT7inNkeWjKmozCf9kwTjIdAby/dU0rAyoor3B5D8HHMrxgJXlts5vDXG4DYaFh1L9U4
4qpzcviCNGLbDLIpW78w/bJYs2LmpyBx+Fm6wJq/Ru6Hmiq9xydLqyDyv1IIB5ODrUa4jhLdxZxT
yfVoJfYny+6mCxLgIddF7MlSSGX/mdGZFHVMIHnWmLGAZ5ZJdB62P4C/U2Z0KtCxogxa0wM/LVmv
HZGLijNxY4GhjINYZ3jQBOsCVg474hoL8d+z5/jWc7Zsj9V3j1zJEIkSWHMrREKd51Y4VDV2OyH0
aqC8HaAKGdfSJSXGQLY17Z2/hFPKyP8+y6v2qu2rwdwizpkKDDbJ0yVpFxEJeskilymZTfdN/BDC
vTAbjHbatAj0pGu7qicLwPHuUH8dFtisdYGy0wuwP1CqSOKJidBshjqeNoO9cwDDudUXIYDeuObd
SLmrnnv5EkuJrPEJ4TLz2atX2CV7yoy+urPShMdkEr3KUla6AaceqFVjM0+BM2l5fYghcix+rokj
IacBt+HOZRgOsl97S0qfPn0xvWauWoBQe3eaSB48XTp7pTSbgy5RV54+TpSbgk2pe6Lwhsndsc2d
2ceK72RQqSdYWGk8gxxzHKbcUL4tplMyctQyCEb4knqMCuSdbedwmUkTx2CMy8PKf/378dPIYc74
GnBZPu2S+fJtoafkZpTRUaqcLk9Gw1T1/6aS6yqzoT1Er5DYjSYQ4sMgHpkI5yxBJzYglfs9Hfvd
TrnriGpXt40tuYUfB876oPYD3v8frgofPZJrluO/64kVy0qZ0wEpxkwePVinwV53xw==
`protect end_protected

