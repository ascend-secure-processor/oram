

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Tjj6TThJhfnAmLo7oIpctlFOokCH0PCTpyCh1pd2bSt44jTEefon49/yKIQIZPVBZHWEuh4TEjbv
841vgrGnCQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kufniTMrhOaDqQGSHxUcd7FFMjL1wRIDnkpb8QfUlB59hKR3x+6ceYz8tnv96dHyLXFspGDkvIIS
AfwaxQP6j3w3Vcio37+at0g4uw71tc9A7fZiEx8sF+Xyta7rk498JKFI4e+x8HZZ8zh++OgLff9f
AuHQUfQitlS1ZStkATI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1ZIScumKuDClbm3sm8YNCVIS4ZQOld0dv7QQPRpx2m5DyPrmS62n3tn47TfwscpHHng1va7uCFlX
l9nAY4KueBz1Fdfybk7k1RA98NtnOBww6JSfDnxRwFTIapye6iIJhGmYJIoRf08A9Do6oRXN3j6H
Hx4uJB/P4B7pnakPcK81X4jBz4cuDoy3UITmltHpw6ia2DQYIlih4LJBoCjIebaQvsdTbldOecSc
toRo0BBTgM3O6jQwkDPhvkm/JpADE97PM4m3BAOGofAvrGPDAudsoFuW1K0C3JEyYkiSZOozX4Iw
DpsUl/eRnrBRUTXsARIKgSHO0WTZR/ndkMVaHw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dZ19IXXhI3is5aX2SXvhu2pkId41bH1ZKB2mCtanVGF9GIYicpFKax+2oPDRel7xvvMLSYRq7nUU
Zqr4PQ56Es//zDT7yE6RPGIthXyVmqDHilTX2HfdgY9vPAQd1WtE6yzbSsvj1hHspLezpfBlrMQS
RahD9vWJzCgwZDhLxfU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JdJxda/MKKcBnKRi7UZe28jwxgzwMwsrzF2g5IIEMpCUXAu9fMvMJPdopsJ6n6cKwMa0ZJYXaU24
wKuQhfg48jir7QZjNc6bNHqEbWwmQlmTfAqWUEg9694i3R7Lzj3PzGEh7Vmc2xkMSAA7tRrCTr4M
Twbu6MuwQT3FkrKtAdlpAC/fx9Ycl7tICcnB7BoCGKkJdxUKzvq5mNEhaw+Ob8xn+LoZJfOGPM9e
FTonoBaGL2AOvAGGYTU1BNV0vrhGXUcgi/3XhkOrwwv+eTeFF3GRQPTYw0rbYd/1sJgZ5VzfAoSQ
0oxeNBdBZuDfM1zMPBiZkBwn1yg9nYSxyOOHGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4864)
`protect data_block
LKZvEpr13NqKpuQ3z5e36UV+M3ItoXGaoUgooP0vmfG0IotrumNvi9NuJffuIsNl6qxsU2gLjcOR
k7fMRG7lDZ9MHEyQ3siOq99+tGXl1NmsufpF+4TyAcNxkNAu7TfhLNM9Bhznp7iUF9drcqCB6pG6
cttijkpGY36zwu+ujqmButC7vo+vexjQKZ5Vo79NcUL95nYPRJZOYkfwRyEeLkzY0XImil52VSqe
GX7/ggxH9rQmC+rlpjrApYZUZX1lCMLTVId5o+HBsCT1AQmNYIv3VeIi+f2S2mKlDw6iFdzCc7cy
aHC6ra7nsit9tTARiYr4fIr1Wb2JpbInpUsl6APu8qG1I7W+lFWPkDd/L4us+az7NnuwSBd//DlS
MLwft3PmVMIjWk+l3iuY7QjkipsfnTuQPtT4ex1/MU7UqlTQ+/talBTQ+eobaFTZ2mldke4szHwC
/Tul9WWFRblR2U394ZyH4I64pyTvvoQRuAvySPRm1uJM2r1Zc5VaF9N0G4rFBOcWP1CW3+64usQi
vVgAxxPN6MyYDICbhirrccaNfxOCMaUe/vNZIsWL6HKtnOfcfzfhFOBD1leuck/EEelulf+GpUwv
4tkzfGlCpn0gBHzrd6DNdEWqbZgMq99gXXSYYvkXGZ8onz7Cbnh8i7iZN+jjSQfmzcTFedDMkGA+
myMDWtmqAi23Qfjo1aHnAjGwqsWPJN/eKWJNkNrj3tsTzaNtxxlVK4S6fx1P925K+nqVSHFK6/CF
Galf0AU9cRLUiXgAZsKSiBQ7DIx7yOXBVeq3RW0hSBMADsGcE2fxKTzPQOvp+gt1prsjt6jQx0fE
IdhbhmqsY37WrrS/aPw5Jy8kOg3YlFcq+AbpVvoC6V0KIVfDAWWMGihMz1XWzgLTYy6lh2ELxrW9
YakkwZzonz/3uJ5FKl7eipwjNZ/N5c1HjEsK8ufTEsA+TLQwQ1X26AKJfFZaxHna1wNr0vkEErcY
gOWfT79fx1g/VTnjKVxxUPLop/EJ3FqFI2ShEcAEQ+kRI8/KpuMB3kxCEyTb61cN0xYOKbwV6/VJ
S1x+tbd8QR/iKqksPBbqWweTBv00m/BJNrQP0mF5sFTiLLDTAsVFNKA7g4WB4ETdUG1hy/H4NoaW
GY6DCDb2HY8yEwWaiiBen+TsPtc5ikLlEX5iHO1F5RoQRl0lRoGwA0oRLw0VZv7w2mxohn7vMhQw
fMv0dN0b259b/VI/nsaU9KaukFJRNvNsECxCj9XKRkGPF4Te+fT5yEJRJXP948Z9ZVqpJ2TkcCYq
XLB4BErzrEzeevzZzb6an8i/i3NH1dLu8I5ahZ61VYOMs15bjJCzcDiWw3X8JTZGiYjvO9c7QB34
Zob7p0+fadnbsagpovRLS8t9QuDyMXFJsJDXJIQpkOcPy4rlHPzIN4znaXw0jaO9rN5zmg+22vWK
aClE2nrMYFKUSCYCgV3JPmoiHLaibsiciB3xHPb80AEeIjw/6uaYjZcSCuR2vMp2TRNQtU6Xivxq
Om74Eo+YwAPnGc/AOAQk6BatDaK17/ZInaGziAOd6DIrrU+KEfkLXHWhYER1L8j+wFmE1jzi8DfT
c5eEbM9MdY6SINX4n9BAszqI+Ia6qIpmcd1kk3kDubQKC12Fc7Wb5hUVejICF8L7E0zTJLkrDbNI
X/UcjwjMVHeMit3WPdXthRvT/xRLOS+Gv/uzbtNXI+4KipkgKA+EVSQYITT7s/kPVdFj9KA/LbAt
/LhROeW7iQyUki7oH9DNT799fnf2Ed2CNXftTYghHKlLbY1o2odKjPTs8PQWwJlAr3zA01pMXQbB
kCNJnahz9mL9lcTewSAsT/F7FYCRjHdhFI7zubTCzl0VKKIpgzRWHHtT5vcZgraOV5iK5zYUv6xB
zXR3Q7YVzu6Q/j15Icv6KCdz9Ex9cv1O5PyM7S78z77x8fq1XiKN0KRWcGx5hsYHpoLIHuzJ/QTY
c1jwPFdwG0cAquFOEmKovgQWGTvaYPy4HrTy2RWt92nXjD+UKa+e1/MAXn6idGezlSVQbmBeuDlj
KR0fAc1ruipLAw8n7iQ8vtf/+lc280Vx6K69bwYZSh4cco4VN4EMwRDKPgbZSKfu5LHxIzA0K1zs
OcGmxMUI2LznHnmj8MTJPA/h7yEcv20k/ajJprLU6c5era4xL4ChGjHVFiCT7X+A35YNFsB7Sjwz
pwVNAzH6EvjgfhRfKeHZ8Yx+JZkQP4RXT0lrxxitjZnrHLHCB5pvAEWT9/50hRzJy0FN83JSHbSF
CkAQFfhfdd+N8t25QwlO3zG3vwjvVrs8PPBTOKF+r7x2kLtK88G3s1TIaaF/KVMWkPWXZ49fSJqZ
Y2KwjgyRaNp4ko6vMCjmMv4l4ey9WHS8bNrPm943iAdViTHADg54QkV1SlqlA7to/aB0iAScaexr
sK7QvSkIyODp9pP4oviVh4PcY9tSK4sRD4lYtEb5zdKqZp5fde4OB/rjcUXX2NRKv/2f7MQjy85r
FDLE4ISlLMQgi1ELaWcUU1PPkBiYE/HEV/gjb70FLume0Hgr4zfdaxVSMoZYy1cn+Q4RrFtlbi32
PWK7vcJRb921Q864SwhUM21gULPf4Kmp5vXWyKv/hqAGknh/JNVAWjCl9jF+OoEEItlyRgYQTdZk
KvudilBFKYIldz4FROUPPodC+w7qgXlFRxEP+Ba0MtBgtSUHniHLjMDYxE75pz+OEDOlG/AP2jip
A8oK7RzFI3+n5vVWlcYfS2Ai4KbYkEWU1KG6BBZUMOtKo7/P3INlXVTHCT0QTzlL2gKm/QozgBE8
Yuq5LP9i0Q0zNS7vGRrf7/UK65LOFhFkPYp72eGP3uEXvTjzcTb3BvH9vR9XehVW84urLhHjXsm+
EB8wz8bI475ObHwkGITq7h44hglQ137rr0BOP29mk7lprxjCnClHNXJgVErq8A8XZv9nzFQ/n8KM
J4n1kSnaVNW3JREQpM7qwMaOpyuTApwGCsz9CdGzrlD8g9vJPdaAKjngcbPugReVM74+XT7Y501W
X6mglMUNjIWS0XuiktZlKU6p7eAwcuMlf+Xum6yLCc9YxsyegroZGknddmuGylc3RGCjWQFx91zz
sJSPxmfuaTggPpN5Dj4LtAUe3/u4A18WLWECVOcyPAG4RmzV/q8lc5y00tTs5as9xQ5nIEfmx/Ws
hqa/F25VjbW27IwZoTrBipclUIb52WCqlu2ZG3wRz7vMWkTGat8kPDCdMU9BEwnu7T18OeM6J2uH
j9S3fjvtwJOvPGvEfr82YjOY7NclewRWfbTaQngD9btQbFs5m+edaaoQHfWxxMJda0SCNF0fiEYw
GbkgOkJ8fpS+CjocNgmEoe7YmENgVp9CabCmd8ZLZeYdvKGt0JlGrtND/fjM/GiIxg0Z6GzekCFl
5dM9Ya9aaMZqAE8sjfZr85UtDeWfZ7m5AcTeo1ZFdjWnM/iqvzinqVd05QaZeTp5rOrT9RN4mr7p
ydiRIIs1Fo/0Wts4d1XSKuGzqAW7oRvptCemJDPilPpxEwpZqSYObo9sX9PbXIkga7buhIQTpKKY
gApZVS5XAQWyCmcA05ybyti27ymAZZh++aT5+qHNV5Sqde81fTBv5uOAe7yZIdjP0b+ZYZzY0AM8
sg9OnnssaCgYVD+8PQz79DBEwAinaXRtxxrdi0t67SsQ0sItS5Kkfs16L98nKfLZcwxa+QSzmRL8
y3E15J0X1QV0ySKGMm89VdgXiMSI58qzHEWQpp0HvxIX+Gmr3VxPTpROysO7O9w+eeu4OUR64t8/
YXl5ucoDjneP3R5xq3HLukDmPbU2oV0eRYWV7pPsRwLGZ/M9aM4bc0ctPouKv1DS+xwwNvIzHbM8
NiZLa9D/gEgMmLsjs/Hd73gMWUtyS9TSQjVLggvncZJ5u0gTJTbIOkqfkcClZqPQhuHKBpK7FNhg
w9jEhCfyb4ZUJI/sXZKBO+SsZzSuD6BoaF0YU+bi8/upsIlSptxm2oGW6gTp2eCBXqL98zBkIdHT
Am9Hwf4ea43lWHZm8Av6G8O5/UalVurQxWamhrOpBkNSgszXUlL8B2EEuE5VD6ll0jK+Q3Ix9Qe0
aG7Z0OQ5SM2NpkurBE9XSoBiFtpvPdJ6ZIBkkmAsfKV3dZTIxKaB2pQOT7HJZDWP5xiKGCpqqL+w
vitAaDp8MIqAd0bZgMMx1nA7KYRSQPlGs4fcAPzhF3fAhq5WMQgKTZgmJl6yT4n6a11snar1xPYA
/cRXwvVzxLyCnUrGn6lRWcVsDyDnMIqLimJXsUujxz2wTsPt70C8DyuY4l2iFG4Mm39MSrZX61e8
gELR0NyS6qtRU1dxvElO9I0gohFyc8xN3s4ogCeBuFwU1vcFSRL4r97S/OvoMwUarZb46JYqZsAJ
Wf4Kj7N50QJnpc3sSLz48SSylyeyahRHCNEQdXoi3vPISfewzxhs8h3czFnwVGpmP2H3ZBoVismn
vR93GEEWyyzA1ZsSQt/G13rBzec1E1uY4YhanXvbQqiufBtMytvk/W7zKN1HlRzm3dwWgtMPJaBX
w6PHZeLN86O9jmTl+seVKnFzZNpzto4IE5O1k3grbKXDzcUTDlxZ1ot0aQa4WYXsqjO/ebIy77zX
mEded6dNLqWEk+vqEkhVGcDwmzpxL76jPmcJZuPeWjBFnwHjxyZGwiJWKEFJXAaXjkkdcZ0sLaJM
ctNOLbdi1ghl88ahrp/8gLoamVghWovz9VF81moq2H7lyrwIf8pX/mxIbEurQVUQWf7Gx2woKYfX
d+RgCNI8YAJu/cUFMG+nchJlchDYF+qah3aytEhTjxvel3R/8SygViG0/Fw8FBhA3AntCBOSYnc7
WLRRqISB3p47jvDEpNIvbxJ7xYgT4oo/5GlqwGjidBUDzSs+mR2GCUPlZqyRcIxuYP/0X3tkRVlZ
JvyZO0HxD+PhYef6ylKfyTuGovmm8OjIraAwGCCK9P5mlsvqaPv2dAVa9Rc1S+NxU0s1qrvsyEuk
dCMZgHgtJKHJCba6ahJ0r88DeoKHePzM9rEJKbe3jlftF4enKYOZNnjhp9QxHWPpeKvvtoGnDx/+
GorWkHt2pszivm4/ilDIhUVT30BxN07L5aI+S27vEHtQYmQ/9kuHK+Xk06622USQ8nJ25TYSuqrt
vSZoH+c0GH5OLTKbcUWOGSHG175b9Bw5WGNn/feJCUWmwvLe6VGUGPsk8U/c6dj56y5vD7BWXcHI
QWVcb7i/8vvNrYKwIoqK7F0pJp20qrM6DKl8hMLgI1Ve3aOlN0NNpW8kWHNPKufuWCjH11INXtcp
EbF9e+s8qZ+rvWZZfb1cOFa26gAW/TAoKtN2Sn05/djA+57kD8NBQB9TlVDd5CXe3PHKQRK/c5h8
iqRla9BtJszaaNbP6QvNM9hJAAVN1AM9F3VFFESrPICxKoHX2HQ7r6QJA+htOxiIp2WllAtF4yHh
aqGBj6zc8krMLrfS697gyzjMyN98u7Ep7X3EnoY1z5fPQoJ337RDy4CKg9yXdXMC2AewAVqjqJw9
gT1zk3s88r7tU4CRCfvxELjOTz8Ev01CqWqmm3Os1m/6sFN40VdxRYwL0H5Fskqh6LTX011c7RcV
RAg4TfttN++i/28nC+FJQ8h7H5VqdpgPIh6sDOtRWvj1GtDv6pDgQVTaHnfZhO5jbs3PENKb50VU
yZ6ZfhtXhwgr+cK1Kh/KjKSuspBIue8DNb5TMkDxXffgKKA5f6EXX8rjNyyOWJk7LDQMXS/rstyB
wGm9zKBGvlcYE7aiADaBvDhbqD4ucZXYWjJ1e6ZaopbIKEtJNk9KnOPs+reUlZITZhY4pS6ysFqK
6QZNzrOkbDkjoNDDsDnyi6pw4RuPDp8vZZ6BpqVp8koy8Deq5ogIWEDv4mQlFBJAlzgVMsOLbW+U
GLDRXb4mPZY9bXgUC+2Bu3+Ai8c/n0J5YIB9jdbfCWNTm4oGAJ3ziVyh4hYkbyO3andOG+k2J9n/
PlJugCOr/ZhZea8EogGS/DJ3UgcBhKd7bIf7MD5F6Lp4Z2r35VxweF+AsYHsCqB9n81BIadeiLED
Ht9Txg7FZYi1atXTiNaUkIOUnGbF/53ZsNfudpYBQ2nduh/bBQGWi61UoyyXh4raktl8GIREUIWB
ns7ki7jdPy1KqqGSUzM/QAHZsg8SNWMWsIaNppTc00QfiHaqVdT7exeWK7WP3suo+JbKwpyKXuC8
R1MYNpbxnee6wI47EHOV4kUGuVToLE1ZUfJ3rvZohenzJUuW4wfPYHjoRFtcOFaEJA2+s7HEoyh/
8mu28uDt4OdM2UBz7gwW313Gp567YF+wEW7idUj+2YtzkGubGsr+1vyYEA33HeWJ/RP2li9k7zsr
yEQqpq5LsFxAuHYX/FNcGZNIMzOvt9opBZB6AJVSrlL4RCRijPLKaCccFFMzmnU8mUc8za3800Dp
jDd2rXwQKf43i0rXhVpndDEImw==
`protect end_protected

