

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hGnkkojJvcH1Btj0aUpDo1AIagcgLc169BhKXOjPfO0e/Un8ncHUolQbIqm7kaik58sXeBllf3lh
A2a42qn97A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5fCTsB5sZfjISFw8+J9F1wKLotE/U74z0rVWldcsjDTojqzmeWf6i1r2wgMEoteWJkc6gwDpeVs
zqQVZ1EnBW5MhjC4hcu7RhtiBy/Tdw/A8lKY8AZVu0Y3hqeCyfa04I47rTwTO3g1BZjz8fnXeQzd
RdmokBrUFn4VcDoBGh8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mG0xGJVeC7nZNIL1mQJkGv0IEzBiJyNidVRWf5c++63vQzVYifsRi8KWu66x8SDyb8zkue8ntne3
T1IrvAh2Ax724Imgcu0fs4oXDXy3REBHlcHm0C7nZdo+DeZmS+VesZbbWHsXySFVntEkuqg08l9I
t3wSZHSldkbVH2CPDDAmQc2FlL8PGrvRBt/OktNWcnfXmZTKsv87o603IpGTrqLUnKU+LG7qZtd7
bVvKHo8LgJ1U3ELMAjxbtA+qn9/tQaI5QQKkiIZTub8ZJNAw1jRTpDJLOtfiuYsffNBmHPT2lqVV
7osZJy37XQWwyGJltPsUWK+ck/poSMGbFthA9A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yO+6+zEb19gn65ome2eJWY+JbpbkecSkyQK4ehpLO6MOjholoP0Pi8dASPnjw5daPnA9UTfGNfAV
ZSG4BUMXnyzg5ZgnHbLvO80NLAYMy7i00O6VNKujCHqoXoWBbafcB1zs1/KBtkXQ+aHmafkKVxue
IbybEEMAHF5RtAiHXi8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bvel4swTvMrzbyxVKyLjgcZYRrbYYeRAdmC6QvYCS5vLiEM9sgXEQR5md9SC/ueLG9lO5mXbVdcL
vhUhkk8TT7YzLalBRvPazAm35ipXLREsJm0G74uBzDOAGJaSm7yJ5zZFQzKC3mwreUKMSYiR16Kz
bo9Kw2jVHqnosMZ3PsdNaNNH9PhwE1Bn9bdQKPtOUGo2BDOw87SY7jkGx5HNa2DQaKft7fyRKbsa
w46nROl1tlCPVaBwrGTFnGoyRc6feQPKnxGxsE/kwCAEun2QfOJl/fUSOvHKFVk8p4t9E1hde7Dw
n191okedGliv7eBO2FWPrUbhwHn7tnH91e34zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13104)
`protect data_block
ysOqb0sQtHIppjkksf8yKyhnN5AM8Roi54RY9fxjFRXnWl5r7mXs/HmMtu1VrGeVchFRSKUuEKww
8j1WBaunKEvQLTLx694kf+8iXklMJGftr2kZ8JBefXt8NECecWK3EPCQUaNuhuUuI7W9ScbayWqv
lAMhZe1CDppgrPlDCP03GohOQWl80qMLA0Zuteql3HP1DPqdifu45QqOPs7CUoetz8npK5HvyZKW
K8XFY7K2FcuQ/ecTJsZsMLNLW+6gAuk19tdBGqgN/IG6mmX48ipBfgD/9Pc9x7Mya+SMFySAQRnY
wUvGsVwQdHKrmN5wiD3NgnU3oeTLldUmb/An4nltDx+ra3N8wLCSTEcDqlWjaI7SdAFLt91dtwhN
Si5OOy21gy/3pGlvYJGJyOyAbIxc3rl3yfvwkL36PzrvG29rlGH63IIYH/BnqNZUgvl4BezvziWj
Bm3IVgvWsO+p4/oucY4Lf6Kr9PnYQjSpZsSaU85alQ5xLYvzGFiN9j5GQGyYxk4yNoxUMIvRAE0w
J3Fr1yS4a0tprY6vqOQc91Y+195SbDA2sFlEEtu4ZDk0HGhbGZEQ32XoDFza3Yveaw6pHwX59O/M
x+RbjNz+UwKqp3mebXlpxe/ZXENw+MQHlH8/WPMmm/iBAosLVPL2uh8YpD71iCcVKHCTGzr025XL
ebQ1X6ycPvNSXi5KXsI4hrc9lV341b12d9vdvWRX5iZ2+sz83E4vmk0INgdylGy8PKBqtBF5hYWz
Y4kSrId/B5NYWwPm66wRX5koZGuCaQtD5AGUCxaEWPBoCQMLy6xzArAAH0f2IUuGySrz7aPASWUE
4jM6YTVEcPvQk/NAv+o3wL7SnGJM+vbKN9J3O7O1dDSBssudWydmQlPkgOIX/SHee3ujMlqW/2HW
ECERQgNvQmaGl+8wMxmgG5k4GHIedJxGbX5o8R/eEeG6Co4rQfnQ9JgnUEhgwWbCsLN8HIFtmdUH
NnEYqfUDWXING+E130kLfasCVmRUhEP1OlkQLG73uF4Gj8HQAQHHrm61NpHwWfEWgut96hff5oVW
fQKIkMQEOJyto55gOUvUfI+IQlGTUyfmrXaaXmh3+uY0iYg8VOnbwO+Ue71PFBV9/puwOlyH1H3Z
BgWWNKPjUcmY4JyLiltRsJ9G8lu3ucxGgmpMFeaOSjjPFbC2yXvgM5a/Wo2mP0HyEaBh0k/kJ1bb
7X6okd3SH55MNpasCVXLDPltlTHOlAMVIQpbSaW9ypuzHKMUa9tEhqeosQgbH8KwUDpnE6UsKk6y
9t+KFa8mj1eu3d1M6C+tc35cg7lk9Dy1bZOWbgKuFiiHEwP6jqtlp037p5xy07vqYNNtUCrM/K/g
WFUna294wFz713itGSQbHT7MJYV21NPQRjkU/gENEqLj6Xpfg0qKox1PPWNLgb9dUQ/WZSeQvTE+
6Jy4mdoE8LnvjisSyMaxmMgj8CBes4lsUlEaRxvJ2gEC2O1Ho//TBStf51kMmdrtN4G9YEpxy9ou
xUbOEv1p13GdyOQOZg8WljksLD0rfAxgmKxjwpxLA4b9YQCaT9uOtPnQdqIUEsXREGoYA+VMTfiQ
D5MJ0Rm+KvNYnKRXgFw3r7/7SSyydKXfq3KHKc00iN9VcJhm0bCV7NCCzXFNCi+7fiUmrzMutNws
HTxOqU8dNGFn6d3bLbjPb4e1uqiylSxK5jxGG9GP5GBH5C0Fw8pOrFqrWuxwnKi7dmJ88mTKO0Q9
rkDMIke+6TJ+oqItDcmbjCjnao837GlJiXMlnyrTnW5waZTMMFtk/6VaJzXmwPEiF8OJpvXg5YL4
VLdSRWJh1o+wqqndyH5UFzfOsll93GYSJ5e28C5V60k1jnfenSEtt1YPTUbn5WgBdH/6cGXA1pbo
KUY5QjPaJU/wb9na/kpN8f7cMTEE4CPk81Ms0VqrvN2c43P+OnC8n8M7+56NkXQ8TDqHAgHNOwgc
x9VVMzDMMzLxb5V9UjnzTmWcqlxQGvGtNZrd83MFBwJ5sraPgC8GAkqSvX5vDs0fkraWIR0jaiu6
x0FLiWp1YOndBx0Tq8nbJBfnH13GRO1UvSP0sySSVU1TDPXzRc26GY22GJVh+W6ZwTqXq1Kfd5QB
QK7MKzIrQNd3nj++/ktoLCkdhP4rZxCAka1Gm5LpGZu/K29hxnoB7W9mLJmz7/ZaWkp4VeqA9SA3
JIYk2Hr3i3R3EveO6AHOpbsgc05LwZu2Kf7mTzh3LErVtpnaiTMkaGqrjewGf1fW/SQt6Fhe3LNy
pr1iMpYczlZQxY5TdmhfGBOlY3aDoBjr7V5gRLS8dXg8Tc/n3rvHYEwFoxZMmI2nQZkujg95kFyl
uCvDAZCeqGuJHWNFFePOs1Fo8e/Z+gtWci40u4g+j+w52NUM0eX3wI8jqcYx1hGVX2ynNcrdKJ+P
P9COc+KY06J0r687QWOWyEqHen9+697XuoaMi8PlMpOquFFQUBvkkeaBbAy3XE9qWuefvcOGbS01
dnipne1FQWjj8IUR60P+OKHcq4aLdGaixiDitZb/CQENRX7+bJ5MAxNINnetfjB/4gLAagnI2e+1
53iyS8zMWI6l3dFZhK12IPV78U5NKTEbwuuWqW6PQGDHXr8b6zS1GZpmzP69kjGN5/f0c5EqMmex
V4zvqXuCVLYRTNKpqetsTSRfQIY7SEvgD3Xxp+qy15kdXy8e4QwasYznBGYfrAHwX7s/A+qT337U
f9Zp1gTYzbTDzzJpfBXC8ygmmD//ZDpwQQs83Ufa27YQBIlgBRENgAKL6ChRFMWolxYWu5FRxZ3j
pmOQqjaY1jIuW/kxGMrTsz17eHecR41mV/QOY4GYSmGAx3ggVkjHRO7LNKPNXcNUQD+WY7NOxLpl
w+5nadecykwegs7RDenXfkXo6FIQzE996uZrQZ+tnmsViZ5Eallt89VTTpL1N1/6C8deWJr+eo4q
vfxqNXO0td9HD3EDR2DiMC8ALMQplntcVhV93QZNl3TAVhn4PcLZWaz7wFhOwTolG+SjL0iZ7lcN
exm6q3IwCUSZyBoedQyxcSPCPV7uoUvZaKX/7oh/Efz0p8Gj0Ha8jCieC+CX4j3dfa9H8VyBdXOC
cuVCuOrj7VoaGSniUj8XHPasmPr8fCiw+2VGstXIc/sTcVIeQ/ddIDf3rZZV1vduHuRoqDgwuleG
6O34Mdukz1sCTl/BKIz8t2/x1Wxs29O/ofLyId4N+gzrXxnndY98HA2Ohi3pRn3Ly7oYPoU3SB/d
ZZByCoRUYHs5Lg/f2hUIy8nCRZOTz4U0KBs7MygWWLfFgywr+wLBjLmHVM0FIHuTYDEsInoNM1pI
VKIYXMN2ShGxj0lWPc6Ki8xOkkCi3rxJQmmqtqsspM639IBRTnyLJQuyh+zGHJ5q5qqiaVYwN4pP
7pOgPO3fm3vBwUc0igvgLN6ttdLllMC1XpzlWlQ/8XWvpU8sU+ce7HtEDtI75iNJgEy+ZnFAqN1l
U0qmm+rUPWr5h9+rIFEeD6qxwK1AbZFm1X1ea91CwiLUZz8or4MoG/QWL++bt66/eVwUntT2GZd9
GB2g2KM8U2kQz7UtvqMNOieZaFxf2VseRK2g2a10GBJ9l71iYcBifJr0p37ouSLGJVXvhPKrjedD
XAjYKkkxUgoycbsAgnA8CcFXbmoe/b/oD9bgUA/MwUu8MpPkYI/a9s7I8qNgCl1Evx7guda3jzSg
8D7qMEYiUthi0DUkIxPuCzMpehtQX8pvmBMZ3w7IidtOMv9Ot8XBVHkCTElxDpaOhZKeNFDKGIHW
5HaqiSuAlZ2QBTGk6h+gNm8kcPBWd+9GHeG8y7Foe83ygyJNgadCPejYcBU0qzHvo3S4Q+Xah6kF
E+EqkXGxjoxcvGzFs8T1aUlO5oumMuJ3jKI6OlZQxP/0jP6BL1gijr90vVNwuNfe/yfyBgdz9Fqj
sESOyyowMVIaRK5SIaE74rICARoiOOwSQxtKv2LcmRvvUoP7ly2R5EWI55940udWhxToU7QzHEUl
IZjn8qNp5rDw7Ll/QlNRSVjF+TBbe9bBgJKR5lTeIrI0BKvz6k4v66N99wf+u6pee1414Y1m+M2Q
YrTOmXnmQeBvwmti7DgautRzucDUzsg6Y8FRPJ7n2B4vWNhRqiGqbHv1ur/m3BFOMAy8m+apWw1V
OcPhLBHizl+jK2DZ9brRK+KYLUqfU3fKJm2eUWxWwYtWYJnjEY0jJD4eT6dBEZ8x0e+b7sUWNn9+
GGhNzoNHjtgRAIVs35yUuYA/95le0JahHDmq/IB07mtUPotUNLLBqCqEvBFHKBeMHFIw/gv+xbbq
Dzz9JrytzNbw09tjLVMP0dK+34hOD2sAaryWIC7LCHyfOru7TpP2BZj5XHTEE13sWYp5f3O7597a
u6jUmF/aw2Zw2cqRgE55pNcv3rklr+e2Ve7Q9kBMkLFlCS/CyCYXE9uVXg2mp1EySwdowqyu6m3l
0jgUeqaeTtqFdfNTyitxeElryG37W1T089Rn2onADGF5EWfDnXEpYcdWBATWDMJ2CuXNQVUNtE5h
O0ss/px4i9CWp2R2J6hf2YxrJ5dkyOHRzJvBJP2v+5rYMPd4wwkdt2P8mhAr96VOhsKHo9Jn8rCt
dTaM3Uhxu8/LmqvKtADoKnMme6AT9YsL7bUpiV4y6a3V5u6Z7UzPBvjus/LmdMw/AmQXI/hfAzDx
1MYT5MFBZWH5p32lo/UO64RZA73jlZc8oRsHVtWMbyCw61aJRg9Y3KAqyDxvdBsA6m24n21e3jdI
RBgp8vYXs9WyyZEPWCy+ULo7+2Kzg6CYaEcTml+I6Z2QwD+3JgyA7cxhwJdT9SLhz1oiijeHnGH1
TnXzSWQKpLC9bSwDW9DHIv9CoEoaE5cbNxOo7YkQRcyFZzG1QByL6HuzqjbVT1PPt+10s/1qh1Oh
C5Zd8dj1Ksu8v4DJzerqC2w5hlO7n3X88kwE6V2REpk0finuqXsjBPozV8hxg8SwwEcpqx5kKEYP
mwkE+OcA+fst03Dg0cW0k1u9qjcSQF0GROk+JSj3HdB33dDgHSe1QO4ASd9be2hIYjFAn85/QYv4
JPbQc08ELAO5CSNXunCvvj+2HT3/UcnL/Wv6pQyuMox9Fxln9kO0lG3ISnEzUU6YgxSYmbeHm4RN
cV91YyvKk+ROrZdGRqr+7n2PAmwkXeR4JD73VQeCLOI55SmH4y6kGlJ+D77jweBUaoisz4HzrECi
Zi92tXP6oOP4nMfI3nt1kMVmY93q0FNGthYD+yPyfGkDGypeguPwHSFfqlrZ+yekK0GIB4FvGEZW
4oBHUDddPsz/xcNRjSf/Vfrc9SZ1hZ1W3uamG95VtULe43WWGXpqQbM3xb/ofaxJpcRSQOPNgeS/
cauvjXJMTft2TGSzP7iINOCXSSF2h+l3jHJS95emGeY53ScoULU0XS3EYqdM5KZ1M/oNPLaJfDjB
75ZJkIj7UifAfgyD0Z+N/hkfC8XLETMw5SYBDHniOBsMd2DAWwhnYCzKWRYpOntMRUgkST1vF3FR
6SdpfPRxb0BgYcJfwLCsmu5+EE/sA0pctltfNHKEV4JgA9uzhZ2Yj35eO9ZuXASzcO6H0uLZvHKP
LFkl6XuX/oci7YdvqFLZOEXI0Kx2xFS/ppsGMrybgvid2j18nwxoVTfK3owOAYrjOL0H4LSgYOEt
DsZqCYcGh+JgDHSeJL0s40Fg/grpzwj8sRS44V4N3ZJpRpUQEiJvvkWgDlflk/+rHGP25UN86aOe
XxvpbTulZub9yfWFcutx8nDeLeHWFOhJHrbs3pj5me/NNIdVAJ/SvPO4dG9ipyjr4L2ivqu0qbCJ
tg5iRrwcW4gQoXwoEJ+9NZ0YBuX0pMkLhxbyRrzoMFTNuC42MTa4juTRI/dCKqjuZB6qFpm1O43T
j13CxZvColcssaA8YC1a7xmFe23JIiCAr+qdqLQM04WJ5tN2rV4i1uQhXH+9lCxwUY2tw9rNo69D
4D+uuqNYjzsVCFAFkm8LD9iDy/Dak1v0F84y3fkUo3xMG6tnx6+Om8carBcAU6FMMrESRIP4prz9
tZ1SaYoRQyjtqxrjQpaEmpbIdW5E1T6FA3iOzIDBlcQy1D3Zy+UYyJhgQh7/Pi99WevzvsmIVjIp
UkT8WRi+gzuMS5kURytJVOH6uhUNKVB0MiE65EXClPRdq0387rZV+8BMkKevTdqMiTR0F1so+R7f
DNVaicKa2oVfWIZbwfw8hRTQEpdZX3zBs6XZgwPF7FMHxuPGhkslgt9Mq5U92LG1ciW2Us8ATLBB
LknlcFWsqHHbIuET2BojL1xr1/XnPi9zBSF5PKA3H4Tn82noe+pXVIcr9+hEwbWEhVS9jdp5hOJ4
y85XjNrvIl7eOQ1ktBxq+Z7MxpHetfvtLrc/vBnweruwTb9d0b0vWGJaWZgKTW34N50AR8UN8jZU
skOfl5mw940AXAV0HgfNxbcDmnBkw2qGU386f8sWGyFFmGvqt1E82fS6g9p0Fd3dc6jvF2BND0l4
/nc/fNiZVkExH8cGl0LtI3DtPpAUP1xdw81gKXSf77P9U52FBGrk3hBYROjxvtmkHfSBFS7M310g
K9gStSG6VJK/xAjXHNmpeURi4UuCAZgid8MiMplHvQyDJn4EMnpzd3Hmv5FDfavEeSu56Z3/rwha
48Owlnz8LZOKXq7DY9/oJMmm6id39iehfilmTpvDvfzvvplwER1K2WSaAKZgcvfGDYLdPogXNpFI
rycq5e8vCjZOYlQVSHZsyQ2639MOukwreyIFSFhwq4YADoxfJavOb+Kr2x0/4uccBDuJ7RV9nuy+
slUL52Qu1Ksh77SM8ywm0uIsZlrA5vk76yDCxwH61+3zqGfsEN5SqAIsHMtkN2fBG6I+L1UnOdz1
V5sTDGFJiu5Eet7Pixy7IG3hI3dzsM9WUu3samcNqjzLdI542xo4NoE1in6BpsUi4j5cLvyplpKh
+QIbb794GveSB2srfe+oigDAKzolfrI8airqd1+ODOJ9vjLUBMlZNj/M7ltRXbVIivP7FpyE92P9
EYRotWT8zKEg9WVC4l1mc2sOsW3E7a839hsCD20Cgu5vWzVNnqjIVys6ZYAZxbcRTtnEv6XrBNyj
skIY26f+/l164eXRMUlAMuO2kZaRT6dy/oeLvz3tS4UebK7Z3xKTlV6df8szljHcb+W3toOINnIX
+Zcbu4Kl1XPIjWk0ReWseZPATrldSrETOKb44axMdCnpldQNcVRW6+PnLWBHonPAmwEhNYFZpali
U0Ma+JDr6pZ32xH8XoFCM3zNWLHSBR6qL7FsYPxuVMy0iP04Jv+zXR0o76DSgIkfwneO4hkeV9LH
Kb+1NVjpR0exSSIe6wEpQFGYrCddv12xzY25EZUZd75lmhzG2ZMqkbE1NVfoL+RuuROLaAz1dGu7
mji33Ck7kqDN+lmqCiMdaOxug9byONmUZmGn+W+W+WR6W0BNrFUL3NGXW0QdpnrgYpTvBn/g5ePN
o8apKKq/eEHYCMnEr+sR4O5J8LNsiqLn+YRjCCLRaTY9memUNCYDXVnGh32iyWGBAJ3vtZE0cRbY
KVlP8F+CTdBUU+LKQBPNT/DhgcG26PKpHnOshb45Bbrr9nNsJxc0Wq6hfH2Bzd+MrQaZtiJsl104
TQZJKL9260soXmA4IHXaut1AhzEyWngYFt16vWcuv9PWKImqRfYodSLRtxRSHMiSsIZbrRwyVMeN
fDi4LiThJkXd6/oOT+HCHmbEqwT2iqg1LTN1aX5tPGe090jPpt1Yw1EL39a3jCqC63NM12SttFap
Hcaxe0BBW3v/NkZyhhuOFd+v3HznhyRxEZiSvqASrntnWZjtUfWI8Mo5GSK1rvzbBHswYsl1+fpS
6RsFjQy3Io0XVG4JQnWQOdryFf7eSpMG1kZgMaVwEHHfGTQD9hfCsPzw7s+umqpupI6FW+D7ck4S
pmcSvw7DFS2UkhpP/EZhfMBYB4mdITpaOEId3aM2XiSkR7m0xdEAerZwRDTgcPu4m6uvXddP0vSr
F5RFrPB93QJqIMNlVxwxJXwSAdUa+R4OwKsqdH/3eeiQqto9xIyBhhSS9tWramrZtm5VGxETFyKE
lNyiQSWrfuqa0SB5YJIfEE8TntylZPc7RVFiRLrwnqZfFxmobfKXe3GZvxl2IdOXW5qljPJS9LsX
jorGnwMqFNIemrk4UC9WWyys7XaCCq1rqjTfkoeP/NJRLUQHT6tkLoNlrOEuvICtMCKFKXu2BJKw
UdQxGQ1xguNf+vgAQcUuTyufQlNvYYWDt2qmdOA6/fwqjaio5vTWA4XFdPjHXgqgNS7croAo0V9G
5nGV+/MPeRMgGVZ3SWJIXMz28St6q8ZgA2HAs/648fBQrQPhmfZt3Hv5xmzw9iKhUvmptqHD4IIg
Kt7/svF9DFy2I8vPisD4JjNBDbUaIWAN37D8k4w9cx2+O0cTIsKTP0tblKSNz+4paCicw8XHYT9O
NjcNXid1XlofQf6okfSI0dwN3kl0DGdmPtWXJbG6OH/Ys7L1/D/eW2YM2d8A97sf8d6SBJ2sIyih
sotovtF98wsJNR8+kLT9iKVH9NJmuXutcpdo7RNo1saJkX6Z6jfJb7qrNKIIEo8ywTv3uIaDMVFW
d8ZQ8mLJMNeH/z/8aHl66bdudBPAyfhaPyUyZtS+ChdxNGqBsmw0/vG0CqJZzcZtcjZL8Bji1isk
0GpqKKnWm2+H3ZPFz1fwE8TOYaawElqDB9cc+sUcPx4ioVxrSGhXUZwT/OGlTdePRefwTS7RPSlk
4pnHQVGKY/o5F22cFj3K/AbeKevbYLYy6Q17++/Ig1UZwnkI8lN2oaodqJ7L4RyJpKIEV9u4cxSO
sNLfEbh/C3zyUp6R/phZ38GuaZ9pRd/6OgCqIBtsRMrPP/LexVnK7LYqyKS3kc6jkGUjiMR1qg7X
C2P1Eb/ybrWeEI+tv/GjNAhlfX1GCixvSWu0TDfvl1fM/+2CF7PhPhIJCFIL62XZvZtgS/ZizDIo
ju5lDhKXnxC9YSH6AH01wAGGk//k9jl73jo/R+6ZN/dbE5xZnq+fO+C4ZH0zMFgMYyK5LYeQUmt9
Z1xALE384n4rJr1V93UDzV7FVu92vTnv53oUzPHFu3evBFh1BkWR80JgEMlJbV+lUpy8GJ7IZed4
GG1p5xqqMo0zOCc+nD+FmroJwALha2AM2hTptWW7ZiQ0SXB+TiVwwdlCIz1I2xcTLLxjV/KrlUS9
HWau6ud3G4bK6WeLBb4rTgRUfjFBYAc3AXv/j9jqrzW0tUznM9slOm16oFMryHXByDqiMVJ/lb/H
umex0FYjN8LwC526sMoa6Y6nALWEelm0trKYhlE6/b1Sb0izDU4DzvTk96A8EPdVI05uwCnhhLWG
NTlTp+SkM2bPzVCqnKn7znvCsjgqJT+ElNKgR4UdbnSk7Dvm5v3KHITgMkEusWiRCD6861SGUnL5
e0p6qyhkiFEyP9yAVGG616EzFXlgKxwZKfJkA+lcPXWIooXR1YnB2mlLCZgJpwTKQYbhN5vqfrLl
/O6zFBiYy54FbC1PZA10+odLt7pbW4fOvABCsfHFy4nAAOqTbYeONJ3sbiZVpMWEx2gkeGXr5S38
SXw9ZK+mhSbq+GC6aCkILcigb3KALYclVM9ICsTQ44ccscJeY1LudLBDpwW6SoW+/31zFp+h/uhw
mMonXaYefCv8vMAbJGfn9h+qsuYEOXS2Qo63wunZPzxGoRpBSphDUPWc2gPRgUqHS51p2tzxjav3
23oXcA+R7tLnbC8bqXSneupn2SIEWjOZyop9ABk0D7Bsh9EyjdywNKZOO0RNAOghLFPNQndthRIW
Z3ukWo0cXSf9d6uphZt3yZ8nPN8lbWe+DHXWeTGLe5KODEvy4W78L5I2lwt9fPa99chSC7er3HVJ
5xYDjaK9NauCUaSzdNSqfJrVmUEbw6SWmaGGwbGQJ7Aa17Ow4rXE+6fbz874X0Gnfp0eLz7zMWtl
Za80OrqlnfXO21J/KW7fBlHvhY83O7Pp8TzitXJG9QS5bmvWWX903PoRt3dh7IpbEpB65o/T3rGV
VaFqLgy3yJgLnqwcdUV7hhAgjJImnXbnMih+BWmB5wyA18x4EenwwH6mFR8bC12i9VXk++iAg4vj
M9KzI3cDbnnMsqqYr5Ote1AM1+1lnf3h7A6EKS1J6SOt+oEO5jk1ZXbXMgoceCw7y7kMPFgd2e8/
SECWQwR0YUlrTe0Oer4Fud9Nn9P3PIXheb9VnML74xwOpOpXoB/yl7MQrZ6LFZBIldbN1LG/Bw22
cceE1nhMcxHnVK3Kb12+OBe8mx57TC5qDkucoJwTt8c6y0gWi8LD3dld7Xfyd+xui+5Xj0wEVBjl
VwqkAPzMOMyuhAMPdiqFDjLDjLFDlA4gpmZSs0p2waP9uP/ScWvSssRxTx/2IFqSUVa91yqyAPOj
lTPiDsE+9TMCBw/rAh9gmsoWG/YqeunqqB9mKC8CaNSSbFATPj3OqTs/6eOgba8daF3w66iIDqSW
8Ln2A3zeuZyy2oufj/4fEHRPWU2Zl7sTY770r6bYC2IcHoOauqqveIHbf11knv60b5KBpC8Z+bJL
tvHFa+p/jM+bH+qIvBV0P5KpvCgxc+EXo08c6doauJpKvi7g9qFFXqmAUxxnIVVCIxVQFv6JNCd0
C5IROQYnVGqY9IK5d5j4xhodcwKVX4oqwr+UmdjSNlHINKh+Z1CUj2DTLmY35EiNoceCGVffPe9q
BQh8RApF7rYB1LG4mhHJoG82RGfrlWcSCVZCSCm9v00+CIzArh2jdkU3dXlriM/kabbEUsy+tXFt
fynIbyDfcyal9ydDAAg3W9547aoceLSdFgs4e3nk8745n49ZyNNULVQcSgru+7JapqeAOop++RyF
MGIMgHfgqIPgCfnw/JNk1Zrx/0R7gqCqFDcakmM+ZWl3LaBA2HWufiJFeSBmTTvwoQLsfRYWAx0q
F26CclAnN4wA3IiNQwYRlm9AcmpwgrS5oC3TctpChO6r50Y8R3z/qi8tphzkHOEJZWEwxM86Nw2d
OuMVqdEVxIqnfZYdKq0tQ4oXd+0EunQijJ0YQii/8ePz1uKtVhEcUli9ReevX31coCgxB8YZKKgV
GDyac92e6vPA61VsUJNnI8GOzKb1WJwJkTFqjN97HiYZTGYGWgrxedO0XfQNwEKR64zRKsIZZnPj
QaM6FywhODURgJThVI25+HBBlLPhBRW3yd7ayJ7JZxI7VXtTtXmVGawwYsHulEZek5JrF6UxQqyL
TvCetT+HKumWWEnmS/RZDDbVWbCKM2DG8ByQpVV+SpK9oJG2JFZckFuGaNENfI+dre5u7QTaEM5C
qiF2+Z8RyDpibTty2USGmGnC44bN2DRveheCR5NXh8o3urMSbjkI/xCHxcaxHx5HakyVsEK5jC9o
+7oEgNhoO/SDISxtr79R4Rxrptn3UDeH3wwoV8cfI51DyK2ZIhqM08goPdfbR4iVtnlVBG6qZB+5
8G379Lxw/cR/vg3aDZhIOpqyfMoJUn/V6txulE7U6iDq8zIxQoRShcP/GZcp8q/oPVYrw7Mr4IEU
uyFCrl0n10rOErUq5BY5NqMfgdY9pq32BJFj9ICSLB3aUNiUEeS1F29qm/Gi2ljBBpdSMbj7USkJ
XnUBGiD31lsj2dZrWll0sKaQn/XXre7YBDVFvYwwnl5hRug355W9wbIrmEcJCUIPGUXkJK9W3E2g
0nk77ptnB08BCZx7RioOHpJPoytBOjFQ9xfxj63eoc8ulrpc1qeWFeB1G7plLjF2qboi60kODGB/
LXkpGmk9DcgTlIMHXoP5TZXTDjRWoA3SCtp2IDer7MA5ES8PBf1rzI4A09AchO4dzGjWwUkHZx/R
SWTRAWvLHYopn1sveguuYE9hTAQreWVDehQiieRQDJhqk4jOHvvmYbhOkou48oe3QtpkDIeJNn7z
9bJOLwcA1TheaFISpVu+3mSDsfi1h3d9ZlkiWk6yaOTGwFjad0J37rKenZQtwWEY+c1LrNgjSbVm
ADs7m9jecPtRREu1818NTbn8oEP0nY/aV3XAbCU6asxmJoUA1n/Q9gqgJ2RcC2MuJu18z3VDsUIJ
HRzaCQgzviTd2/P3FWetlxZW7U11LiKtUl/6ykmSHhz4bFO6JBf0aFYdWAfopQE1K7VmXEsCjXSu
zZUvWa3NprlFd5GJzy1jsEAwamhZY3Z4vIN+Q/jAD5qm1/Xe93r9G1i1vbtKZRV69P8PaWIqzi1l
Qud4LVM5N8Gc3IQ4PwGnrA40NRkI8yDhJyuV+dAtzlTsrIlakP8fGBFOrXqjrRq/1oLMPBPvsnyQ
UmVTDlBSJX479fENoHUhk8odrO1915FTDGHwnCZ83wrOKmMKQdIDX1v9j/iYkIR6SlU1JZPqH4E8
I8OTvBmV4QNziJUzCwAD644gBxyho6dx0UsABamB90uzuzrSQEATCODjI12vLIITV5lhlYvlH7VX
bSq4MQCPsae+V4kIfIh0Iaf05SlLwYGHvP/zRVHvlDMuyTzFU+pF7gCQ6mwkBo7UBEJiD2FfGOiG
choYrq344hC7/BitD03mYIAo4ePntytIStY/DkkB7bqoi7Vie8VZv37MkWSc5kIGj/5+4EKBwHeJ
0zITFVsbtP0pVfiQFN+ccHaTYqA7ItzXdBvA3HEhtItUIguzeKRDxlbDe+sUwtymuQb2i2H6uEbA
gD2QELLKDafYOF5tYpJUrgwy/NVObqoX6RKRA9+lJnVzSmB0L02+YqbKGt5KyZliVM4JmM8fPuPr
pOOlSHh8mWMCUJ9HDpD81WUpHyWzhejzBvRWVtPLsFMxIyfs2pYHTjVj+40i+h+Iy9EdyWiHMkO2
UFpyitaF99/ayJohpSzETZt+QSi3T6uHcnPAjFz1M/RT7tRjY8pF4NtEcouN9ocwOTQcC7LrJcnW
yMRU/TwPMot3mXiO1xcErupTaWd5EzXNAFb8V19EhKvhuABvOkkCHooSmaMwb62saz2NVaSH96/W
t/djPZHIBnUFO9zl5R1bcW4+DLJ+Lsrg7kWbq4mpdcTRJ3qJtajQsU+kxhjX55/rZLW6iwCMSGBX
bnkJYswLxxTDgZ55G4uxusTs9gHVChYtnpsjYXi2Zngdw/mdxFVWgVE1KZ9sYLqsDIyG2wwkWLzB
BE6hp4GVchH+0ZobLAe6VoBn4Y4C2ApEPlw7tOGWzxkQKDRMcOROxacBcGSSN3aOcJde9L2+9gRF
ReVl528uJoRjsrpWc8jL3NidvI1suGVdW1uXA4EDePAb39vppKuTZgbA+ROyw9FSUvxWE3C6LoQO
hybOm6dM1vcsP98vkJsj7WOUogxOLECILhZYSnITFXytFqa8JYXt6Pbb/CCoVBItHOt/VC0m/2Sj
tDE0pJ4lnJvzYNc8C1+E400pCSYEqtjVBorLWJ4yp0ixgCabPFkelJhIUWIWGs71l0C9it8LwlNg
8VrJ9/64J8m0LgmWIJsTqyKetSjX8h94m+VBMDAnXh1pVWrl8I3UlkvNr2q76BvJ5WlMLdTTSGBa
MdE6GYvx6m/CAwz+e/yh8XBVwvyBIbF/MsnA/IejVM6jaCuLNA+336v48SxMGa6/DYljMIorsWez
qZm1GslYiNoyTYh0yVSHskAaC6fT7ZH20/vcW8Pr5LrsKRdPfZxoGObkUYW4V1+pPVsWYqxrpay9
dLEdnfyfwhHr9CbbOBhPkA/EIU1pr5gNlML+BIOjt00HD556t3hfCrkmr4HU565ku2WdBycehXxm
p8FQ22GlCLJ2DnFKJHG7uohXA+/54GcSMCYDiToe9sMq4LslnU/0CbNjAQvmRTtqSg7TWv2LwfLU
uNHznTGBPty+5Xk2aCusTtrZUXlMkGHNRc9XOeQihegBHcTcGXYsc1CdyWZmIrWbc6A1AVVfv+Bb
e4SnJD3aLzFWAKZktENattHU0rn82OinRnh5mS1ZFqwjR/9kH4EIkruvco+iGNHsC1OBZJbavS2x
ytvtMAoGeEi2KMu+0rD1Wlv994kjFQEoED2hDyKNmlNkn3tH2VPstZZu3djxe2c4w7pLtMN09G1A
Vzh7Juf5u3jmkBnn5EbgH9liG1KuILuW/OyhjG9EoRaG3g024prIGDxIrAF4uhOzfoGs2pZkkEk7
Qj4QaciDRwWPsutCAEwG3RXhSdah24EPhsUKbgX3E8WS304Gth1NmjpnRHA9he0knQTIaxsRcbU2
v1KiKlRFT4X1dLczAJmqG9ot2R35ubV58taWfHILBjvXEgrGNj+anK3QqdmubqtbKZ0i6ZSG/G+t
ZUIi9phYErt92omsjOc3GhiOhqVNW3dltDvDej+UXeNnsvJqzcbuiNhFgXNo1d7ysxjxeo3wXBHU
ce71pwPuUi8iTt1lxBx1iJo0uTZHM4ikDcu2m1mzQzCA1R4TzbT8YCKRTciNC5QUS69Hd2qpozX1
oTSeWeutdhp0oZuJwIna+oPoCEFLslEapKh0mFQmHnfB1mFeMdZeYPQDjkJaQx3qPjxM43jvygQf
gSL0VC3iZAwLkfkztzHcXsfigKvhQtgB8z+sS6DnbKNR6qCPbfi8CmUBKFC110JgIA/h9SowFoDj
ErJEuZ4pg82La8jAbeIi3GE9Nna1ZZinBQa9zuNEx1Ile/kr4x8HpotZm7vqA1tzgRRJhTnuxi/s
kmeUZvApp2kV4msGNbNk+FpHZUOJ2FKpE0GFFQl5HYvdm3yu/IrS5oRJ6VeG0DxigrvET51XPC9E
FO/LmimdpESDLht1OVxOs/JcmiSQfex0N/apx2AgtXTF7M2BqDIj+rHB4WKCEAnyCHrwndTqzp9a
nf2xCZ4SXUguMZnHCiaDjHiSWFDa6rp8k2RSVclowftMOWHP6t6BUOkqn2zjwCDKK2rAn7g68p9D
qIpdy5ZLZctlFDyE0vlTKsEeGNXM7+VvJ1vBFiVDoa3IldqQEkEaewACz06+2CeOL6Nb5BZZVTQu
3rNq1hMG12b7pLkNHrDzwU7JrPyfzSYti9x4tRis6ogdUMzupS/jN6f4Bud4S41VOnO9NeYb4cm0
qlgqtb7sJpaJK4dhL7wR+iuDq7cXd5nUKFgmbH86z/s+QCpUZu9LEh72eBO1FeXBzR44zdQukW5r
3VRKYpEy4WzfTfczOFcZL2qgFfq12TUs5598fJ0OatMGkCWXmwS/k1C4kITxWpYSDWd743HGdkMu
ebDBrSYL89HYNOByZOsy+c/zPTGxnOIBXb898ByL69+u4tNEHM3PrrMcymTuUHYKF0rzBxwIMr6R
AAKfJjFkYsKHsPXYtG2hbLaNyZBs4g+JJetTK02V3wmWXSlcBeLLiqgf2Gdteb7/9ImXYoCM2tS5
KHiyTwcqbZFwL+QT5iDV65scc4Wx5JdC/GXkLgrT7hVDdA4Dpkb9NytX8iECdv/njkKKle3fPXVC
6YxCEY+g0m8SkkAg8c1sqjA8m7/ZbUwoRzGJAuZyy0t0f7TQr5gVHkZn0eUQNwaUAqY2Vb6P9lMA
dhPwXM90MDasKrjvGEUh7klFTTQqoLdpExuPk7UXS07zsRmWxamGqXJv0EEr31QVawsPg7gY/rPF
HTIonPwVqCZh+BklqUnRL9qGLLLvHTwxNhoZwc6UTY2xxQArYKTJ9zJRJ5J/mwCbgN+dQSGx/AZZ
cTgH4CRyHK5328EpYr2KGYVUIXiRFYtIDagl37EdBsumsXtCqBXw/s9QdPHCibllE57sZYCU97hO
UztIEhSP3hkU6KBSFcRANOaxlZY4NSY09/DeiB8vHALlMH4hkHWBTyXh8YiPpEVh1lbamKgP/MXd
PZphqcnPSz2RP2Zmhzdj1v6RxvbrNiIa8VfpSBdP1rUtNiBaj1BDFfeKJT1XdWtLNLy+oh4wBL5Y
kR0kIBMMs2jTQh1MKch6+XwB6KANccJCBRxqj4SctEwMnvFR2b1pgGWoc1D3NBmgwMlDGDbaKG6u
xiGfWxZSrm3rKvnA0yOMfG89E6Bjlpfr4MqBDsQbLZMke10GCV5dj2Y7aLTgf8TStdEpFKMt+6HF
W69AfQ59Jx61cnSFt9PtwhTqrpQfODCFAfFNflRDBHNEoW+XN9ue3/NGUz31bKO8NwRxqrbRYYtS
0bhKxnVS8XqaIMt3C4tiHHMoXwndD4yYsnO3gS2yxbvdauArOxJ05euXlS1DkGpgGQCWCrGHnRue
tED5BaNk3NX8vOntqxCyB0g8CNzTQw+g6ZNzVnw6lT4+XVmGWfPKZsxUkByBC2TJcacqfYFNq9cU
M0JFUbvI141xVT+Gc+EDYdoOfVvQECffZzxUuq0azKC558g1vIz5OKKw775Kh+8fMJGAmWfudKvX
BNKw5nrDxX3s4vydkQyAogLlQ/sZVlVuvNgOGSACPEZy9panbj7ipnvnJUq1zsHFQCEtck4Tr6eW
ASNaDcbb6azA4VGviffRILjCS5vVbtXzaRiF34Y+8kHsmSPz9BRWJudcGiVlvNFatzC/Blkxx+jq
VkGT4gF86KLshOq33j0KVBFsUv2H7ZA8HuU9aN1NWpMz/XbZVbDNb6ikfHYoNMQHUp6mDpVGDd0c
VPhpPZrX4CmRZgnQFw1BB3htN37xdh4qMI9JJCbCJaxw3oVSC6XMXN3jQ9NusniWkDXEN9pzaIgy
ZLx+g7JpYCskYNKXe4N2mw8wLeFAw4yc5+fUdv3yzacvKFi8SmNh6lLXsP1nDaUom8pggPsYPifS
mB+8qBoPOrpt31MeImjxNoAJ2cCz6Soa760rYNpL9up1LCQ+crfUM5mot1Aswm9ODMJrU2S97gtD
JqQLqzpGmKOMDguQwYbTXK/IWZ4MEa/HpBW/Nz4WNmKn9LeCWzqOIXEvWqtXOE9RoKJu4drHm9Zu
6z78OcP7wBiyZaaRsZqCzNjk99DIyaiwfJpbk60XPFp15MyZPgZKHHQgc+s311REfWteiecx3zFR
r8ooRkOmKQBBquCGHHJFnfcRUn+5loo0Wie2RlG7cmknDaip/ocDaCy/CG0wyyWoiTeR8P6kmPkd
Biu8LZP8722A92wOVqc7CzJNlCQGNLP+0/QFMAUyessmSRWcyCw0bZRL0NyUwig0tvqozPQbx/bo
D0PuTtDacK7MIK4A9u6/nwCUup5ZhnCdGPViyA0skwUQNJjTla4seMn8JHZdXw7+zcbomlLbWkBu
E8VXKJ5M2bzVqjAg4HpAxTmXwcCBYTh9yjaEBXAVLdwdn3fvD8Uz6BQGmR0nWIKRJbANFXb+QQbY
k3+GArNe0TAE9D0t7mc742G7nAyGXShBLJgdw8cOhmx9m/RJiidoPAPT84eUzERxB8i4skWJFe6t
VVHnxzrmrKu2RSZVKYaOR8yMhJrRyIIQuPMeKUoPjIDUKXN7hMEGtH18EwnEC/Bctgyp
`protect end_protected

