

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
maG5N4mcxNMv5ki6e25fu3wzDZm0ZTSzlFqL3Fug8tlkkCQuH4dhwgjjbU2JjtG+sGIdWDl4oKws
zkzQ6HslEA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KR1Quv/2+0ZW7Pet6KTsx5opy7Wi+3rbIke9CQGCJ7yoNHVXOqYjWlYz6znINSCOH3I5UuGSO0uS
nJ+wGAzv+B9rqLLyBb+VoxMDx4pGx9THQTYXhEq7LKvCeMNx9hO2zDcBJuLtSmrZh3FOU7nyE9q2
C35VPHOq2Vs9fd6O5+w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mS6Plnkb+x5/4Rvsi56Z1CtPEjpCD9vPk2BCfi98eB9E+AEQC1ptthM1O5v7E8DBxXfSbONoyOut
nnC4h20txdR44l0MPxo8FVucsN6/67mHSLMg0jRCqcAZhUGkVMpiYF48Afc1btbnoSXE8jTJnh2x
+TYNazR3k35kFnHwBuVsv8svjI5nOxutolrhQ3rGn/xRBD/sI4l0+QFZ2cZznjJtyegrdJVoxMJA
AnM0mbl2i25mmP2CmgSP56Qjly26te8W0x9+yYMGShwk610vByf34BcGi0gHVPKcPjsgR6OlRTWM
xj+9oHAnqMOCWeRqXN/ceF4+ecHDMfx6D9Ib+w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DqWipD62syRHsY/gUzM396cqzKm2gsbDUqyq5R7kromixBzPU9bVU6CzNsNCiQsnSg3/Y6zBz4lJ
dliX2RwDE6+FfPmvCK8VMySdgbq9XrKb1mVGgWraxHRy1JqG/MeJzox6x/LjOEQOamRpre2Kh24w
JvAE/LxI7sFizG/pLLU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X6IBtaOk6W7HSlW/D5aJLoctHrM5bNuZSNxOFnk+5aflG4etsaZ/qhMPWADSwSUX0eJ0nvNp+YOI
cckeTEaO8qV9fJuXfO24cNbXqYzW8Nrom3ciJIxN5FHpiq0rI4FbXMDLNAdbS3c5efscoeym6Lif
7OAZlg1gWMP90X1PpbpbUQHtXonnnNRSFTyGBEKNo2wfWZOHaH2llECSLauFG06kdQ842CjlwJaF
IchPeRI1/WVXH3pab5q6NhbM70NBvSlNrIC37g0F3skvBHBYoZe90BH4cX240u7D120iiGXWP2CR
r9rRvUUJ0K0v5UfUfHAu1nzSot9VNlHrkz3Lqg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103072)
`protect data_block
FQJX+sDnZUX5DDtP8K1UQNgBUndn7nlEsZ+GdXwJYXX9KMS71kVpweDlN8ikIXil3aOtSp58d6LU
w8ZPT2+HrioYlh4GBTpQk8vzDyEl8aRFICe3v0IAeSXKFey4M/2+B+7n9AZ+sTyzry6P+MutPAS4
3BHao4AE8AcW8/QH1Aozcs9zytQIABw1oENXSBRB1H51sFD7arVyu9uWUPnUwGRA1E7KpCUl9h1/
LxHwo83xxRmolUfQMt8JbFFYsgR29Kwpf8FYZFJoNjzTPW7dOeLTT5TabVI4Nrh7GfA6JTTE0rk4
nv3+Xj3JQLLKQW//Dvo38hdImq8mxX5G+YWd3j+ia1hxOhdtdwb0oWz9xwpmkHhYfSTKxJZEOedN
otMcMB0IWNO1i/FsJAvIsDk5MF+dv7hmkZ/4EI4FCU2P6HgwNiWOM4KbZJSZG18ng5f7+G/VOOmk
IiTBe+cuf9nhq1gBOfeXH+Hsd9wklahpuk0B5Wh2z/QufxVZ+uPrROa59Hzxik3w3NmJkmpov/z1
7mdX9rajKECKi7YUNxIxAGtGT+e/2P784SBzL9zgv3+d3aWtUy0ND28pccTKgsBkhLsf6D6us9ry
ADS4iLJkR4xh83PyV29dWmNlfq6jIk4s1zmVLiDuwHBKRIJteKiOOQ8Olx7UkODvV35eyVv5jFNr
ckiI46CsgiYR2pS2HUleCR+hivRK1wjYhsb/Rd27q7jwUb69UyzwiVb57Q3fx84OgpxGZjlDhA9R
jofkf0lTkP4dfAXMFRDqjhhWZikuyYjjegYAQ0um/c2tlmcqgkwMQcMy2J9echxh/nV9Y4vucDa/
5zW2kEyiuxEAwqwdzjKBKWTMLEavJA683WIcIboCZfQp3ENAD5/QqP2rKjd0Vyhve7qnhrNshiXO
j2JGL/bVZtFHkhlvn/lJLP918OhENWfVRnY/Slr4/K7/lGHnip2MlQAawCbIDElFaxqS/h8/8pzY
LRWAagL3FBubExt5ZM6PcmePtZzUwXAmFnf9bUxYQQm/jsDHQ3iD7qY+7TfLeDzXxImx3avgSpWi
nFazD0DPSD6Wko71qTseCG0/BWKUpmbcQVoCOb2+0sCS5hSEJjE7WkI95Ze6Usdq1JWo9Yihrxpn
0E/8yfckEW+lgOURyTbwFtADn6OI+MpWOoddH9ZvWJ/dOYHc4CshgU0s361XymGsjCPlnuoPOoC6
dKAxAPPdPHXQM+xcg2Erkh5YUbjGFNaWGpDJ27T1QNXOmMqaY9n4PDej38uuEkckPqQihCTipegr
NLPhtHKZ7J7kQk6ICa0pmeYMl3fpp9q8LSJIkwFZIVtd0kFWnEuWJUto42OjQYhdG6oYBin72411
nyXK7heZIoJG6Vg9XQdf3LbZKmDARGpQ92X5dap/MNsxObdhNBJjHGafx3lzB9dOvsq51Npj9qVu
mkAE4ALfHpJYPA5lBqAI2agcK/IxA9DMtzTwSqphXz0ckos5PdJ53+pDzcgiCDNi0AHvNNtew60K
jTju2FSQP0sSv4oNgT0AfuX4zzebTFhqJJx8P0rgVWgNRPKPTVzmFxBz5K4JauIOb4Tkmw0RHs+S
w0gk9W/x3gE4qzX22IR0iE8M/UqEmRlnjgIVxq4cX3LRsxhOjXEMCurE2Z5Saw4SpPOWTP3BqNmw
SsqQfgb1MyA5t3lxjJiQkcSokEJGWLDv7X/FNd/+R/wM2nbF/uF04SmbFxjOwokaRbDstK3y42x3
o/VKC3HFx5S5w+GSAfz8IPzy4Sh3Qn3Se7FRBXJRQVpMxFfgsVEAMpa+gZFvxsAA9tamMnwHCqSX
EwXwJ/9S/HwZ+5cEB3C2wER90uNPQMw7SctLBlM0rST6bgOMYKyhfu35MD7KA+q+3XFi91ZaA6A8
KoRqwnjprfPhv37IkJKhmIRKU4MGsXEppTXXh4QqGHI+HbYW21cqB1M4BY1DgMuG4OeOhD0s7xJP
ex1Eze7Cu8d92Lu8p3lGBisgvD+/kDMnDl3u0x8fJ/al6znc4EfILXNmxP1vxE8KWLT6+jRzAhbo
1vtOJUFI7kqBFXOFZbv9OYy95SWZ23QhxEw5VcN/0WYT8tPkleT8VLJ8P9faZo6zZTx9l+KCj3YG
Ia64FtQwRTIspdzkeZeMbaJiXE+vo/rC1UFSEDaB6Moz4jlFOuBi0UIyNgjixb05kUsIC5P+YBg9
FTssNKjYq+Jd+MD5u41tkD6Iu4G0AQ8vynkCmmqfSqLlmjS03WG8/83YrUOsySGOmglpzIfVTQUW
bjSVKEgGEc/lyI9XDvF4+XHyF0+dFnAYrv7/W2A9z6hEIp7U5UyCEj/QeXj1olQ+bhvKbMvy4L5o
EX3pyNBi/obpTMG3GVbR1z33Zlv4w9EEb0PiwLDgKhI8pqShx6Tpcmr7tvgvHx8yGQlhRc+zWHSG
m1HxTvqp9965gOfc3VSbCSXplwX5ed9y2d6q547xeH9qw2Dlq9nhewAWzLqmV9hMcOkt/NTOwHSL
0AYKmZNMdemIqeXCMkhrn+lu9v29Z54zDE/eakwsCeGtzR59nhEgl6oVVaVV2s7iSdKOglWA3H+q
C8XGpSEIbidVcOlCyRf6lgxyGIpqGnLweaHGgZ+d6V3z+ke08Ze1YwYK5EGZMllk06mxuk6VK52X
CD9C+vpyKvrki5RjdYWONpKLvWmu7A2Z43wcOgbAPGMXI3dFpkZcSdJ3CUHhKcsztNQpWBrMBSdu
1ZtLdEFm7NyHW2dx4BBVJkB5GNgHAgz0xK/4wMFpWoZhjveAU+qRSReVYtTeEFWQoxtG5adOSyL8
5NtSjunFB7FZAuiPgmY1hYaZMXebsHu72OpRB0yx/7hxIVia3iCzKt21xQYDmC2zQriJUux2i/oS
0ast+Dzvk7zhXQZ3G22IY/yLveJYL5XZFASrbR86G7i4gQ01Gv8f7mS1gISR++R3nsKEA9x8B/BR
+emfJv+DHj7CjlJQm7AKxSKhAJ17Uu83JOKhbkdaCfuV5n7c4IiNVRpKzDMsPScLJLTrdU3au3vd
xkoAtIFAEpYuK1FoTJkFVYeJa0cpDXhA65e8Zt+bA3nCt3phI2s8CHaet23tP287Q7UWFCaszDNy
CRESn9IS7uUhz5M/c6gv69nLsqOwTeby4t2iy+h3Sv6tPAaz4azwc5UbX7iEOem+iaS+D4j0qyfT
UlJBjfDuxaJMz+C+svk1jaN86wTv/pUFhZ7R/UBdYoxSnLoCMA3y6gFda+awB9v0wsIdpfS1rVKE
WRfRnFAXf10U1VnfyMap5lx8owJ/mspkF21i10SQYGaSplhSe9BPlQ4UmK7fwH0mb2BTyMqHTZ91
fdZXzUjPXBxYdG67u/UsTUVW/QhXuobZJ4jqG2Sv/ENS3Hu6wGiUUOtFFRasfdm8AfTCAB2qUS+C
cEF/disIS3jJQWZvxpwNwnZQ6kXCObtQdvGOd1kQ4oJX1zrhbpHrm4ozrQPR0ZK+Hd7KZqZ/TFFG
06JRXEoE8ZF712o/pwkJLSnJqrMa5GZZRvLs0oEj4H93CpEU6rtryhzcXQx3P/o409Hd2Qr1rhLT
nrax6KXYhWCcAxwbGJ61xyQS8gYZSdURcsV11CsJJI9eOj6zQyvd8P7Sru4L83T6GInb0r3qFyCX
3z2XMsLYioHiQoC4mub7EjzYGYX/8NibhAfqPDOT24mQxNfzPlJgAgumsp3zzkq4sdHmNsPffFhp
elI8WC8Xfz4oH/snrwbqKmyRRM5QxMa92NlW1ypvS2sGdyrUxZuOwwIguPOPqLq41Svmhyv7gede
WJU0RdTH0aGLkQmH2uY7CfYKRAe0bBBzOh0/hnwqqCwAF6zXeClMWDe2+VPrPSjXgxuDRxOMMHSR
09Q3ib+q3V40Fci1COZiKNTYDvVDseOMnNSuauIVSup+ilCmbXMzYwQONT6LS3FAWkmXd8tryuJl
JE1D4y/oYCNFSFvi1tcVXA4BpHzus7+CqZ8gf4ilK3Wr7MH7qDzGr+yIZnFV0mFVeJFHiOvstynQ
FXZ4aZ3orAbevLzMf0623DCAf/PhO+cMnkYx+PtTSL/YDXwCNhjC4WV7YP/xDFEywkoHcLjHogXo
mimun/NXBGEYyMScferlp1TD+zQD77K1lJeO9L5iUMq3lb4AJxxOnvuxHf13HCUfwE/+Int6O36+
vkaic2zzaA0JwxS7DpScSfDytVOisMgV76ALtBMJ5xDZ+DmBiMtx0uiwF/p6UAJiq4PrIQ1NLdCP
PFxk2gCX4eracgywOhcuhdqsOQxJ1a35YMAmPHyayEBR/Nq2gQ3mcERfADRvJVQriH1hY1kPiCbX
EmQt+pjeooU1KYruOogCxMc3m1YL74ltQyXazJnZ/lsFgIEoPEQMx2wGxafpPBOWPRKtqmgOhTZ3
wTOjZ8qbUui40WI8aa1YAAdUXbGco8swJp3QpW3dYNx3jiBKffscIPZowDRJAPM3hh772D+WEkV+
Wvjbc7gueCnVRg9Jp8omTFBZv/7AJWLMpmGXJAyfWu8RUMHP5vgRdVqlQEpj3GbaNDw0glrvzxu2
+BBAfr+0kbDFHbWsGum5y1dqbi2aNhNGRJV0pllv+lSRAfy2cYWFxEkqxeHt3w20ntRMo+pFb+Xz
vqXlQHzLjCTZIUVb3WawCapaUC/RfPuGKFbsVYZ/Zo3At78xyF4Iz9qByPbGZGwm5DcO1G5Hk6YL
Q6voJMKhrkctrRlYD5vdl4YCS6R0+gU/avP5YYxXhv6vOdscvvnc84fRXIW35vv6383imKCquzt2
OLAN7wxFR5i/JWogifhPQHOS2Dac7lAseajYDQTn6mRJJuFAfrk2BXpCeEaW7i1yzajXrz5iXbBU
4vFRChKrLk6bXbiIJnQ10zl1SmrxrJ7qJtSiiSqG71eznh+PNUbzNe4WzGDrbTLejhNPMUDcktTI
yhtFiT61SFw5JDu/DNXTWCMdMhJEf8zlFN4HUFh7631pXb3zGPLuis9tSJ57o3kAoRAm0PvXWQav
x5QRLAKWw1KsgyAQz+y3rQTE6nIzu5YxWipEueD0mBSbgnXLcuIN7ibUtFQ2cjqFPly8S9APHI+e
J45guntV4deW/ZaszU1sf4biPaWMYabkrDelbiC8Bh0KHqRTgYioFHbVdZuzr+qUJXcLCV4oEuNW
2tiCPeWIwQZoaWqhZZq4eSVhAZkzPQpuRudMLanrJNtKfzsQAudrZRTpsWRgjTJFqXEzugziL6B2
SOESFbF06oBm2fvJ+nEO9/cpNKBGWHnVV6HSrf9jYzs2h7YLxngm9JRvcXFswfGktsnzrBS7s7Nn
leribxEBVVFHUi5lDM+np4IAyf5VdDRqwUjr5Jk5pOR4kwzVfw7ksBmJVNUnHGtkDDC9hCSpUhAQ
mUURSOg+xBYbtSn97nLfYQs6HZUC5SfB+NH0jJ3gu7nEB9wC4pAGkc6lAE2DRv8C08frlk8Ps09C
H1hZGJqTtyzMty6MTABy0GBxuWkIsxJgyXpGzgNJQKBa50TUgD27XJRzywdpQhs5nb7+XGhiB+to
pWrQjJekyrfZxqUlrUh4xekpFCfhQI2uECsduvOCeeWRvHQj9AYhciIDwGb8qPObkdLwy0j1QMrz
v+jBYI7GBd1ZJmXe3ynN857+NgBS5X04SZQg0iHve8NrFjtiLZYVEJM9UFJ4neRy1m7UYL8bzDAd
XzfFGCj6pXpzm6oPcoxsxu2KGD6iVoYFNAHigHGN/MphvhjmMm0HZOArzgUeT0vU+ZgGCXXvaPOV
HevXxFuFqfHtG5nDinMw2/aRYAonsN6iF8vdmnDSqLbS1WwalEBE5/YuzuYzb8t7ybGQ+yByMXv5
DnAvom2zlwb4Y1xo54ZMprC3q7d2QiRDnHs47LTMj2zFqh4iPysph+0MnnQMX5NTArpRrrEFmqXF
XW4copLSmqjMSwSwSWA+WBNt2a/RSWrbeGEcXWkOxJe4WDSBX6Ka4eUck2FpExERcTo0iE7dlXS5
Vr6PU3fmXKkWO6iBGWPQvA3V1zgZJqLXwQC35eDSci+LzWmbTkkOY4y5TrwoprHWR2Ntx/XO6scE
jd3DLp316zrVHu45CJMYvuDS5DJDj34bO5bhXWjCecWxv7403mSccwVJv9lXRhxvqKfld2j1n9eG
T9u1q82hyFZQWcGf+o+KeHP4eRvbvNklJEzuu7IVMefrzsQoYg4aWubPa52aljTyAQhk30FR8gye
xhlm+PABGqLGYv1Puj1qUxIxG3b/il6pru9H3d5ksKzCbRfdDdrdypukBoIpMOYA/R2l8C51Dtc1
0i4E/4SgqdD9CY34LGIEvVFKgFa3ailvTak1XZg9M1GiHxa7wBnVZ0yt1K368XSzuZ8kB8EjyF9l
meDXADPLx1oo2GlF4IMYp43wIBNBdCGEbe4n3mCHy7labvYRkCy1L8n8hM3un++Cpbk6uIW6+9Nb
kPJnciAyjPMMc3oyEEmf21+ylfKGO1ss0riZ698T0fRYxikQMmKZiSH4SNBVLIyLuyYzMas/IVkt
Qb1IkfTSG+bTC6wQmCsKOEX3gQqxAI5+mVvR/3ayPpM7rvCJZORcjGgoFt1AF/tBfU00GsEjDBFB
+2j2N8O3gxAAaSZT3rjiUoMui1PdD+rLjpI785OoHwIcnKp0IGou/ewaPeoQ3bdySYCrhQHP6KFK
QudTW8HOQGb0IEsvavLdFvrTSQtS704C3oIbPbvW/V4kQ924drHz9y/SV5iOdOxhoovx3ztl5h5h
ODmz84S9Oeug3BxJqHYo05WzTYK4W+2TYamiyhVOpW+7KAFHyHct6m3yV13khAVOmVlxgx8OVK6w
/0MgQpHMfoQhXaG5jeZt15B2b5ZuzM726W5yU047EzgdtW6jqq60NnFtT6KpjpBUQmKPuRAfV9QL
HFVauWsQHXTc7ZxjOqSvO6kE8MTzy9j1wez2PFGwkyKbANwosecL2spHp4nIKOxd8Q/+YABJZJiD
klbitwTGLjggXIDKjzLzDLlKQz1qai40zYYTwSBDJ041nyPQccsiZjojfSGjCJE7/oJjMUMroAzf
rL8FiUvgvpgD14JD1wlDqnKrOu2UlT9++rH4sj13zIPLwyK8yTIoNcb3/fNv3Z+ji37hB6+5o3V+
JBStuzoJ8plP0fiNksoN2ZGYKrIbhmu+RKL3OPZ8IkNeRq3S0OqdEG3UO435LQUutt+bkuqoYaSI
xFTzrPB0M9S0JFA69YYjCmGbL92Qc5IafDM9B6wtnfJtFiHvTAYeh4WxbDDr53YhnWRBPdnTy3rz
E9UCZTFAROlQhgXLG9R/wqsZRBJaChxpSjqBHGtjTlxXpszHEtP1hQ5LMcTDMwhVaSihygWJpvc7
cc+ZMlkJbIsj45jjzARNCPRlWixNswjeKroYx0Fh8UtFz3xY5I9jeCuF7QUo3ypsR1X3sL3R4WrL
f4s7K8hOada0K416GA5lEMlR27rCKa8vlr8wtBL+xvqAwXiK66m0JQCT8K93qyZ5Qm/h7CWWfl/C
UvKkhap9LQ+R7RsUlcWgKc6TvFRAsNePSv2qcA2A9kmXK47vqQgGWUYRuIGuVuKnWAho+utePLB/
SauqwopZh8+jfcumJpMfBK1YD4PZhks38+Gfq7EwhnMf/u9wD/vSRaUkBuN3D9fu4fSBrAHSoJNh
lxGV9AwNjcAu0uQIkhV387g4BYCJ9VBLFV6eaNohJr91wlH0h1d+1VsAWCWePFQ58RH1IvK/P4LI
g+ESq5/+OV5qcTYrjceGPopKiMDXrWSTtrRjBJzzM7uh8TGRJyLujDyqYrAs12hc/OYhHHkCipjy
hG5Tz90R1VHnYLFi0SAMNXC58HlZ7Tzkg3n6urkmNTr+Z9O2zE003dqBQDtsYNlm3z83/RBJGqHI
ggdahRamrDxdphbyRRw6MLKm3WNk30GlJVD7mWe3GYA3jUeLm11+0KiTwlQKI5aOkmQdGM4BxC26
8s8IDW9OxAf9rLiXLkPumyXoqvn1owE4qJw1vIH8L7zHTngxZyZJdCE3dm9mta/J1CjXMZ/AtsVB
7y/zCYdk6N6GIGvzD53uO0n9D0xZBpnJ0d/Y2N8+pMcWvyxEGNgja8ydjYKoXI7Qivo1JLZRcv3H
zR4zJOWsDVMACoy+PFziajlraCoJHQTLtd1zfsAUYV++/AUAAn03JMXf+lqSdqxvo4nBUOn9rwsX
HRu9bbI3MjjrcW4g+b3gQ551aX32U55RO+yGKdGskfmE4IGe6sYgHxlAVhE4FU/cisCWeG4aF5MI
p8OZIK/jBLkwa76ivk2QKTiKM7JqbMUHJHEhLffyWVP8xoSauNixlnpcGg71NOndzW9Hu+IQh1m7
NCAylKnZTzOp38HybCK2NOM54DQrhOTJ3lynnqfEMY3OCtGh4pLk9baI7o5tDrV8ICmbzXfVTTlv
OjfkAdNHC70F3OsnahO+RIhNrZ8oDobf3/xru1IsdNDnCZOa/fdH/iT3ebqF9KwM/Sin+zEq5aUG
UnMPpgnIhKEzhGrWXsUelIinScCPrIucsxFJsWihQuWMy61JmgKPiX8WGm+vFxeGgAOgzkmWeC5d
0OcGzeTPwuxYJ5ZoEMJSFRPcggWY0b41KUrafzSGfpKAYfIOUa0DtWsj+KoVtrR6Z3Xa7WnauwPN
WOYa4wizq4X3yQP7qtusWh/NqiIrHhy36fJk3lSQPbyKS3iT9aP6ukFIO0JYUDq4fUK3mYG2YRIE
WVL5oZF5kdrIENDcCmeik0EvLTR+qZCD3WDPJZOE7ngj/t/+Vg9DdrsRgMWVIp3tvg7bURZoXtvR
ju4xsklcKyWmPmAnWuYxZauGf4MPxCCCHM8cC9Z7bMJ/Inu8hao21auyPETzzDeuxJwxyZ5Cu0dR
Msf5v1YGD+0k1WxZU9bYPa9iFNxaYnYvVoN3BHh0BOwNsxG5EIR/TfPBQd3RXNcmqwElvYQl0RwN
jhaGYdOItELMsUvkrpWFlgq+w5/0XY5NNSOMqYZJj04uMkF3JMXa45JoKfwhLVFWpa0sXx/Smf1m
NoY0i5b0qQg1ALNpO/TdIpc+ZK0YCLo4XMvj6uuM7XL0pp3sglkGcohnl9fmhyv2M11dOtuURUZM
xBFnViTx3oFajWd7DmmHwuS8dyML4fMbGHcDeHL6HNrcjJI8jAFUeof9+Xx64+846UBj0j+3B8M+
IvbIbyhMeXruld6s8b41Y5NSmlJNM4QkZSO9kBP3shLGN+/ZmD2ZyKOrQTM/F5NP2T22l+LHEWS7
TUFaHeqCAdzezJy5V82OB/6BRa06k3MPrQ4LgKvpAUaqewP4ZC1QUjwWf3jjfpvX8sbJbnHaBhvu
kv1+gF8Za4gPXJGlQdBT3brXjOCyEHowSyjwfudhl+78FPV/5mMhdST9ZsVhNhfgfTGaxSYXJ1dt
BiNBd2MYXck/OjbSqZD+7xYhffTq2WFrp+jQgOBzzDEqT1T+WCAoVyc17Erg87Rdmx4FsoW58NU9
+xCDkUAmkZbUwcwA32ctBfB1YteDeVhwaCzMwevyjCQwTRsumZBZkGnjT4WAn35unx+p0qnDqLgA
2eVUgkk+WCgWFtUv5PohPXLy+z+ERlWGCr8NYfRV5u4ZrtEGyOXVEus1NRQlKORnOMZ/kdsU8EwM
9JR/WzbceBhDEwYUQmExGfsFi7o1QC5bgMxkYd+6LiCHv3gTt8l+UjFtpYCknuyrCJ9B77Gcrerr
RHKMSWgucZkhOBsZpzN0onWg4imk4JdhpgfIcGaLYf0M/ZNOLfcp+LkdNDW0I1/rzsCfliDO/Exr
3Yo9FediWXaXMFFUM2gboyyfOBD3HJxzt3TPXNarz/gXAYX1PMl9wvepKXGXxC90KPObJWEwEgmS
O0aKCl6jC4TtBXDX3bFd8ObTA/8PGo7Cqr2iZXi7aR2oFQI3xLYQzZaTnPrNNbkC2JY58ksqkPQX
WVMZkDF1ZVPYOP8uXI+mTmt1YNXua16ym1JMukp7ld2wBHnyZPWSf7j+w+CkFmOloKiA0rMNau3b
3a1qldyG91uUe6mffzrmzXilGnTUlohfC4DARpJaGdbn2FW51C88+VxrYj4MtfbUBRQztpPSWbjE
yexRcz3sYUh+4xrVWvlLExIeh9fSvsxhl7v0g7TBIrDJ4fglt+UUszYGd6SiYmwzAJX11wTU/Pk5
Ls6SuT77+joy1v9NsHtw/XLAlacrMehoKAWsgYOi4xxALPAg492ewIsXIGbhKTJ/6aB5s/AFnZNn
djWPALVm3Qk6OhA3jEgMycTGgJyU2OUJK7InQQaEmbUnV6iu9vA9YKZzVdxKnDJCzRrFEPhJMoZ2
3w8bTay75ji/nRYfkNQIHh5HDfAxf7N20s5O0lQ0B1jGWtq5b2RZLC+I61Wcg7tt1P6eEvjJIK8W
7odFTQqYebGuxKVNmfxpZpy4w8hVwqyP4YuV0KUKTRPArWFG4YBeswrrCkW4Vk1bNh7accK+RHip
+qlsGb7N8jkIwkBHHEcPF8fE9zIYve4chj0eMUKqV+/OyGedjeK58gQEwjCIt9e2ReowCLbfkdXX
7HhL8RMJpZLhtnKNc/wkxfgsHbR0MrCEcdS/iwOvDiPeIfW9BzwDwSAifznwnQASGg9AzqetZ9cV
+FIwjcJBOHXQzZsnIcBfzKnZWDxLuxHk2zwlDYTR9ihNDe+nc5UKA6zcQMOJFir2qk/2CiVVp0AE
zFX5Z9lQk5BAl+HYzHC8aKP3+qSxXK06YuWta1PYNHodzPuahBgBDM7zSZAw90Kq3WS5UbX/IJ2H
7Ud06hUtEDz1C5rcaMULcgROQuB5vYbbaOf/zePC6NcSftDTXzrmr7r+xg8xcSfWdbTi4BnjA0wb
VmKZxMYlZf1ZL3FDP+jzD+MMwfsBSd1AK9TDcn3hFfx0CsMkfYfqIG8+wMS8dN4ZmL7aacUanP/a
2eU/nuo0Z4orv5XMXeKfBXgoPAH13kI9q9r2DAqH6kVeEuUUaDczHT1BS5Gp5C/s6IZwh69FYPm5
7YlcYQLGsCK0LmZp1eNf0UaIVoc/9DKVsVkZemv2dJVGU7qyE0rz1b+h0StCTdb0/Smmev3W1S+N
wiSTOMdXxAAGQX8RvsL0AiiXORYXsCZf6DNTNCeGx5lvv9zBkU/MmSN9Af10ofUra6lOLaiMoXHb
VppD1YQt53Cg7wxHtqGlGjrD3gAdZLaPqGfOx2FKVFoGKExp58VPMr9mdvouZtD91g6wTRs9KmGg
pzO4DaCcYfiM+vYKpxirxPIR+nGdKG/5V3dXD6bh29XYe7SB7braW+b6rnl8y5cAyOtfg1TG+ZUb
2BtobCNWr/17kLph8pvHBtd5TPAdtIFaJrzKlGeGPrvXDng0SDMBvSL3qkQehGg497zQdd8bLipf
AaaHFH55KW/WvKmGkIw9uT8FISxs1khMsxgoXL9odH9JcgI6gOVpAHBWkj92htIi1GvgQ7fzbKpm
vgCqrXIZ20MaqwzmPWjakMQPaEsZT135sLX5996++XYq5XBkcCf/LwFLQ/rG9mLPCzIb6YszVSd2
FZiY4LmbIbYJ4i/12zs5jbZFpu8YQJ+WECf+F+VEH8T0oWhUwQ4NL0VGKscXvKdb9/qAu5OryI6d
VP1SRvLzAcCCuVBubq6PJbyeQdFASyM/gXCRq/q94dhFzz8c3w7lUdb1fTqElONkIGuijsK0pFKj
Yy7ir4myfSSFhZDxzddUjQqLYQjNEgTUIYzdDskv+NJ2Fl4bJnskQgKEjLmfnD+Dg6xP4RfDkRjz
Urp2uxrTufXhXNZYIOg6B5Sk807fse7wPPbBbyV7Cw3GUC4BohNv3G4WDj+YiSPo4FvwwVyv74SE
9d46nIo++kbkiUfkdkhyrzIJJdpuctOTHq0pKKm4lXFo9tKvdQKsfsaBWYPHv3KWfhhto8dqUmQA
L0VeSlQwSD14G3M8NA5fj/TX2NWmDQc9Az798IFEc7iXeXyv5Y53vqhA9AIF4w5iDboMOXnD1OvZ
TEPsXMi9w5W11HR8C2hY6qr42LDeMLjXHr2myvChQG4oOaoWNedmQQ4yy6HpZJC9oAo5HgpmwFj4
iKs++yNbtHg/83jvu5xIcN+8eK3NYGn0hAnB7sUaLz710LWtAwp5gaI8gNITOuWkgW0SUXRW+Op8
GKxCUGw9r1tw0Boy8KADKm/IIqhMOKeSXF11ochUF6PwOuHOIKZ9VtdaevPLu6IXmzDcdv61iEjJ
pyV4x6SCfi15TKMs3N5YqKw4Ix9pQjcMjrNEcg9CVnWr2E6MWbn8CT4Hh/I6rkTNiawdTKgiC4ed
IrKanzHEFzdP5EMAPrpf97nN6ikA+wG5ktnMBXSoW6xPcMfNEQykjPaLcwFU7MYWgy2QDijyqvkh
Oms/SZDK4on0rEU84aXG5AymdKss42yZbB7P8dZ5UPowoVqXp+viTJlhv7CStuXWSO4zYz0uL1lj
9yn9AE6fHVNA9aNVQtlTCHm5zb50Tiyqxzs1p5VW8Su3YQN1a0nC3ZpatzWrBwYVmeVOhyWdFCto
+4X+G8iLaycTN+7N9n/M/rfx+X/ucW+hCRW/AKrP7XbVQ59oIA3tSZ/jpHkdA37tzGLGu6OnJRjJ
qfLLZBC4b0e2pQBIOAO5CKHEZnEu5usIEqUR/jIe+87+Pinx7PZbRXWoD6opw03WeSB+V3Uk4GgA
6IjJC+2U/I2jwerpPTZsBH6RvDlT4dPE6HbobtbUViQftzKQNzIO+63qBhwClbkqBcYPLH5kyRF8
aIeh39UmDm2QAKPQHHi32zhWZvRyJtVRYcHOyUKRQFwCbNACdpwurCDYLmqZsh4iUdXYJ2HY3Ygk
+Pq48p+8uXBy1xGhy0kEaTZiKb65cQCPFrkURIqDMqEMNMhBKH21m5bEnvKUjCnRu1EsvrLHfn7k
SArI7oGUvOsMOmmuGxAVQ7NaTmU8hQoyx6RAL0rsc4qJHWxRNZtpkWWY0wHphFIv3Qy7RTD63SaJ
X7nyVd8uWVNNvDBt1po9uWDQtGX/sP7qGmrlkUblnb5eidNmRkpEX4vU+lI7sHKmLSEDIXMPvwzu
I9EKviYAZxiMQsbVSwHmFrk59IKrhxhzG6V/7F0oWLK3qi4GH6hMlZVeKsYWXJXVJzxu4RaeQqpK
jDqIpwavFnB9GV2uWk8eApmNcUl1/QVTBxWsSJHiYm48vbIaM1SjB8hBGkmetAIOfXizyEN31fib
VRaOio+Ej36a3e3hZOAcof7P+6nPlJxIZxGGBgOszX3rO1ZrhHRnO9HNuD8vPUVXV3yH9ycy02Nu
zsNX+cGpaWnsezy0FFUeBxzpy5K5BaRP/99IQycc61lD8jzI3V72mCvYbxgHjhKYbPfNNebTNDQ+
5sIY1VbkuuXyss7ZS6FxjF50SnQpM/DsY0tXUulVhgDZPcCetYdr34LxTk04JVVo+17XqC2Z4RU9
IqYT6ehjm1W3uQcDC/bEVvRYAiWBhqIj5WFgrgtWCY/gc5j1uD8gT2gYLCtL9ejrdYKtcVJr1V6R
trFhSdwRoTZu+WroSXpu6DTL9+Gpvo4pEOkMjtyejdCe4FCv52T/Ttk/HrK4Lcf7rbqaFk83BS07
ooain2200L7/hemGHtpx2M7raHRyXMlIakikErbKOMXCQNUN7ttGHhYAxyinGoUGbAfncac/l5Mi
0jFbsZCmHwUTt6KPuq5GKQm0AsQu7TxPd5C0/Hm/Nue2AndlFgIJslGPbA0d+Df0H9AHlijwsMdU
XUAafmC/ghphnDlLPmK7U3gmMSrNMEobKeub/8H1LPdVsLntEhBgujNyTibPkaTEcpgqzcWWBkAl
440iWsdQ830xo7ETW984xYmpfRDwd4iXua3NNjQtbJEVC3WhhTOaB4mm972PI+2trNNyC6Wv0PeF
hH7o7d6zAdA+cP7fEXLXXpie6qnEa+Nq/uspXn5hcB2D8r/ZQrdcMPd+D91WtG6iRU4+diX5G1WY
X/Ohuzs0Nis0FxSNppwYXnuhkpz4C5eXKKA0yyRjXkuBRw/mL9CvcySgfaXKrqj/ou8oAL/cyTV1
lYWAL/fzyH9HZAqTZRY2DtVCanj5H8iJzKSaWaKEMyQBYrPdxoQ9k+vVij1yuqfJxLVCMgzRSTFw
bOB5UT0Hiz5p8KkDqMuTpSH50fczUArdIh0PFiqNKso/kGw+9KPN/TF+Tee5Ri6xQNz5ByBwaTNZ
vZ9aTzke9sRKfxz4cNq1Pm/lGIizbOn/hIDo3AJJMUEnVseCNJzywdSWYJbyXrZA1OjTIRB1C8E0
SCSnnkGTu4D4/GSU3KiNVZrcpmJkbVlrVYpJ/LpXwl3ABC1cjiBFyV5zrRFY4cgWetyM1i1AQ1gv
20K6te7RZp/IxpEhiH5Ivb3V+9p7HHAhJuuJW7BIQydf/8d1ROWCf1UjyXR3OtvalrW/Jm/HayuB
EwCPNKCdv534nmrig9bCYs+ArNhRLExY+2ywtljubEVS1b68dY5/CuMW/0mS0/LbsqWjD4ZYxwou
WdRztY9WT93iftrhrlKLO/7qjqUQtcWKrMVWc6MHYktJkc0ufJVWvi9C+jpOK4QFpVas+bQJaAqs
YayPYnRVgq6PM2uZzGBMKec+MCfpiMu9FAlb6tH508F7r9LXr8mbc8NHYKL9bdUaNk1IIjodh3NE
UUx2zuuXb3MRz2hoT5mxP7vt6ySWhY9sw04EJKqgn9UFgLXLmrJTfkpSZ0E1fRQwA8TTakr5pek5
3XVUwyJrI/d9lah8X0bHGflJsXJxiD5Wpov+NhTJ5E4qsy2OFZNTEQtP5EZ1bQVI3q5zqyy4jw5K
7VJN4OiaciNHXtGXzqcCuXBEHAMggM/3O9vwibfTtb6TvD8DFdleI3qO6DhxuJYL8k6A6w/sN2IE
sZtXPgaMM3TQoUM/9xLxyC4MfVnj11CISkE5l2cQFIfH382p74Jy24J2Cte0rhfzQ6NQ+mTRjzZq
ezhnX6lMsA6qZMcNXDUSjhw26aBitTEwbBbaNISuyAC9ZUtNpnSIPoV9p4w57Bd8o7k5xUNRt1R8
0Slg6L8rieFGpP/7I4NVPk6q6lCEFbh1UMmq48DBkWv+fOdOmtJ28Vp6mtxxqhpSI4V9RHdfB9Mk
UsgCUDDIxhouiBn/BR7VinMQjsbpsb1yiIqv/AkOOWKndLsS9MiiYSP4I+YVZ62u8ovHzu7j0kWT
DXxzQeUMLtO8HL0rRYhmrV8Uir/2nCyF6GEDyNgdqDJcACD/sG6AOJpChTIIeZi1H79zH3Oc9XQV
UwzJ0H13f//8TeH0iff+JYp7ExIhb5plBbc4kt14W4RNswLVPg06jeiOnXUEYiZsVGH9bEJ9kIJi
NXZeA8jI6OozZDjShUHwPxKEMwan2NsO9YpL2wLGfpQLgEls1nI21TO81+GhvenoOQ+q1QxSjw08
dtEDT0BJw2m0+ktBPKyqK1EPmodEp+uquKFUniyVYEmLu7wnhWoWY/0ABO74KiHJv9ysE9olQKTw
4wjGHi3AJLWeJA21qE570Uxj2lGRJMlGs8piN9I0J1DMPN8W8TRD5P3Qp1ezj6yYeGAEmvEeU8Sh
X307m1KGIMLSpGcJk3aYT7x+6Dby6EHM1Jj4htzp1NjbMOMa+KBDN/cS7iiFAgOhfSmMkZ8kuWgx
gH2uanjhSXfWmAGtobN3KFIaThMZBQXoYG9swmAD4W7dY5uoR5FHb/eURCEt/05M0dQjkp/yJNVK
n36AVuBm5RpF2goQoIinRbJo+VPlh7cqvnYuDwN8q/ARvsCjTdMT0vexQuhfrTuSH8on8mmkFY+Y
C7YyZGIfSwlAfEN/loW+f3A+OmKvOaM7fuHGY3DyQon3GH2S4tjtETkCe4JW60zKipaxU6Ms586x
iQulf5ZNAQdQZ6JHjvyg3fMgTFfPHXKjEqY0mNdGuF/94UgKhsi91qRieaurzRU9iMqBmuUCMV/U
Dt2CGifoVuTO0VWeMOg0liPxg0ZSqGxw4e3I6k4ZiUepaXrCoBRMtHH45gNLfpNvxEFNDA7+3Jvz
gsf4BFtkIcM7YQaeASja+VqV5Rggcsu7qcgMAGvVsEQjzohhkAzAyhr1/LnKnJ3yz5YDfeOFL+hl
9Y990hr998mZNbHzSJm+vvN28H0odHEinvpfkVprpDVaw2d5IH6AShnHKBq08hnE8KKw4Aybw+DY
TKN8sq/n6W+8PfwyzyyyfSCGbXQSloND+RXbKjx7qtEUIR1OckrTuMhomtRZp2MvzfTaynfOEqLM
VlEEQzyamJFla15teC6QHJ4cRk0cxVzgp9gIBjD/qM4JhgQWHbb2Rzr6OIXJCO6hgOki5bynjr1U
t7mgQWwcDkeY/6MB6JuT5UQchF5GyRcIiF4CHvjfML36yG6fvDOHiTbyH36LubZsaJqKK02j8UHb
E2XJGYMjlRjgGcOOjF4js2AR1liND5GG7TmiyWU+/inXh22e2A94qhtj3aoqlG1yUSM0gyeuRH9A
0rOs0s3QDIRm3oe/HvoFEr7CNGj+/LrGlBi77QvHRUzvnLjq/i+y0dzznRUwV9WPeNmQhGh2wnMC
DbDw8ICtG50PJBG8OQdmqVJKzN2YjIZ6GdeV5JYNtf72HZAjl4kc/d7Ye1+SLPd6EqQjD53u/w8X
dnyLYo+Qh4mwvhqUGxaPyCLwBFfTi0sRFjDT52M6LBZ1zLf07kVVGhm0RKQA5nB1lVsvN/4THRJ8
AFwwhuTDe+B/pEMTfcQeDufzf4ahWQwOAip+dKfTU8tuOn7RjQgWFkDAQbvKoF2LSuj7AsaBZ2gG
/iscsN3bWqghdHe5N5STun132zTSoAqsFszTcrNuWWSvWvDhzo7x4PZ9P6GCrMXsN0gYOOPScGvh
s1aX2BdMTvCIDxiCJwmNM7ZuzZ/3BzEUwToGwmXUXUSB1ZBeFQ/Vvovag0lJFMDNbsuNKtfeYWzb
Ywvz+TCvKI5BY6iddwFj6Pn7UGjCXtQNsJoqa7XBPtCYlh0iJdy42pke1j+FTsbDEdZpavxxmzzm
NbWmGsSYGLLHRyVKSyy6iZsYotVuoCEFj+hSJtYYYDhc+8bq7M7SEHkDybBG7B4XXu0qJjImYV//
viuND4b76ZJjbu7JnhgU0TYOr8maX1iMosIA9Cq4N4mt7cIlg8SdAl9Qp8UECzp/lRGddZO8qPbv
SOQX+ttX7wLJETmXVL9ekEl/w5d9ThxPN3yB/wqSpNOv3ta6jyGTwe2aWF8B4mWFFJmuj54Y58co
b5iA89puzlFyxoSD29AUr9H+QwadnZ4QNtdfsV677eaB5tMqTmmgvaUMuL/aBDWvkaEMoRtND9K2
ArEnHYfHWtsKwQsQI8mT6Ps51rFU0Xh4wJq3sORwAm/mZVblJQ6s6U+TcXfCCnnxLYaqckX5nwJI
v2MjOUae9ggt2g9VKCJd+1grboPbOCtffeX0uLB6U4AixAvDmSlynltmldnh38e/dbEksCZCTUkS
8xJbORgGo+7Wmm3fFXyHpaLXpTZixkMCsi3/i8pQwlIIRGxQm+qo7m4u4jEl1rTOm0TWc0ZhStyQ
AmNG61uq0Sq2bJxRb//dfj/knNb9RNJwdyTFVn2ybftFzbO9DsOpJeHkFajsH3BvxfmIf3K6tCwa
TdboLtDzMqGa4XNUlHAbWT5/ZGAHc/5QKC6X1specn8j7Lo70Qst2nXMck80pTt1OL/W+TCBLBr7
cmkxhD5NWhoaUQ3EJuWgrMlzWExhMwbHvQUmEfUxhDmPSqp9zSObQDTtfbJer3oDAWtQEtG0yssK
xBxzSGsQmQqtPq/zu0zmvZEY2BxmDQgbRd677NDhRKBINsXdOM4Rtr9u/d2WU+Oo/NEqcOyj6h4j
M3uEWuLtX46p+VECALt9ck+cNdLN6laqOko6FXoukxbMNAAFOak50gTfIUs0GX8heLt7RWaIr89f
6mDkLQAsxUHcnZ2gZf4Fz8IWbac/N9IEDeS2W1/Iwl4ZxLTwgfR0xGzj/Y8ZJ8xULvg6cbB5A8lV
SCf3mVEwhNqGirDg4uvNl6ZxCtAZfYULgba7HRU4lrBhQ4yeLvKTxTIaqdPQenzUmhxCs5Kseb82
Ez5afCamoKH4Ht2VpY1BxZ9noUd2a7dAS1jnHD9fN2AU5Xblwp3amBcPmX7PppwdbeRQAsHOrPH/
vwag10JIkKAG3jERA570K65DoBTIL0OfHAaN1gQcLFhGJ5DIO1QibjX3KnYvlKt1Q3+sqXA/JlvW
FgJ7jpBKML1qSs2zExn8OYmQ3Uljjjnn6KF30ugK1cQGHxCub4CwJiicPi/aVB1kK5njIYILJCWT
MhDXGdS8UgBKbGGH4i6eSQsNCmw3ZRp10wmGN7AbQIWzTWmu3SdtwuAdfJEcmkIZ+8k8FGHknmXm
5dZK2uP1aCYpZWHojc/yQLAllbFT5UR0rFiVgVyI8ESml3aKn4nsXZx8jJ1XZxuCvG0s1pk+KtkQ
DX6WYqAZr4yDpXyANrZaMv6D4Sge5mR7Psssr+L91fMHX2jVk3uBDump/vRkamUX/aMM1RGEQPIQ
HCzkPCnTEfyV8uDaG81s0LelMbcvx4cSUdUq/HCKwprNPQFL52dt6oQe68ZviITueg+LtQUc+H+P
bIku2LR7/Knh4LGBnC9No4PpNlUp73mU3QIVbXL9TEWJTiYOOyfjcokEC4pTUD/vknpGmIaQ+KFq
V2cqA0TKIko7JkbO62FXLDUx1qN1Wz4xlPOVYl5j+UNmTpCRKueJMgIrM7untpllV6CzC5vU9ZWC
z3G5sIjsSd9Q5Z+n8u7MdOjQbHbkvPncejXh0mAbm0kstzrNT6i7EOz0QxxNfZsaqEO7D3zcGvHh
Bo2eY/0BRKATsLBq5D93ESBBr7GGwPY3oDqnosfIzJWoaqTFcNKo7UE4wEYB7egF6HcCI0HTPwzI
zcLq3ovM0Yh03/w32sB6e1jaw/rSRfeLcBGxV5PzXE5bBC7BZKwqdnAcVp+o37tqvCaWUk/Eem+Z
7xYuyv2mgrhMBTMpXwYsQG8TpNewTpB+M18RetsoXEUmdHp5q+VvbKnssM2yyCl7kWaB3oeD1s1B
CIXv4FWIpPqWq9tfSaedOXa7a5TOKDgp+HDeZi5dZB3XMn/MrDgVMVReG8hMMW6tXbMpIhwGhR7s
K2uQjTbytcENDOOWtdeyin1KbaYoDKSnhI1iBta40bCmiv5rTFMFsylzsn/LSCN7PJzxYDBWDa2j
FUFe/WqsrxvhevJeKSkI49SltfVK/BpArEXJ+CH9w/rzAQw5eIapt8NwtsVKB82tWw+UKjphj0sM
JaQm1AWgmo6LWJ2jzYV+lgS4HYfjS82sVQaGTdK3EebIxX9+mOoSe5qF0HUYVITwAQr5BbezTuPs
D7rHHruxO9eqhG8BZWw5T4oYqBj4EBAZefoILGJHZVWMtwiC1joOcp3DEVSpF8Ke/l6iRA8YBUbU
wcDVhFv8fQHyXjpvCG/Mo0v505iuT1EaGgEMMd3jXgfa09CBEiXApnLmRJkWu3lDDluLfT2dct3T
m/SKIC36PcyPwJpKfmWi5N3th4Os2dK3IODhmH7B/967o5NcyH/yFcr6YDgkQKLTuJzuGK0auNHU
+gi5TWVFrWUUZYH3eWOkhjpmVqIgjIyAS2bl4kSZWUe9MUULSMhAl1O+gM0mlSX8RuQPzPeDcOHw
JQmIOKtOONuM3mEbr4wJtOYtXUytHt/c7RQNJQg1AmKPLDyN8PgYNWumK+ryHQE3zvTdQxW6yTfV
ZNA7wxKcxhRaiIRl+o7VI+CXhkuyjgduCn8mSsnEPjLVCKCq0GaNAirkHmVZ7k+qESCPgnc+lbBR
z512I1naW+3/9pjyWZUdQ0SYIDnBtGljoRgQbw+PfBPr17kEnlPXxL2c9FdjYtIHKnDZZwO+wCW+
28WmLGx5IdrhnMTmfQduAOsmV2NUPXJ/mtkFpTVdEPdP/DcE1zmxr+TBpKrFySXFYbHNjRsHuyfp
VFFqb9IZal6o/Q9CDjJrrQPlueT6JP6PzVy7IpxFAELEHxOUSYGHzvF6/l8wbS+/7foT8lJhn+a4
ZHYS3wbT7RiQLCFshzpGx7Cfn35gByezneKyCvwtQAFExCY1TTmTCJr3JTcbgI2odRxAPMPIy/yJ
80Zq/AUR2a5cvVSD4jo63+rAqs71zX/IeOahgi47HUKv4DIdKzZps7RxbLNZm2tNxkB+w7yj19GH
qU8QLXjtxDyQViWkRMXO0iPO6LN/xnuY0Bps/IvDwpOmczX7cdoxEJF2EtYeKcfoNFjaOqVOuQlF
i27nqViFGBNQl/DsJhwENbXEN2gR+tsEM+v+X/k/D/l2ZBhc+gbeHT4LvNhahI95qCcsyBeASoZA
qAZr9dXS7aG7sQ0N/cx1aDmSVDuyy4TlJoY5k649QT5o9wr6LlBbc1l5ELaB/+ly/W3NLYXN0GW8
pP4+642NSlzjQ8JqExOqSL5IvWR0Nrsuk3JOgAov9gOwCW4oCY34ztuV1iBqNAgK9Btd4fZYq9Sh
9IRB88inihPDV7DAtNh0ICqmV8e2ge+Lnabt9YNNz2OjErQCet/S7Z5E8SjjC1s/4tx6ZZiqqNc9
Ws6jR4zkg+mUSEpL+lvWiGy5ehrZ2ut7I67YPUEQutDAnvB/UwG1n6bXEFG76eWx8uBWgaGldZNV
GbUr9+/KcvaAQmKLIDa1pp8WCr+6HXug6Risv1NYTibfFUBN42yG3/ThAhFlbOhg7BPVIScOd311
GJkZHex3brXTQhoeIcLFjJkeKcyf+p/JClTk0RMxvNAudRcPJPJj2TM4x/dC2byM54eb6jBe/2sk
Ro9lZ8k6YTekO73yjvl1rFVb0USKUN15cORUqhexq3APFwlewK1B+I4SL6wXNpCryrNDkpjHXg6C
rIVDPvy7tR3VGe9Gd4w/Z9xgcNvb0vYSxr00/jzI54j4rQxBHhMgU59PaIQ6HmPQKoClgtlvCi7J
T/VkIQmmBsHG0RQ1UdTUMYa3WrYuujI/0F6tiA5RLJQdis1JStUkCGzrFIj4TjP4d62LHslcIkVP
0px/Utg5ur1rYfpwkeX8tm/PAzJs7YrrrMP6W4V1luukNEXBbIbI36qoDHxoESk3EysD1UDd9cMK
vBddn/X4kb/aPmswDdVPNtoXBTUJKJejNb9mQf0ri5ivB76LprGLQALVWF40PSS/tsP5VWcbytNB
Q8V1xoJ4X0gR5l9rgtSvjP3KLdo0bAUqLtMrud3decKbQTdwrc7iPweXSEnQM1IJ2V6sp5S7aaP4
oq29apqZz0slVpWxXyknaCYbDmDC/pWN/psE8vJZ6F8UFWUXhKgOA8nsIWpKkXOe2w3ywbwQLBd+
lr9zuVVlarZdR3O8fYsdpQrw0K0ifKRma5L3kk/9ykLeW2uf/U7Zs8siM+fFhQnnScHbyHaRte93
myDuGfyOhCTG3dTWfnvvyLSBF6WPgbKVA6lxsw/l5n00imVDEsBfTmJNydqb4ewlnbnFJwcTYEgQ
S56kOlTB+/f8buEvYH3XI7IFK4sENcs+Uks0e2SjNXh19HW0n42Z5k19TIs7iWEWFvz+dV5FbRVB
xL1XdtCOgRgnyK4hdWahDs1oHuWpFQlFcWEs+Jl42qSx2zsip03WuQOZLFXfLE22if3Vbd/JwWZ2
8Fdpow6tvHj5GxlFkW2kAl/nu8Wq2vue0esOZabX69K0Cfg9OUKlm4P/dRJE46tmsRmW7ZEAvrCD
pi54aRp7Mec/IcUlhnz5k7sya89vdxT75mffyjkjsbAhdgQiCMbt9uTNsbz8VFR0H8oUOiduimsD
hO8Z2Zg+fZoEXH0wjzihegSTWTlGtCt3TAex5TXRgf+ujMJVRgY4ecYxVhETLPKLknJsgWc/vRXZ
4PU/lQY2U7p9oihRIALuopUBgHtAxTFGpZVVfr+QBgq2ZloQUMJisDl2EqDGF/xsybZn9XFR82dJ
go/DWx6/KPhTuK0ODBxVEhfmmNjoLaP1NUF///pfVTaPMuY8WxrywAmNsVFLgND43kqZjuhkt+eq
so/qiLQsxIuQVe5pTOa5E8EDwrSptkMC/8/raYzmEJB3V4c6kCHU+7OXVEc0RT3oBFBymfeKHtPP
BBc3GOGxHTDcbzj0B09cOeJGqYdDYj4/ndj91RRWAnoW3Qj5XsYFd2RFc7U/TzWatujtYlp1u/0J
PWv8iHKJqCmjPHUnY9NG7Ry96UWM54pyasBC+YCn80wWVtrH6rK/4p5oljr4fBqJWZ/3/KOZJrKK
V8w8ca5vVfwoymEW7ysx2Lx96zz7lhAaU6F4V523287WHDcRuiVcMt1/Uk7+gnwCC/Y60OsDPe7G
iNHnoW6HUR8pgJqCH28o0GO7lCans8hnXMP0n47VspiOpThYup1U3qgHy72/tPbAmoVI2FFmR/dY
ZLxVrbIuoCV0JHfj3827r5lNMEwnov5y+2xFP5haaumWT5rGV/ArHXDJK7ZVEtZFXcrTnmfo2qrw
4dIZ0IrmHcCuUeaR71MSaEWx5OclE9LyOkDd9wBUcHRSCDoVgXxWW+Yd72vJH3O/68uzbETODQFu
3gYBITT8j3OQPIADR+3b7IuA1DEpNjjKY0uDfm1mB3BiuMkb2Jwsr4jWwhz13+UxH+mQgTqQoP+x
ENFl7EH+jcPltzoNwo0LW41zW9XQ35VljDiY7eCtCoi8Up6gfP8ud3iUe5VOGutZKF989YGxy1FX
iZNNGXr08MoqH7qmeyGgnAza52zxyMto5q5vUstjbwOfvvrgUpCUn7KY17micTfxhkgYG5SgOt/g
EqQtuMtrYJP1lnYI6pAMW3AclNIDddAyl8iR9qJIlLh8dcCqaIaVHzkCDaGfikHELpxYIoPRBhWS
9QHduBCsAm7/F9f5lx/RB43yIeiLxaccPZMhAsXyAdVuf3TygThN8oMRwDxSvYEhrq9SM8b9YhB3
xnZF2vNclVy5bzweZ/c20C7KRyrDCFlqPJYiJW4oN/a8H8nPC0smoUNA64fy/yaubERT+PvZWGgs
gBm3eT/u+gGSyA4bGYBmYJrmDqTFoic/IIr8QVreUhiC14xdWT0sIvucnJcjatLJVGz/iPoo/jo8
x6ZtTdAAlXbuy1hVFWjyKAu0+T1pkNFEuO8MldXTjFwaD/TTXawrxqZh693PPZ9bB5OdSaKNirxs
9q16dIrCmwwJubFHixFEbnf4M4iKeIcltbgywtvDr7S12VnlncLFtiD84FnHZJgu26pqDprVSWPS
8V/tJi81wL49pCsFIPHh4tx38NMumwMlojoOjdjzbmcfXLHTraGukrrd+NBY8Wahyo2sNJGR6UaR
Jdhv6sWxNuNoKFS9OuZdl3TdIUUnahsLuEo0t+JKKetVbzIK+pXm1KcH/nF7TkqJnGhN9VzXSw1P
gW7g54TbsyprfVe7TDXBj+jLL3TLOoo50/zV8monwp18NlJ8AfCNIAqbTm+PRbptdJbp0F5VxegW
SW5GbARoNx0BoeprRxg3dWwlKxpA7UfxRyXI+Ro98sa8LdZNcdaF7iJdDb4oiGsR5V7Mun5orrBl
ThzDhlQQNbLXKAlS4P2A4nLaY89lZJNn0kqaD1F1dpYZx31RuKVHhI1Kp1eK+h6Eeu9gU3blQixr
oRorgnZIIFrQrXNY4RdL84MQxYSDAzKF8B/S9eyfF/muVRu2Fppt9WScrSzf48hr86XK/1Ul1bi7
5CixHeR/hoNsKQFSzpGCvmIkfnc8QWsQEba1W4RPYxgLHjf7rsJCsMDz+hq3GaqDuK1Qszq+M7HQ
ciT74tLf/8Ulbu6IVQSSeESyGYPsWNKGmBIZH8LWxXHiaCmHAbwTSRPQeAILJh2hSz7hdX3R4Mdq
EmGAz7e7sKI8JZacYPEAZ9YweEwxz6/GTjS2zt0eX7/8rx1FIdEwx1K1DEYGbq5fu4mvGnHjh214
y0PjBCHJCCg4YWbQAu5kpjxlN6wUoSVbAPuh9adZVM+i1CrCXczBM8sN4VEf+oXieJXljscAgB51
kTQzMIprG/UN7BubcSJd+42x/AH4XKy4PQe2Xf+MJ3GaY7BJm+q7IkZF/p9tGwNu9FAF5qgmGImi
2RT7lTqlZGVgs8VNtfGtFzET9gr7J8fCYZjq+CuauiiVUPJlIZHBg1VwksvBYc6e2e+3gpv1Q4zt
HT/4dWpk8Q7CRqOW1NpUcXgnePrBgGqFkqv6PVbOXPY3D+6mO1rt4XXNXoy08ZVchLdrBqoC5fOp
jvoRuKxTJhPCORcFJgPqvsYdDCI8DMzv0h3IQmcisebVgIW+wL7rCQ7/T9KL8e9WM4N8FPb9asC2
mN8g+QPkD7kX40YXNwX/6NBi3sakd924ycXgotJEFoqQUp8eRtW/WKXNqcr+sBY+1lgzU77N4GYG
b83dW7j6W+WEa/6j4lO93geuf/rUXLSKdeGfNmMxzAudB2bbaC5ycQG5CQ5wdv4DnvWWr40/26zw
rf6DWNsmDY0Ip/RcCYx6fWcZrG4u0+G3lQM7TeYQwy/20I0vlKcaTBh8MgtuEjV5+GrRpY8p+BSj
qxiDoVyxiJyls9y8wObIBTKDz6bz0p6thAQq1HmH6MnkFynVJw1J9alzcebDCsH/J0lNNO69iRpk
h4Z/+7bx5VEBsqH9FkXv67ojveRsnBxPxBaS7QJKcQC2n4fsDZ1b+WbXcpmQ98G3Qu7b0NgrCc6H
xmSa+mk9szdTkIP0TAKMeFFRxXL/DPVho+Zcb2+7zYposPdAO+/Pcu8QJRezCCBXbJfBo9JnKgtu
M5QdD5T3slAgUHmagUTjtUyfxc8Lm25oO7ZX0qpH+fhXnUBs0/PQq5uKyneylQqhj/te7V3KLb7N
82EaHtvrkROBQGoREKjXUv/gll4Sd5tLPuI6XZ48PjkVFDlUsEzFIaIp3mGfCPOhAe/j/6cXfa0P
K9znpLsBUZ7W/qpvpDFkSdeCGplsukJNBLpY918Z/uKV1Kz9YHQF/Y7c5laLL6OYpophmd7cRgms
4LfqSaAZqq9F1IzlmMBYeeXHMyC+NR2sqe5o33p/io9o/vJjYFl/5jLwCDHffIQnSWLVlRy3xDjD
mzep1fsGjtWP/4NGgY0MhnNnWRbkDshuT6XAcmdaerDb/DeOyd/xCzSyt2oftTY7Ud6Oen+IaC13
5uB5NTnHWjTTRKLfNHBLQ06j0m3Div2FQe9CbQKuum6sAkXd9Jvs2TfH2nbxuBcpoSdvjnXI2ahL
+eNyNfGXRgSU6+rGEi6933x7/objY7FKNt9xYqA3yyMyWqR33tTtP8wwN+vufnjYJMAQzYqhklyU
pDjVhIahO1JSiExC2JEqlC32WC9aL/Q0lgz9i+vW2ksT0/VWLOlsovpAVxbeNkbSl0ABSkOzRQ/K
h3lE8OCA+0cFKd4jfzKyayJ5lrTAt/eYLoOtr02ToMjO8iGZLlDQgYB94zsUJTb8Lb9YmNLSDErD
tYhw/7T7y1G0RvL5+DI5FELiYUHUmyxQGKP+8TfwzOmPMZtvvA+aGTEQhKahug5zw8nT5eNFQXk5
xOnMHqi8RcJX6R1gArUu8iP1Xn8i06RhGlmnfzxMbbAsfJva9Wl9YRcSa7YPndfeGul+vS3Tk6IY
sW76YkKkkQ7NR6Td0Cey4i0P8+I6VbpLzcELhp63f4GbVjdoTI0rEXGfTIeWMCbNn6lK5ecbJvRQ
DQ7djKPrQf4GwiFw94YirvZztAxe+OIHXOEv4o0s5wgFr3dJDc+QO7is5OdKGFu258PApjUjw9za
9xmezN90fvfibc25DPGECdveZrlI+SizJgDlxjm04WsM2hHQCV/dbtc/Oztn+yhiH+W4MnnP4IpX
ab0nBLBPiySH7UaIzM7KzgKQ2vRPTf864NMrKmAJjznbIQvm6sU0rtvFK6mK9HdgoSIYU7FRHBqE
C/PNMJilzvNNXbd9VczQUMzihfSBgdB1lVXoLhw6bFazgjYIElrnuoOF9uibyPtV9mKAiRiCnidq
pJiwX2ELD9tUeauFxmK+T5sSfBOFPu/gl5Ew6yTcBHtc1N3FakL9ztxlF/mkpLguF/V1r3KnN9Pz
a19CspTR9MzJjxTrbmK0k7e3eXntHO5qM57BRWTLvBlLLZxh1Dp13CJ81cZB3L5gix0qmVVOnP29
W2berttv9oiGCtGibsFcQNM7pJRdEPnQRel+hJD6r0iOubkEmLW0IIE3gLWFh1r6tPprUZFhJ0MX
bw+Nvzj0sW3mQdRporYnPeVGwRNIY3mbPT44ywahzdNihRGgBOpjn/NeAfsU19OqUCTTJ085UUp1
D9lZulpS4DfEAryyUFjpEcTv1s2JShCoCGOPrfa58lYwvE7CmcT5pk+t1xIAHWOWSSXCDA56VfN6
+rNkLluG/mwc2ycss1CwLpfMFaETwqULW8htc33v7eAJLnciBOC9SDJAnEAISqaYT3JsE4jfuUih
vV7hTjoiMDWCTib2tA9NJBrjN29m69r3QL5mRR5J6oooZPWELnuzuYy0qjBc9DysDyChgbQj5DQP
lUuFopHsbX6D1dERtwGVHjYtqjaUGF3X1C0+E3RifRPGtT4FtmIp6QedKFlIV8/AIrcQ1Se1Jsym
FoDvXfvZ++QOZANzxw5bSTNu5liyhkgvtPVYHqTc4JUwzPOKpRSEpooVl6KwmeDcwhcLbw8MPvwV
6+m/0nl/GeP9zyKStj+s08tNJxKZ9kk5fD+uVDYc+/IGdmpp4puwons6C+9fpCF+9idEC8N7GpgJ
tu2nRsZCrITR6kgcVgOV+qLQoZiSq+jNP0Hdt9zaNWT1B6Qt+F1qsEmf98Kls3XZyXH6i6c3uZWM
7O0lnsNYJhS8iTDXreMmcCza4xSn8GGCy+zQamkZcbmYHLJZ1nUTq+FL4ej4am+j/8jg9VmRjVMM
ZIQnkLDRobwqcYY3yejzwvbXTThLIHI5tjTI4zmAk48hnSLT5xakFU6UNse98EmaYf8S8u4KTyAn
R7SFjdoTRoTnVFlRsQEFVx2Vv4Mpozm/RgGj803Z43O3P0bC5/cBbip6I3PoQ0SSbX2wtHBD6g2Z
8KzN6MFFg7TNeeKITEdAl5QV38oAgsuT9qxh3iZq8hbkXkeAALsdF/kA527oeGA1oioI1dLZajF7
yq4fgCeRFxNVJv6vJNjqzhtj5mkXoim9asdO0g7ybKowtlwLMmy3TQUXZlAqAxTcTPKvVwoJxXod
XUo/34cZzkLvSgLlb72QxcL+ED6XJfhTNFd1c8r253l2B1Tp4jAqaUSEncJJTvCOHFZBZElD7LSJ
zyRTBux2KyOzxMY9PyTmYbwv7q5FNPvolNIG3cbZnFMnJKwK1HWoOugvw+H+x4WvkdePHjfJXgGX
rCVSNHqHCcEvNCB8IVciJ6CAbBY/MWlftwX2ifIwJFmRv2I0sQOO9oyFgCt6EUQHrcXAehUZKvzE
g1KpF3ty++uH8cPoRALSgurpGXxQ+UdYgrhzMYrfw0CVNqEXU7M1AN8kOoeqUSaxDRdMgEz3LC0P
i5wJAqXqrmm+Ovq15GcQbGQBoRwYpTv5lDF+ETchibm+lBLGVzkeJebcZw2tLYiNyADb1tKhO+Zz
rDtBx071oCs4L5r8rvV+OLmbsZNvYwidzFgz4XFsrjZAJx8vAI/pD09mhs4inzLOaztmi3rAeoQs
Dl9UlS0Yenr+hVN7C3kwUYq9FTZ2E9Ntj8PzvlXQpAsTYkIfYhvhcAAnaCgYvqso6Wmny5FGci74
IKk1vmdXECApTdrk2kFtYalISVd7Ix2YVGONN65c1F/64wCHDdVZL2UqT1LwFGOoFd3ggQ/w2wfE
rUgzxX0Ajqv/jCNel5c/Q9ReBRXCaZdBoqh6wU3pCi68jEA8pIuO4c5t2+felPMPZSeJlDW/flG8
KzsYj3CZe2E6HLde3/tSmZur8e3Csr2p4ib6dWn7ixHUBVkXYhwPUPo2WjrvalH5pBiVynYSzHqo
9W+m4IKyckyQIuk4D7PSXQXHc7HmCeDCpCYaQw1aiOEVhNfYGZtqDjHAv9yn+Wf6R4WULN7Lo1/b
ybAmtTjyUp1O5rHvOUX1keaBwpLhK35LFToOqkDa2lUUOk6gC5oiq7BpaAU6GDh6wuYhxBwRI/kK
5d/SRKssXmviKkFwCFeXwLO7bgKbuE+drUk5xjHvKbcgzi0Zxi1bwVtCSJPcd6J613z13St/hFei
g8dI7aiqPV/pDvmbprBQcNmoWndP9bq1gYfwVWWkBkt5Vvtmfoq/InCjtPkDbQpV90gBGr76ymU9
VAxoygHget92yLAivqtTiSesuSW3e/g8EwOAb+dhdVYtioo5Q/tytSRWhbAOBoT6KznuCQgbXJxQ
tynDY50r3bLzox+2YbvtgSbN8gp4ktRbRuE5b9HuWN6T44AKZHrAYdHlUvpTa5O6IHnYYPfHQzp+
TVdWjI7RzmlO3ro3G6WzSe7W5IvE1ULUUfgzGu3Zi5u4E5+7ZFn0AAP9htY3uXEErUlAI5D0G9fk
w9H5SEUOnY8kAsQXCEyKcYFF0lhO5XdBC2p+841uqEeNE1251r0v4u1kgKvBkZ0QdTXgIvbxt0Q6
zaFZ0ZSPIElXvaVuRuLyjhrLzlo+EEIy8nwtMULA1CC/JyRWaKT4LAsRuUspqHiteL/meurpd66F
0tKRp1q+R/p/mKOnhPMczaPiN6NwRju1Est3QTXRD+5zW6C/5FNfQrNTnrsPS+Y7aMNIDz1lJck6
pIzLPwvVlExjWu69lNjLF56unREAREfJ3ks8LjIU4b7GQ538K0ti2fvwI/fop5hCPc7HMe8tAaar
tTxktTpQlH4g/Cv9EeB/k+aF1TOtlreLAQk27NcFQon8Z3THLwmdaPKP69lwFPAGljXmKBkGZMj/
gKZxEX0qjt+wPecS1iBBvln3hiN/XrWZWt6rEbGXX4v1NTHUwvV9y12M4HI0EXI9sm29W6XOsGzi
BTFYMc0TUXf3dQtrnVY/w3MSWwTrJHG6hoScGnMBhk1UKbJxQvmCpaZqoZB+8Ud8ZVWtotBFtywR
6ovpor3iSWrSp8wgRotlrbd5S3N57BygDg/X3XdUKtH3mj3tN4IRlWLhWwQBAceG4dX6GwCUchfg
KU2o70CMJ8mjDUKUXbfMwq5sggHQK2f6zdl7vWHlkUyZsGWngEymF4PEA5E+u+jD7oFUU6LmNTRd
sqglvgORcpy7j2sjmnMEcNflwnCMb9i1eznUcDEfyoxtXRbF2+Rj0fTTCdDKTjG6sZFF5c6iJpx6
aFcSEF1gZBEzVXgW0mhsNkd4Yf59Gc1nBo7pFDmrbIV0yTa7o2ymZ7BHcklffE6DaK/k6wRHei/E
dfNi7AsD4uA19DwR8KrbtFmf1aA6n9XrtIpqWYm4bkLYG86dlvmUGRUrDC1nBaMMqvPSB2LucSZ/
qs0M+PLuR4huyQYMANBnX4q8rIvp9PIbMqtqbSaE9gYUAqVyGqRz0fY4XLdKYeWDo023ceISZAQ6
r+i6zcgQLTXjgkELcvjGbtSc0KtB3+CwJ8Jf+XfHz52zweYQU+S/13n+57o64L0ZHKSyObMw08HP
gRM0L9ncMnxoCVepe7HTDnxoPljEKjcobHCnKRUEqCoaUX/czLT8nAgrrZMqvzcbFLfTw7XGRR3Q
Pf8o1xFDuJDUEnUsRl77B5j2fzjND1eGFcnJboUCYTDSsn0TdAe+oaOAOhsYbKNT0/h+7A9n4G0n
xsIJyV6lczbpq0PIbIyI3m5mMw2zCPAlqg1DqxRwSpoJoNGjdp3zA0t1q1PZC0gPWnbLKkHtyrfo
dG1of+25kBgnKH6JlZNSdI0pEFBfj6n8TRCvkCPex7lgX7hRFrQRax8m2gAnF2AqgfCOTRT99qNf
ucgVFvbgGJ+QP9ZNR4pCFVFkLUIg9d8+UcZMQPnRRxuauuqdgwIo6NUsqJE8xzNJaLF1nlQ/DY8m
SG5BI4tVvmdSXjqURmJfALhJVPmEOB/jwieoo3fc8V4IVFk8w9gVMRxVoXrneEJrr4QlLX9iaFZX
YrJi4mHv19Zu6PihjqzqJ2gkpm9d2Xf/kYmOmYe60iwg5dB5K//xjlyAo8t57Cj7oC+f4Cg9nHZs
xLQv3sz2io7kujRUCBSupPysWqlTs/vM1Saxtl73U/C0ZWdFxjsfelNDF1m/DDK1BC1dc/yXV1p2
vZZbIoYEeCTVuef9HnTEwy2ldyfVPyftCV6Td9V30hIVViJGgX+lYFFS/LjRDDIdQf8FfTsiPw4w
7rFoK+R6PiFOEIs7jlgql5j4VSU2bxdLTYn/+5T3QX5iBvNDNKzXFfXo0R+WYDXsnPT1jqvv9TF2
LFpUh4iDj+6NxMtZB8zq6WdFEpslk9R6BSJE3AEYFqFCn/1LoiPCGmgRwNARZLJD1bVjthAe7hFJ
XGLyFyC43znN68opknx/9eNMdovTtil6pC4IqkP458DSFSM1yrESjKV8+PcKzye1yGk+Gfk783X2
AxP8nHdu692PT0edFl6h7t8K8dSgKLJFwOAR7WINNif8gAbzT+hMeKcohjMuvp0eDnWaDBJ78dRM
6P07zbeWo2ufXoQ292SnDP/bn42Tl42FgkiSSXpTJArqATaiEqztETo7PFG7rKSTf+YW0NTOn9bK
RUZoBvki9JHbW15Wd1Zts9y+2cQUz+c10pZebcQXUN3nrHBSYmTbOh5qbhralasUbwkObZ0FlNFA
mISGq/LHOmw5CKbXNZiQ5EKuOk/E/Lc2ZtpN0PsIMaN4nOeHdZ0UwepJVLAfNQaYp9uHZ2QlJBnH
PCmcf31z9V1MglGgC3jq8o7Fcw84wluRiAb6LH/3CL9RYYYB+4j86hiFFoT+tU9Qby/QOVYxGB18
ZhhDMHS2li6CdUPvubcIEfvC3c4MlU+s/XPBOtmJwo9Xrk/SjDx3oiK3ByFqA4iX3FURv68fNs65
vaYNFJh/beJnMBr5YlwqqUKIRbQPdiU5OW9/+GAp9Lwe3woShT0SDcud01QDDS6nHFWhLfK/JZ4m
2yid5PdI1F7Sf/ygSNeZ9Al9gxMwS1tjXuJoKvm4+v5BfcMa76DwVkUMmZki6nB/B/ziVHPOBvFl
0NpntJgmNVO0NlAnW+z6GkyGkwxr/HJYg+vF3CjDCFjhVPk1w4ON9CDKWuth4DeIjXufCf3dnsYf
pcJQdILP7l0WI77vZJuG7veLZUwu4LBRVUsBF21Ms8lValJAFxodXvejXCY+YJHd78n9AUwI0YNK
bKWy85gu+kVp4SFGvtT3ZF3J2nzvSpCyIl6oLe7BrNhUqvvJbb386zsOOGFV0ZCRWa3DdYRTaP3J
HOVguXrW9i82hqqzKkeWTCY02DobB2WSV2Ob6rXzR9rN8xx/lUfULwMlFaj/FI/8NYHmTYBg2p2X
sgy314BWfWEvMhQAtUJFt9alOS9zP+h9ByOwF1ecLUww+wWC0rGQLnonMoE+DNVKyNIX+nyZpu6c
4mKWrZCm+JiZDa3LcBf8ZNzDKBOlGXMbXauuKpCxf7KyWAKizAde12hykRJm9Y0s6J5sJDjj8Mlu
CCZ98veRmEqr1hWofplbhz6rwuhTXH7JLgittoXKDFZe5U3ngxRBUeRXb1ju2EdvdPlRSDZhaELF
q8FLADA1rVltCD261W2WNRJUtWHDg7KuMtGzUvVmzFC5IGUuP4D3bG5krkRV2jrhNfolUm5S7nzq
h4A+UcBXynXv0+l8VTPS0q6XD5WbgbnIXwU5iUsJsF9CLflk3hml9KVAy0RHwjGzSEVmuwL7GkeJ
DCDHLEWrjvTUvClY/5XifBgB1BpgmhrD8joOwjc/6F2enNnJlPRVSxe6M1QWoLwWG52yO1V55xDl
jxyE99GsnOw0ZflyHhk1lJNFFd5qnsFHGKnavLDBWpjKCPsWxblfZighTtgYOQiq0RHERqT7R4Fo
7S4sN6G9+cr1rwtciodDeHoquaxvgnImE7aa46cb/S4LdxO1UsXaQUXdrGh7Rh/ybzZ5LI0FB0gj
UVbQsK/Bn0erRu2jcpOXNKn6CPJFUaDBqbjlyPhwZmnsaPsZQ6b1+JeYeyVNTPIAVlmKMnkwM4qa
0rB1KUUZ98IeJC1C76j32AbIHPt6uxqjw6nrqk6lOjOdm59PBRlyS2jhXKF5OKmzBzH/Dr1xUD9n
EpNFPlNuqHZVKbz0wd6umCA7nQKDUvpXll7Rth4d+Q7+ZOhuxcydnjYT1Zt48fXRQtGNZTHXLLSL
g+u/Frjs6fFem97lOPAISaQkzhMHvniKpr3KK9jamWm2NuyaRnBtK8Hw414HBEbqPYJVOeZ3aTwe
ySJzkjjAywyDf1rv7KIlBlr1ZdMHVMDuYKkBEtjRrJvJYg/W2ezaffjKGlInEnr0IvqIleBFvBvq
jsJW/E2iToQVgXhS79qqf3LknO6oR/8sqM/VuYXoj06E1YS0QzlmwnZzqzCRfnhbDKZ0SA42EBwb
LAzWafaCGASz9o6X3m2HBF8R1+mFqBZ1X+ZbDMf2WI/EHiIulnVPappcumRUh1Ct9kJNOHA8OahC
upQFdVRFNFgBqZ5NTtbQ2KWUMq3gsSvnso9DMzcyNlh/M/Fx/NNo0nHLlgScykQQ49roNLXbTx0K
iBKFGUzBk4wgjs5NFECshskFEV7ZKtxUsIvJAKLLhXsY/AJ9gSQJLOo2ILaZnvXyRj0hJGGvM9GR
PDFyZ8sU84L0PCXq/iH5y2lIQ2wBVzXtpIlWX9oze5egxspJaLV3cUd1/E2/becLlmZXP5FiFgMs
WqJEZYuaSqAlFbfBup8ZpjLoHAlbxfrw4jvM+tQv7krRStVDW8sulfzQ3jh4YJHfar8SlRM22YTd
6jhoRabMplBLSr8EthDhUsuSvRmqIzzooHhL3vPxuA7PdWQHi5JqKhwE4Z8AhdaSAEQkNAVV90A4
9wl/puocBcKwI2CIMdPw6exV+IdNMgKEK/hBgbqjFUHrWG8i4EZwPKn6sR8Mld/6pA1kQoMCftOK
ka9TpNU2V/vAC8xO9NgeW1Cgc3uwPFbNva//jIwjM1EhKi3AK9MBwn/gnLbxgou0gq8u+8Iksisr
s0NxrqODf2GZESwJEsvAjzM2+dmM53T2JE+OBlkkmG8I4wK+cHnfwKvih8IrsuT8sb62nlEU9+YO
3dfzV46HZUIrvEiqNkm18aWY2We/UWvsOWIA2A9nxfdA4g9VrS5xnboE0GseQBNErJ/lMbDWm+uu
apuMO2ihTpu4DhwKRf+9xXQjyTPglaYFjaxYkApsejEVrRCiumeFRQf9Ir/z74vJ9dFpBD1hn8fl
GtlDzGQ6oMZZK5pd3XBJIomnMQeN4SZVGVnxQMPh6ha/+HmA+kz4Bavcs5xqYvnrWZW7ald1MTLf
yOAJmWYNmEoqN1bGD9rn5noBJI+QSpeCtxenawTT3btmKMLBbzkaCOdMCtiNUlZgoLZUPp3/RftV
jP8kMKdJAfdOjhdu6NCFatRtphIVE3McSwG3S40O9V7sdTQ1erQb9lD2wMLht3PU3RcQJa9i0XRl
8WGlsPfl6O3Z9O4Dt3MBoCpcB9ht6YO4S0aVzQRz7TpIxaT7K5DGT+jtybLOry0s9l3kMn1pUP7U
E16xQQCvriY2nT9LlcAXsLp0kTolMyqe0jhW9UfiExsZIoZdUtaLIUAyKO5aa5/q3z8I2zqzFMYQ
dmtJFoVHz0Qv2O0CQYjdZGtFTyZzXbjPEVv2Hkz5q6JuG/lCoCay7xNPi6arJdeDOxMX0G+wrj+5
3Z243vJ4KHoLcXhtJre+mVsJLkPiiNODtR8fKuH8t37dMzhiTLNSQ7HG3b93cf1lNdOFztN+Suej
AkViOGTofYx27PTf84a2xu1308g+8jYjESLiU2CUgCC0LClTEongCcL40PPDoqLexNr//QFLLfPI
cr1qPPBJBGuiXXwLY88zUJ2aIvZ156KlGHv0oNJtdR1y3+rR6V3eM0FPntjWQ04J8UN/N+/4y8w3
Z4gIFBb4va4qWXOqs+fSK3PQ52KctT9SALJynsqhMpNA184qoPDx5JKruawFEL558XdXOZrB4Ua1
6+RgM2pcUkG+arpflhCTmEBRFa/0yxwARciPE2SD8wcPs8sKxWuGsT4/KXNSX1sCENuHfYbsH8al
LZlmngWzmixNUp8DSrgaqqysbE0BIO2bqkonDkSy5kwOBjUxnqRy4CnMKTDEMQR+yWTrrKfZzxRr
d0l0VaSYR95Y5FB1Ra8rwmdgbPAwIVz+BnoHhYeYnslgysMEzYzTBtwdYwXmoifRtNcneoZOC9DC
5+SzX0fxHJHow2ZOWQnCOuAuvoh78RdcApG9mb0obFJ4A/3q9kYq94/ZmU8GoegOrjNu5BZiNk7i
aDHnbXhqdldufUj3V60a6Jym9lWAiAPTXrN24gRHXHK7lCNYgMWQZ5IqE/I2Lgnm1Wph3r115V93
gidldbL3R6BbQ3eURgnRtZEIjU0Zovy6dln0Qk6iJBSpgp8UPSYJ8z+7fzBH72j2wUiIM/c06rSk
YX0yNS7ngi7W7ZnoGxe03QdwwU/i13rm96rAaXeAie55+yGpeqE0lfiR+e1phdQ1yITcGrsYS0Zi
oMyaDezwhBY6wPpFGqIcXAjggQoCBvnTKzgUHPACo3sTGrJSe0FdYZuO0FPhCIIOL6r2NC22htKK
5lh/6bViRMS2STxBlCPOPRnaWzjsgUJxSg8j1DoxRiqe/1VtU9TiKP8ZNPKDm9GMyHCiPL1j/uj4
WrH6jF9yXgOLFnZp1wbiY1RuqHDxIE5hYiAtCgou7G8b2ePvLEN/GWzNYVv8Tg1qkrhzcDqAflBx
sYPi8NbV8q7Ek3YX46dRoen+UOiG6jTCllj6LHyW0kXXvuX2MvrH+WBo/IHHOTCHDr+Gxbq+spZx
hAO/3txc18QeDNxV+mUeM/bcKXuQAUjJn+utzLJakgeGdDGrY1maKddyxCeHMmNh5VNnCiZaUJ8v
yBRMYcrkl49kHrua4BfJqbEroiDdpxksUwVCGBV0TEdy8RaAxDUShkQ63rD1m13k+uiIjd0bgtTw
AUXMlbtJI7SfBDOtEy1zuI9BmY4u1053j5FD43/XIb3MY5yGTigxotZ3fSbsMya3yJB0EIeGAUjI
3ouMZtQVsHzL7N0EbqGhNwIXVnxYXWtjfKU/t8fE0EZshoixeR3Emg22wJ4GsUqgASolT8oiV3JA
ufA6ilDVTfO/r5NzNzlJOs27nz1DJJQWkUJkjGWFpYoKopQ4zqYEM/W1XPpUkZXae2SL8XP2lO9q
IvUAeTkfiTX2YWZFWOCnDSOu/90S/99yPmoyQMMG6XulAoDgb1jSX8kjuFD4+6D2WKKVKkRCOcHc
xeV+LN6PKZD1P9FHhzAy6HMsM3DF86gdU6aX+941cCbxD8b2Xod6xn+Dx6Vin2wSlKfhn6PBo2O/
FcPr2HJilaxAYblmybF+p0WYjKcWtAAvAYqkIdPDIF1iLIMc2WEbRUq0QBjqCcx/hkvrbQY2Znlu
ByZ6iZfDIC3XqFy8OFnRg61q5mfn7QsNU0rPP9IG67+/+hjNG9G0SW2zkN8XKqtSMH1DP22FtVbs
2U3JbasRWD1I4ZUpNck3tEOQJwTpeM4eXGtJ8fPK3mBhU5CX8r0MympoTJK/ccBrWQnYene0SGjP
OrFxhXxJk6LHbUyg31aOA8Yn6p2rCooqKWeQSYYZgrnneGShUPZRT7ykhi6VI5bghNrL79b8qAjL
ga9jJm8+mpG46IXfsc3nWwQEQOlkKTshahfNUnW+1Wnkb8McFcwm9tkDi8IxMMHHaDfjOXu9FX0W
aWf9caowB33u9Z66M2BKXkr50rPCnKT6rsy+FojlTO/hj4dGzU/WC/GpCYFVRcyDyod+airwhTTi
DA7yEG1ob8i/8IdKtRy6yZbiesezmk1pwsBIVuBw1+lZPbXMaKlcZ2jnjEFj0CEpiuyhGLvl9K+Q
wfNggDrWWDsZmfOlZckHHk/zU4xOJbXkI9OiajsjYjzsO1aNLKanLRSOtIgKshhh1og75BeGbpDA
1TPFJgSEyx9WLmY6Va/QakHGgtRnamQwQ/wF/ALghxpBIq/FN8YkD9IQ3sNKPIlc07YFHMil077j
DijROAiezBRwa3d+Uy3Dn7Q2MG3AoxFTa1bayBnmshRB1gFGZMZquM8NkSNfmH4OowynCnm4AxUx
D5jQsB9xZDfE4M2YzOaHYKocJriJj8r5u31hEX9q7+XKsJmi6gGurkfpwczl6mbtCYa+0ljvnIoB
bgdWLtUR96s/RUajxKy5XpKfRsAiQEh/79JdFkmqf17ZX+IBjFPchvTO3/REoakQ48txFlPDBaEW
fDpMoQDSu/trZUVnmPPvBdG+/Bv/8F2MUyam4lmmRyPeyzZezLsyx9wldsGMViJpcX0HKwRCw6ga
Wbq8cHNvO7+IDLjeW9UZEN+SyGibl6+9BB9QkUsoIo9ZYleqLSJAzOI8J/3HLXCYUWeR3BuP81AD
CZYJ4rH7TkWMdcFXQmtyMwtEMr7eFqetuI5iiRDc1Qo3ZraKffKP0k1z5zpdwEk7JpeRWPAJT5Mz
EahB3g4zReA+JXStqT7SjLl7NTW0a2ZlpvSYIJNzIEAtcjdBTQZHld1odYKQrzSv+rXQvIjlDJFg
gXE4pipTtvZOVZqk/kjGfegbGrbBGDAIi4gmovtZYtK/3laLQOhr0LeODnT8H+MQBGMwy7g8cIfm
lWvEOMceNLA68JudraDNjoKUncpmW6kjk3Lyu4R+CkoJnq3ttNC1lEsxLg2HI1T1Hc+gxkXUwZMJ
D803l1wZp7OaSK1ZUDPGu7FvlAGTT7x01Ow+D3xZTYwx8WjFOQdoI7DqQg237/gOSp2g1Zc6VgrH
IQPXEPt8jukzQMzRM5O2Nu0EQHXsFlP48OFdWTohoLF/CEp7Z91/0etj1XorqnJm2IKaoDZLGguR
vHcBPhEu/GPxY1bwCARdRBUV+PfXoFrL72QfcQj+CiIxmQCDgrl2txEcguXOjP3PsE9IiuFEuzGP
YZNmY7yuNaELmrKODFJWFEgAm1dnp6m1PludFz4rYH3wHbYUO+dukNI5D36lg4JVwj3ww75MeMlK
tkVeEGL5cJvzXZYt14a1TOrg8Qh1SKZ6iaHcp1wW5Rc134KPzSbKCYSlWNnS9uPyHwioD08bhj4U
NucxzsqCnzPN+u5kyLHLwQGSl5eFYHUskEqnpFtu5wIpw1ddxBuUNTHLs9sakbW6HWdUcmtnswtE
cSYUQoCn3UsA6cu0PDCtONmZOXE9NEViIUJwqwYsOjJG1t58anRTiqG10ZEavN5LKOAmJLczqwSo
gKp0IRZnIo4O3NckNVx9xgsMPq0Wk21z5HNASvlf5fCcQj1Dl3/yX2cbWrCPSjdG5KwDt/8ZPfqP
nPpmFmG4EbfVcrWqCR/O+dHLMTxJB1SJ99j/lEfZoVJRDW5xJnikd9sUbXeZToua4K2tIRgJ2tNv
C5QFjZ3CjUGgLcxqEsyEWYb3dprSVNWvMuYmCJ8AEon0fOpxoj5844xo4wx50z7at2wH2APIGaJq
ni+OL23N3iuBtmSt9C+NtJ2Fw99SVeLXCUV3/1RQWoqP14K7rvP5ulJRJmY9DABD+nba+9GPu85x
C2AwsH8ZCukvJyjiccEHVx8+hCZJG+MFwKqSwAr0tsLT3CBVZ112EGsjCFtSGIIC+6fKC75tae8o
9KTEv+hNWL+tXn0HRA95RMQzQY1yZKifwdOLtmYJiZrrQIAp+pTUHTwg6jYO6ds+Obd3xqsjnr+E
dwrv0UJveVX6N9gGwzkNA7y9/Dv51k1NBymtHki2kIoTuZeK9mFCRaYpBEeCrtJJtkxL5jYZTnnJ
jgEf4REExZYLUonqWJC6FdR4RrmeoQSjKwRVmzgzamTLP3vgWn6Hz1YHvbIiwoZLox3O0KGiYDiK
5ppOJBy2FWk5XnL/Z5pUx/tZSS+nnQRUu1k0xi/y4oY2Y2ZNTULCBzmGnuVAolYm1l1LbhbXCXR8
Hb5syNAy3qHKPpAaC+xjO/DrJl9unYhUfkpdUbynlct+gtG1Fi7c+9Vgkz7QOCBKooPppBm4v9ZO
vAKmvEPb91FA0lYDfYz1+GjIy9e7vVTJFRVRNSHRBwB1LfboEnO2yohIM/Yk9Qs4gqunzhcJSPCk
XObKFF+VNoqZp9zhvvCtgE1g9rlobd60FZlqfqBnj7cGm5SGapUSy2j+KVpUqQ2Z6VDfVmagWm8z
msvsDMDHdcbQh4rrFEmdtPiNin/XFXmBNG6235uJU0H7Sv4Ou/8CzhhC/v8tfQ3JU2O8/0WrJzaQ
Sc2/IbhLe2rCzPES7QOI1UJiwnP8o7FEYURzlY1naiLIXXvi1duzMKAdk7dEdyRgjlFKVNmWR4Im
iq7PVdl4vesWhwPL6K944/VPhWGNxzG9lxUDWANwU77YODjdWT5d1QXBoWNG7/udfkAtvIKmrKWH
K62Ao9/MaffPwGwWuhCNZoQcQhw/beGZcQVy0Wm8eiLSOmgXy/ekhfMrSYplsqvJ+ENp458e7ho9
8XMhegMTEq9Ahga3k4HW/8ZpuzK8Tiy2ss0SWUi3qZgQ8lFsJor9z8FEPNXZ77yt167LbCz1i6Ua
jaT55IUxrHPRe8HaBCuXb7rD8IOWEulML43wsKuASRvHLTk8Yyuv/XmloumP2FVmKWrxu3SQEcC2
ZqQG7U2NoME2PydgWvUjsToq+xJRzVzxFgBkPOmOGJ7eZDFDOlUOifT0dgi18MP06WoPtQN/kY2B
ML+/rifmuKCS6zPYAjOjhvT+4BvHNo3iDFlIYOIUaVndTx5qv28rH+Hbeg0BC6zxaHMWzKM41dbf
dL2Jp1YLP0kuZO9E1NgGGBUAiiEpl0FRrwTSZ09cW6I0ov1cXrjaDEGE5FDBo1hNEXbWs15X2NVh
HtsFmqYkb8XL/kJIaOvJVn3LzjMJizP57c3KdQYVYpOWFY4a0SZ2wwSbbU5G2Dl9XmL9CN62rv/y
6ubEoN4woDnnCEWhg5Fhds/Tzka77yYP6vz1qOsG+jjf/Pq6Fp4UbHzhHvqDRpejCQshomzwRAyb
S4iQQ08LK9pr+mSaBy5LSGYfFer/QDwO1AjoiVOTdBeQndzo8tCNY3PkWShZNNTBSj/l5ogtsNB4
LRUMVa6AAtdNApO/K2W7EaK8Ot7xUVlaSa7mf7BK87BH2Njjmm+YbawxIKuygIcqxEqNz47ssP6P
vit+Ha1sjyiSeH6dMd0zPbmWvvLIOGjEyAQrjljIRHzfBN1T8nxfsZpfusJuk1jEK2GONsU8vmUE
w1yzsslHi2lV71DlvAZJETI8X3xbhI0IrmqFVX9NGpSJSwph98WQyKP7Rba1IObQUA3HFjIzKk2d
7KzsdNQxJc89miMcAwwVBG5w/QrGgeQlL/IwA9rMVe6u/nxY+v93CpVKfnKCO9y4GAtIU5cBI5pr
80Qh6QpPyi1cbSupHYBVOPUgU+ooowxzwW53dpsQ91Fp1cMByg7sZK3xND91fTLzUO4o7YBd/8RI
P4jqg3UZ1Y6Ld5W8NTAwtkt1kNogs2nAivDhFXjOf8L8i5ufA6+LcxVdKrnD1MB6DhQGrHKZqtmQ
r2WYPX2d0HK5UIhsnv/Q+Up5ZFMMF0DZtGARyUlRk4UdjAvClaMjhkNmsVAA/gvolFcAC6CHxkzo
k1ay19IJErurVL9jQTesReMXSWyvxK/uXf65qjeFmj5KOazaMozYQLRFsMFzmdTU0yaDN2OLytee
VRat3Y7IbaDzUSOkc7tFn/Ny27KiyqEbkFSWW8nASe/ToSwbz5nbSlGzr/IE35yDpyZ4ZA+i76s6
q80tIwp47MfxXxUOQY5CgrQJfhm8TfMGGMZD200Gqe58vX9dOucJ91oPtgLYrRWw09W6ACoB8Ft8
LSx6FG6ITiR4JIyvoOGymLjgIsn2Rb02LwMMs/LNMTtdjBCrY6PnEAAJ0U6RNBX2RdtfMwVTl3+4
w1FhlUQDa3v68oH8CbiFUdQPvJAaG7t/D30gBvUxBl5KVFh+b4Q6tQ56IBuyLz2Xac2SBYm/8Cgf
cp8gZUkkkX3nbEcfL/5gUeavSrL3f0dNC5e/+pO+EZ5DIuU2FjD3J8qxbw5EMhZXzKcVngl3apvM
dY3b5R02CcjSO1DjP7pXrWiuRChRa+cfSx08U2JntRbCiysF2EGVI3j3RDAXny3VLOQPdU0lFRiB
cLTU8P1+VRMIHQ42wzdiBPGS9tkv13H9M8fK1IqJp9SXpS07FNQrfa7rpPvBe5ORrYIDM85Ikomj
Qi1h8PU3XQCIohdnRVv4Xq9TR/fjM33l8qwFMjn7kDLnjHGC30uT1JBEti8vQ5kUxtTHGi6/prF8
iLpPbtKF5wc2fXueEYwMSEO02fr4big09KTsVNu4E5eYXy38z5q0Qxr89JL5wmGOaLLRZodg/BVc
YpZBg9OwKPOXofetE+XVm+ukltzxd+OoLkzzZeNce5R1qIiDm7xCjniyJgfh54/hXDW3s2AWNKR2
zsrR9BpVqV+y0AmMfuAhv4h1AX4xMIDVIRY2NmjPgR/kiHFeMFOR81y+TP3u/d2UzXqSL4xL9OCN
7PnkVVQzH8NbX+yxQ/N+l6y++oz6b/9T0ab/P2mQhnUnWcESLFF7u8okpVe9QssHROgLdfYNDgBQ
VW1f+AfbHEGoR1QgWOhdpY4Azw3/cf/nDm0UKrdDs0ckwiGPgYO1HiAOdv2D3a0AeTMwCS1fpiMb
Wo0aC55tSR4W3BJUAemMl1BnjQN+lFJMOEt/7k3yqrSOnoxEZuKtbffblnhdJdgAv3RD35Dtks8d
l4Xy917/Bu7kQazQcHodG7Qe0bd9ieqixN285e6DPuOpzRvr0OQWEyiqRgSN7wYNaYqr+KTu6ZmB
f2Jnz7LFUkd+lTgYb1pq/EAXICT3c5jNdhNLwONkP60vJiEbWa/d+H7rEvRc/L7mcKp0ZarPZ4n8
11XZZPMD9HnufJjfK0u6r2WrsptVTiiZ0QNh7q9kDV2beD/4J0G7RcUw1apzO0Q5Fdbz4CyB/WVC
GB1+7X7Y74ACDsCQpiWN8PS3S59Ti2Rqy/HpAwdQUlQLXhjT7CEmnqdxeqnS1yOzRDTRu65O718d
y/GU2ZQHkmb9Qt9I0W94Iv9FQhK1zoARGN70wJroWDISGWaJXSavV6u5AprSr0cuBuTxkpEdL8dc
kGF3ggSTosc1IcCyVKx/XIbrGiv2EcqIzYfvl8y4tHQ7HTgLKO10BYZ8STW+Vszl4KAFMvZ2WPNd
//zSW/ZbjrXu6BkhsDDESQQToWXiuH26r+NAO5j10t2G7I0xUXucMMnISUApIQ7+qsWOZfn7ahzu
cMyuVsJek9uUeahHqjYiQMwgUqZCi4nY8b98UE5IxHIP371vMqnL3w+emFnckl97QeKYDUGITzeT
EoFEKCgRe9467zmQf0mV2CMO8K98+rafwEbph6G/YJ8EiBEh8pWkfR1sTDGMGeB7jURZHtQGg9YC
5F3rSz2wEES48evGpoCAFUZ1D18qGdteXTGlkU3pjz0TN/b/KLDV4WACBvMQYsmzupwlNz7ZFNb4
SNV/MGLF6IE+BzMmkTv2/iWs6OkFJdp94uCULsHI9ZNzl+OOhtnpF9WhnBP9dIHxNikgNgma5sS+
AsYSR1BvBAm/vZDDO2lDDrwIyHzkKHPj3J0MtzZrE1u+O18vdrWF+T9YLZ1K9DE/UfjFLiPJNgco
bjtRUGMhOirzhzA3vf4KLOpK6pslRa13nBYLw+k9C5sKQ9RPjAw9tQ0OzJgsl9yCgn/6s9G0mjgK
gWnXur6IHYLMx3nDH0mlJ8PQdB71Ej87O2dDl7wGcyV39bqiaw8Cf6NRcQNOmlIqcvkCzM5eN4J4
QVrb922fHWX/5HdVs2ud40qtIpu5AEhSxvCl/ehnd0GxK/KSjgMCJE3chbjFJs6tzkQaw3W6YB4u
4baujiwUaW6pWQsTbAydKWNTI0VCVBeQ0e3QHeF6gvnii8uXjh2ApkmWC3nXp3oR4XVJhcYkC9JU
xTrQ6CjEo7XrX+ZWlzvnbQX57B18EgJqbA2eZka1zDA6lV33AQhzu+0q2rdHNrHsM2tUXt9Dkwot
SV8wHchh5RAdLALps7pH2viwGuIVHxE4Bsd7OOqeD8xvUM29sSajSO42p1O0Qaa/Po6qf/9N9Hal
hIPspwao/hj2hJwfuNCav6wqXVR/mXMuIIgwWu/S99ss/B9v7Kg22eBTxe8GDI7EqnjlUuywbc0s
JCbdNfmfm8nuXK9LKeXlK0mAACfk4MJF2zFboOAjjK8E/KCPFG6NlEJ/Mw7HCV8jRTgZZhL9419b
S2gYLmUISUI3rWt1Tv1+qbksL47QOHd5PlKQMRqod4iCTOpaKmebe8tJXqYTeiSg5qcE4rKERNV3
Snwd/bZvYsbr9VjRGpRw+yRdl7xHHBxUHpbeZjupAbRdLmDJrzV/z6fhxlH4ufLIyQOPd9YaYpur
gUy/ql7id5XNaKp5kPTxSLXxvc5Mwo3Y94uBNrfFw2dYt9VEnu0cn1waP4Ux93tivwPaHyQlCv1f
JhxKrDMlHmuNQ+OhS+QISfUIn+UEu0LCgtr2EDpZG2LNt4ljWmHG3U+nP5bG4CgRME7shFMV66uf
rxPtKlVzUq+sRb6QFQ6oSA3oQn1Osca4itiYVwyp4ZNxR/FqoK9OJPo4HSrDMXYoAeQHKlLXTrhR
SK1lEj6IUMpnphpQqrSmmPNb+IY+6So+aSjBbAaVPZoK0Bj2pUiRcPYDmuqGsN0wzF28w84HAdWU
O9U9NQtX2FIXYW9ob+OAJSa9KF35wD6+Pe1jzgN+qnolkO2z/5Z+Y8zNQRmqCkRWGfc7foa+7K+c
l7qS5UGPrR2nVKrYBdHBRvWcwstxMXu5N/ESlKugsjTIN/Klo3vJMZw4VTWUGy5A2ZuC2JBvJQsI
v88/hdHZHbKtBx0is2IPsz/DXjMM6JXYWBmAUyCdZidf12xA4Us7ntSUQHOCTTPU3hjs/4k1vbH4
RpjG8+bV3xnF+9WzzpKlrSwYHA5Xt+jqC31zzcTYZdBryPnoomPgBr8YWu/nWqaM4fQenbLVSMqC
Pvs3vyXFlTP7Xvtc7F3Wv2lYoichDN4eUdtUG/9JIZ0+I5tVBW2EV9wmwT0YadGa39cCkLkbW6rL
/pQrr33wyUISJiULLSaEmOmcMQKxk27vklKkhYOWmXYUXomNurUPQM8Hky03PWb/LUmuZ4+IbrOO
PJ9l5JyUDMIMniePGr2cgflm6YqNcTSNJHAKzuONdfQs/ik9EkpaYhrF+5AM+tT/1xh7fh34dY/D
lYH0gWX+2gKHY7T5ZXPPsb6fWNhgvyooGCA4ShguHBOFe41dDYlBzVH3gR7LCfGXsoSYjRaAqUk6
QsceWPOVN8EeixAQl0z7EeWfHabH6m56C5mFnfB857cZIVEWhcrvm1wj0081sMaiVnY3iSUS7iin
r05E9FvQqUptRQMmOOJXE5gq8qIa8YNZRc9vLqfFLdp+ED41CHeXUwerLBrrFb8rcti0sLY2Xm1Q
F6U2tTcLgXT8HWN0tzDwu3Qmq4WMyk17dGJdtzqZvCanWyYZaN7JIwIFbU7Mxj3QbehVH0v6Wwcw
Ft3kasetFEHrMOy6asI9rhCJ2NGOUmOqTKLLAIvSNkx4RUBBgTq3F/jwmcHbSvw+IZcQg7m3D0CM
Msa/fWmQJwepfXBQNw5qLxT8it4SgtGHU+UcTGkxgIfWI8G0LW3+4PAi6xYVLejeRjtus8OZgE5T
vWpcZnFijPI6b3Rcvb0IAJ9sb9AD1aCWGXKMQg6Pqj3M7cNTRqdM2AGUWIdI5p4MhMjRMq3JqFa7
5BRHHwcW8p5UPuUhrm++RutWViUKiPGeRokdk2RuXyI4akD20XoFBkqjRK2SY9aPISnXjQnnNK6s
l363U81nbEhVy4B7LmcaSg71AC+v+opiNHy03cOJJblhRRWeKpdK3DaliFT3LUogTimGynEg1SMo
s6Eglw1tTp/IRCZjwnAdc+PnjmtqKdAeY+STl6+fq3HaXzoOwC5vNVXUd9tHOhcfRQ4hre4+qRlu
23dS8F2h9B12zAONSfj2DtMF7aYaMLy/5pdV2Mi8qtaWNj2v7ENmMGMXFbBV717U8DhFd3RRfvEX
OEaZ1O/NFfdngqiGZRuMv2l3ZsmMdSes5JLC5VaTIiNyGmNYl9zqAzc/H5SOJtjgXhMD0CDPH2PY
KVC/cJZ5h0+w5tgLBM3y+sXwgR81AWJGeshkK4HYghsdRCvGdwDYw2WSe5R0fRz+Ytl06p5aL/HV
Ek5OLbj911LkGRpxMna1zQ2DeDY/pd1qoLxwgV8s6znAlxr9eTd7G39kJfvqo+Ov/9U6Vh2a6W/J
KqcMMLXb4IptuZwOCb4DrvGI63cVzXK0kc6zNVrmrl8fStSsI9CK5vA/9reF8/RhqzgvdrxKv+Xg
Kuo2AOl+q4x0DypdxGKiY2lK4mMHoyJny+AMhQMNlot9geZ/0fT4VJfJzEebXEt6Ku6ekZ0nRTsu
O6QodAo7YEURqLFXm2Ajq16pvBZIT5uTXtLp7IqHZzuvzyImwCFp7xJS0xuATqngpOsV2YZ0BxIl
Tr27T96qZL0NNrT2p+/P6MLHlvRHhBa+UXcOpTn/RBhJ9Z1ZbsKyzT16UE7wHXakiv3FVuSm+3PU
6yx7ekWOXEvetCM1+yR/Gl5gQg4D0cha9dA5hSlGbqxHbO0Zk2zm+SSj3g1PZ9lHUd8OW35MioSn
88Npvw41jfZLBmHzmn/r2dVbZGbXGjaBWbZXm1GaeZoOoZONgOoS3fKpQsvpFdubUP7VXbkhOLso
M8q2MmoyPkt89V0LD5tcGRXSv3s/7+27UIVAFcLX/CaSfx76kS7W4mEtbWald65vYObwFq8O9Sq5
6qdOb5Q9FgCLJ0+ITSlaKtq2JV1CZRzs5edfDvwcJBJeihEAH/flSCCFKkRvYbhJdT83EW285k6L
CKYVZqrYLSb/UxPkhHerDFISY0ZPgntFBAafE41VWKimm0BnY+njqPjYFbZ1STy27E5hGS41BHqR
FaazMrfudu0Bi0uC6jSPCyUOpgr8LNYALWUIRusCqcukjLj7pzzM858SF59Seck3Z52ZGQXon3Tf
lkRKg9z/oq5osu/Uwx6Qi3GYsNd4mR945rBr70PwCRzktfvo2Iu9LQL2ZweJaEkrFBAaUHtsprWq
zaaKoiiiB1zJcsGYTV7PZpau/DnIZyb3HmgF8g4/d4WsqLdJBLgQs82/7vVubIhB1cas6EFtLYOs
Z3Rwg8wlv/kDJvdVJIbYKHnLFKzUfFE3mVGdKm7v7eCdeDMs6zHKJrKLBSPhmugX3hG+rbEjv+uI
7oxCmCg3tJZJ/nRKxgTIKJdXJqPOLUfGUIRJkb1TKwRpbG6mOeaJA6sppsYDsRvbNe3n1YW7/NKa
i94qyvwyyW3ZNs7KwcpkUW1BNtp3djrPqCJ9asjnJvxDJgAkzPJU5+Y61NqAr0bztngItItgJWJM
wGKL2ez8Da+58EWK6B+tKMtByjTcphU9saN4YXPe4KpwcxNrN0wsWi9O1YhedRxggm+X7SppLFRu
kpKo9wggKjdltbiAnVXLToca0kqXNZpwTXyvYBcLIp8/vp0U0wjt9i4f2gRzlMaEE7QSbuaafl4k
hFJL5vvsF+ruXghC63btvKJTHcuAgKorLngdXBB+0/rXp+ydaufCRHCiehj7IynjOVp3/cPNObVq
bitzp6mSU+Htg04bkawgOVJ+RMVRr0OtkoleVreOvzGg7tciIguFaW/v7zrFLDaRVasV271RSG/9
jEySAUteDpiYkFEiF3RKGNskZh2jRMCSq/xtOV2HI7bxpYPXY+v6yKC5HWve8D+OB9j6pljD/6R8
DC6gi5D1aUxUjNS21hWnzJuKKcyzr5fbyDnsJj+K4QFpOk9ZcPzIQCK69Ebal+uzDbgz9w/rlYvC
JHl8/lHqythK3oO0iZVI2LL+NWTBcxj1Euc6Z4+Sc0X93Z9Ag309YqxDSOG+b1VIcMjfmerWrYb/
jxY4288r6d3b/zmh+Pyeu08eMQc2PTkoQpZ2l4yHwM/xf1FD+lR5OYdYFd0o6hZC5PZATgloA0ag
klqLSWKyrFQgJwcr/YkdvCUcvt3hqTi0V7dasRVhTYVwcrgzn10mFtnFrjXN3agMFQ2M/4if4HWl
SX+dWwqK4/i5U9+dA4XxtPh1A+nBSopZGHDEiph0pCjD0VRdkLYTRcIRXQPxZmuENvhFsDME4BVV
2nBWSyTCI/Ar7xEgzKP3SF3MtHFxBN00fpaZCARbLhOkP2blFdq4EAsLi6b5vn7SfY8zZTpWijJ5
+PojmcKKLffVGltSFDhHnK37+6Qk7ji+8HM81EC7c2xbT85IUX0Z1+7G1qj7xlgaODiWgn2LWIDK
RKNak+QlSnzBVv1+WvSURKT+dVqnCHYSfZhacuzgU6UnW0RpyXzOsObQOlrxbBRPuHfE9qgV2fn4
Qyy3FLx7Zi5xzKJyERms6UduGIvnvQ46MOcz5GfEzucMiD+XxQm0xu6vK7G6mLahMAohwQHlnz0U
pkC3qiRjskyz9QqywY/QXyB0OwoVV98azhIRIHH9RNQrUfcmI6B5QrJfps7mkLIkLo5vLlvVR6fS
HGpEIzMdstXaE27grEHjq5sP8pKWl3To1ULpkbonNNk6ESknhyh9Kn0p5gceVV/pc7cC5ZTo6+je
+95vWzqvkJfc8LYtVWDJd2bRHvZAF9vcH8K82H/8yNz0Utp7XjaeHnsiYjEF0NVqX4gbtD6JPUyy
hZVdmKZlw0tfHBMaxidJ/ItaA2r9tkr5hVwT8aBgSTIq15mOh9HM8I86AmtASK6sbcVeOhZOhlhI
7FjiUQBFygg+4XZpEGwyduB2HHgtO6P5MKrvQ+xDCWxhfnEFwIrChC66kTUiNyA7wL66KZXk9GFQ
VbmF54Riqqb4dL3vubUCRn96uu0+KYiR+6y0Eieclll650jZp2B4zUvdIXKWVBdGRJ8KO9tMRQff
gh+lBae/khr6sIXd/smdTt/ZOjy3jgwSVnJbH4gNTBQd6CjYLN+kWWcQid8ljWrbCD4m9yPF6hUh
HasPuw1oSTpV9igcm2q4cxOoEdWY5wKGAkPV7YrQBeopeQF/uS3RIORk/CUxKpvkUwGDmSADsN7l
sLxMGtON7RY20rurdKQuUodSLqcccpFsSk9Kk2HEUsxBcSah4pNDLC79Rxqt2wo55CZzSkfkgmgW
e4+C+Tw96W6pUWurWj0n8P/wGlAV9NOYWOz5jAg9Yqz1b8Nd845EmdaqjEoqaeae3ml15qH37Ukq
ZEBO7PMhJZdlDNCEWdC5+jHBhnvntiU7nUPpTd44h/TpGr6yXAaE1IrayCUSCOaErNN9YV9N4lzw
3/M/hiHeZAEZPFkz+4OjTE6pNo2TMdT9kSYvIW9lrAPDMhDicC3Ro+Y+2akHaeB45HM6DCT1Scaw
fq4HMiayzXfovd+3nH9DgF7X1LJzJ+F0advnvSoya+LFgC8d9NprYTkOGEogsIDLko54wOSeP7er
iXDyenGebzX9DgEx4K+NCIu6hAJ4P+rt8I0mGHEukejuAaoDEPJhTPFgt3+fUNq+NwS2v9pQYMxD
3PeaetDKDMr4KX5naLELhVuns6VoX1F9wt7ieFwD1rvl6ZPF33Uc+NX9UXs5RMNyFhF8IlbmJ0a5
E97WvLhthecrecE6xjnpkLNGt7bXiuuJv7ciyUz4c3igL6u93UJtU7MI0jJONCWLJ8qzx5iyn0kX
wenggeHETh9LRXzKNaAjr9RTybt3Czv0z9KHIFbm0usYr2Du+mq572ujiP5M9cYV3cTsDpoHRMQ9
bR51Q+X24RNjtbfIV2RTgIP8J/oAaoHnq3QH0x4FNB+FK69Owr5KQEze4m+sAA+fa+FXTSI7NPYw
UuYHCg/7peSmVzc4hvQrWMP27lg0n2Q11iUm62ZSFZq1LgWbYAuJFsZt0m79Pbdx8lI9eWFhlTO7
DU/RrFxM47Yhnhi9rGBQHqB6JG6T4JK4rFnReIqd+Mnbkn+1ioeNYHMd92rBLtEx5SVMyC1WH5us
DnG0E52uGpwynC6mcAsKpoNgSK3p7EHgAz/m5MflFzPdyWIyq/XweuiyssgvfVfkuWWWvOqSTwAb
adu2XWhfHebvCb+sLZ8K+zL7+rYHs8FGvKDCKzZu/mZrIbjEDnC3Alwf1FVe2QK53PilObgZ55HJ
GhRuk4oJMuWIrnwJ64BwCsZnHSf1On/MF9qXemiaPTkFp94JhTyYVayWkQGJdbbPvbKbK6RbrDwZ
49YwMciZbe/sCaxBzv8oISLw1US2jxRS0ksoNMEhYHPSSX6z9XefO2HX3tnOYv/tG5grCFweOTYr
ClFSNV7cpyd6s9VX7C/zdehi4RdtoP1kfeZaiphNOUx9/fnztu4wOndDGATDPBOl6V4jeSiua4Tx
h6XPgZ3K4aVZtLzsPa0wzfxMCm4LpOy8r7G2Pz971i6YUrvzyvY5HE7rvdXqVxQnQIdwBBOVhY41
LC3LgkpMMYcxyNrHi8TN83fW5Q19bHy2CaWHB4ZGSiJ0zarSj7pAS6B3g7GGnwkl8YjSdrFK3JsR
sltUhdzRIZ+LrnlpOyYp2H6gsocRQWpg68s/t9UVv+qN2YmEmwTfr6aXWCrhFBSbr4S+QqCWDjyR
H+2mnNsYJmmIhvJxuSXEJdtUk2bOgxXROtBrTUSg9pYH3FapeW8TC1KpYq67jlmcOJfZDQ5NNt5U
O02+Si84G9zvgXtkCzhLduQxKGRY1vy1A6uo5MQ2KC1Bio0oXsd8cfH3x2pp/OfjXdlpPodPQ995
GSzqNj2Mex24umyoj71QzUevjGOhQ0QjNhvDrrmhMKzc2nmbkekuxsWVZsEA7w+lFLGawtm/4JZH
avSENZwCgUrgltvfH9oF/feFE6QUU37hNdIVp+n9DeGuSrlgnDcnI25aUIrvy5lYCpPhzWoYzjz+
Chbu0/Icm2Gu83rv1pQkQHp+rARiNXcW5OY9D0OE0mfNY6ctWRtzzMSbNeCLzBHCy0wtBWWYbUqQ
4a+rzgigzaZBp7ZRiDzbjJwkfPk/8F7b40hP1vFrwsWceYHMe0tTSJwPtD5L/mJRB08N0MAUZwjf
13mNNavpUup6UwOYvRFWOVAKL5hDbu0eswKxjn6bQqTga1RquYpFhMIR3SXb+mhebK8pV2nXex8d
Wz9r2WxluPfZT/9DqQ0/ruF2Xa0cikLvORc7/bkXSZzAK598uF2kmmtmjotPHSUnMykMG16Q/uvQ
TK8j7uZBG0z/C8hkfhlsHsCoasP0nFAnjDgU0QWwWnw+5cbYsJTVK6kbIafEknMnaa4bwWQY07u4
9qdeLTXmML1aoDjSEaQWWirnmtUgurusIdPjSUST7J1gAAIkyUuKqmrOOGgMuhO1oM3APH6ri2Ef
6HlpE11Py4E8BVUrRNF+8rBAHE0cq9Ai5emrB4maLxKrAMI0STqny3nqSpwtqX2PwQjBtljrhNCQ
JIZoRgWyVj56OZrHDpcRDAes5EhxeAXLdmL9cr0I4WHJcffeRKGkssvGHVFnglDcuFLj06ZEf+6s
J3jU8OkD2oHLHU+E6CYW2l0taHh3dmYNxC3ld/Xp/HrHRLvMP2bDkfcM28fmaiEop38aACbJtvJp
l4WAOFEW5dkrGHaHfv1X7dJVPrinyAYLrnTk9wrVhwYJ8sNY8u/+YS6+c67NDycc5LpF5v5LIdOI
nNy7DTXurhy5HwuzoAm7RhFMjt7IIcNgHKA9iBWyI5ZV7eJlUvs9ylyDG9bqdxallZjvu+CuPKuG
8P8t6TTiAbOpfwHdCJ8JZ3biUA1Hqs09vXcOF7Q6diRV+jd6iBiXe1/svSNbK9IFdnJ370Q0zGG/
7ZVKWW/o1GTa5UOCzxu1DUQ5xhAtU7yu5VowaGQ2+c35fbv5igg4BCOhbf0w9vb1mnBBVLuaqYP7
2NjUHfpT50VVl0vUPDaZAEF3BSGVUlYmlV+E45iV2/6iDwF4h4V+A3jOVKXp6kKiKHZfRYQ8dpcX
QezckGnEuRNFBo9G1rD76bWr9JFmhd4S7CYs/XBl6F4eB0kAZ8V0YRxghSVA/KASo+d7E+CIap9J
UgfdInR3qTDfab0nn/abxcrRN3X64MRs0HMHTvqCbqZTC10UNofttXJgCMX4b2mdTg54ov5Yi2A4
XrO921+DJTPvr/yNgRr1dpwpOEX5ju1i+swjKEP4XqdFsGuKxxtXg0Xd4o9IkIBxDuYm68gZaIPC
bi10R2b7MBPU31zvKvn/rPaihw1GL4ojzwHS4Im5lWCGWDpuqtpUhIW4tdNNYyH0b9ZxvTXapKYz
cQ6ZFYNCFOBUVQcV04mOHSdzhV6Eyjy0xKiVL5P78BKbLuxbe7TnfCP0pAhakfzdM0EjNKDTReoB
nTYNYzooqBnTYN8aIiQWKqCgc9aNhKxUIM+kIxkU7Mv6pM7JcrogrR/WPpnxW2QMDnsWUFK4Y3Qd
ITMYCPWcCJNo3X2VT8awbBmEpySPHcBQXyPziyFTO11H5EsgVxFkCuCQk00lWz3nsi1h85df9rU4
wgkGpLXwtjrD71ylFtwg0EqQ/8Qr8fPtum1iLgRYFWbXoeAny4+t7v65YvsM8N33zvJT6lLpP9TK
b8rc0M+I/Ld5uJbOOYoFlRFNiSleIgMd5PmhmPpBDZb65eVrjUML4sAte6Oz4P5sFwE2g62gBoZx
goID6VPJMz8xWur22dEF5It2xjD5MZbCX9C2SNI2QtodiRj4vOzviaIj/wq7JWwB30jbtRJBDMMn
Wl+v0DuckWIiuA+tb5hhamkQvK9RUCWuiVKLaic8eJ/0d0WTALCO80JFLZP5kXvZy2O13AqVVTYJ
WsJf2n0DJ+o/DhPC1+tBNuiD/1En9mxpX9YmlmN5kNSsIRi8xeOxzwMnN+EBL+kgxn5EvFLNrB5v
rP4Riz53q+1KYDX2Fz50fy7rNvLJIac8viRpXo6D3KWfamlqkQu8DSS+Bf/DKhoFYkPn00jMGYl6
pFTICL9uDOC1PE7wPv1rVr+q1/7UFfjgNKNfd+uP7xL4lnfOLzlNcBgkil0HvE+twdXtXh2Zjz+7
PXqGezaxKsRYwPQb4Mkuj9/G8qrEtzpVB+G4LVsCk+4cd++eHgAahL25LsQ6oa33zcM7AxFigsXk
xX6UtJZwBSlGKvI34dAbkeHKbgTBi61/srjz9ve0d63bXALIuhDyua7/IYZ89uQJ9AUyRfIPzVIv
hRu8oyuyUuDTqK+euIDbNiiGfrQgcXGzwsQt0AqPMFYed/1R+dmIKin3Rvv+9sZcIK9xze/8gFqL
9C4heR9tItxqVSVlsS5Jtykv3K4VsEDt/tWyNbL2BfoLefu6/gjXUVmng+FXhszB9NeZ+TL57UE8
TorGmQku/wgXYS8KEVXQW4pqLG8CvnEkEuJL/IVDs5o8R2dcMpZmB+jVC/67VhFxn2V8Oot7AHx8
vxQlgL5h/pqkN/CjHBGicAWPinvgh0btem1rRZZmqlGeKklxlIyDLXIIm2rMwlERMXUKFQetFBTC
3NQUC0W0xdvcOM7nO3ckjPa6gs4dJbDNWfJ3KeH54qyUEcn+e0X0UbJCEXAnoE0i+LcrxaZFmCmM
z4SL2fix9zoVHP9lhqsy53fopBxDoISYLhpKvRAaegucpxW0LuVidrEj8WiqWrDhkBaBAEp8dsFL
0cp+i9sskjLqoE7J7K+g8XDE+/SQtrQX5JLP8IyAU/Vrkee4SDjLrjZGPv+chTAVvzXBCgbpBpdY
bufNp7Pm6VHHJPLMMqPagk1RXO1FSgzPvbRcmGFKs51oQdoreIBuCow++PApW3Qn+hnKQokEvL/m
1ysqpSc16bLdQmODvGjQYqxu6vwP3/GfVs0QiGApMqio3HrjrmEFz0222j+aiuGmIL1Ma1LBD8/v
PSVkcEmSHyfzuBcBU5vLvuQNu/yue37ntkXR3p0d0rpj41+klHev7thmtzTKAfX3RGLv3nz2LsQH
hTM/gcyn4Iqkx0cwKiH+ye63wDSS8YlKybFX4CiecDqjm8ah1+dct/s36eiTrR32xyajvAUKqKzr
+mQ7fq7ppYXqO9gWEdmyYZJ5VWYolCFNYWbwLrUqeM5l1nP3gf6cRQ28cEuiYvnVVE2PiMxzOtaH
CwvG33Inf9IPN/3ujB049EyCsbWn7RpSOaKs8N3kCUC6Hee62M//gMYj0HD7wStTAbl4AcIAOFyr
zqRCrQ1TqZyDDi1aBQ65dmgHJxNnwzuyJ1UrbxKTy9vH7GSpNFBoUxfMkktiKoDQ1b67990FtDZy
9SuZPqepRLHCF+d4iaufuG6Jmn9minfI8Hu7fQMI63TKOV7kmUAyQSGMGYA/BCtkxziaZqEXmWsM
R4QYx3vQIpVzwYpJEXGJ/PzEaOJAPQiIaOIG/Y5iY61kEGjnkwg1jlEwJllPekIx5JI3jLm75PTT
IU5U1m7N6RBawZ4PuMRRDlns40s27OTLgTXyOajcfcem7iSivxzvHVtpjhPVlSpapkOvAX9GUb4w
q/iSEqS9TwF+FF+Vic5OoxtsLpGZvkK35dy/Wnk2a2kiTXxeB4FPB0Dnk1XHeD8uRIoKKWvVkSsB
6gaOSvP1sgdMuGYirOyRT/LaCK4pc1kWCTAQwUgSwfMhMU2cctynUGHHQNfNCSi4BCndRo9i8+8j
696LH4ZJyTDInpEWztTbBBFSJ0WXfzawVyiHJjhcprLe/LvgAKB6WDmohwUx5PsUsNsxOXMI88S8
nWlmjhNkNiM8Y6FSdRyi6XXKlX/9HWSi4tsWp8kkwOjRL/UeTq0o74dDpar1TOoR1/aVmyPelIqj
I3+Ha6TSsR6+0G02MhGxVEtNxAvaMeEX76+gHPJvgmVbB9IeHimHd3cXSVSCceIzHfqw3E7/XLWL
c5L+6YPrI1tGuWszCgwdCqdc2lFM079Nrodma0NCYAJ1LWMvVU/ANcYQdT1DwMd9xMlVOrGfZ+gs
pZYQNy2h/Dtb1qgCknvEnDx5gHbRNn5skkOU3uoTIyEzf35/FiPXs2evstgUTgkWVKSH5Kdt5jj3
fvPq7Bm6XkYKI5lTNr8trNzvghcwYXkfhW9ArYwqZdFWYrjH5jfBZeY1K/9CpCm518ts378PtjsH
pXvg55Q9BQHrUZYJJI4Km1trftrZUhmY63eEI9bvG/iuzSN/QAdOhEqK7CfNM6kNCReI+U3R/dYh
sixZ/tLJHlMtPyZ9ynccZBzW53+AQySd9OBX/HUxlG/XyLBg2N+bvdCnTNZvNypCeb6f1ssS8Vw5
1Zvt63+/9ux2U2CvXZcF7DGeSoBKCHrTH5+SMStvelfmkNrOdBAAO3+TRVary/uAgit9hFKdrTdl
T6MhfhcqCaVgUZwywcjsr44yxYgTmNmA9DHFb9TFnSyhmFS2aqzxHd9c1Ckz34mXDcSaUu9g+MqE
wTWuoX0HCvjAHZpWyzVzbKpX8Coi8PuT0/00vL4yPPou0Ahob7MZnxvQrMH8lEAHn6Ci4pA9zll+
xX82xNE8TjPA6hembucx4UUguUdlXkvIQ+7T3l59JrZp/ga2QzknoksMZGgBkPSse5S2VqV5kpvf
0iiy9gCrFKQVy2DiC5F7ZSevtDbxeAXWjpzy0dOycjgwjypSAixioywVYjrQjqN+rut+yy9lDxO4
gd48UlpvAkNIPXXl4/owUy9AxpoI4nOT03cW8lbrv+hxasAzLD6ERez+1uPqaLG/xhpJr+dsLFr1
4+GVp8s4sp+JpFg2yH/r91M5zLcgTk8mdj+e5XAjojNUQTiVWAigCiERwNWlEyiFjyq8UmoBE1pt
4H5yfZc12RW0P5ynZPVJzbJppfeRurn1ewAjdq2ywDzTr091PUHsL/KZvfziYir1O+ejil0Fb2GM
vYwVdqD8hg/B6YmAZ3rNUYOsZF5gVBUNXnXFUuyY2GscJHu4p7DagGTkkC+DgYfa7jYQLHhkHM+3
BS9C2LZKfvpzunSdWlM4cRCZkffoJIdxorIzC1eFyTJKQdxAc5qnUlKBOuNTlFMsMAfp229ivOZZ
yz0p2azIe61aTytxFaE7AEbSThcxiAtYp11nvivD9TD+VB2qSfAYoYzGSZxHEH9vW3+R1mJxkZjf
HsAU2JdHw6GoSxrxShGKinTxw3HYxndQ3L0z8Wvc1IMzUYfd//jV8myWNVeaNKjcmQf+9j87d1Zu
rVWvLwgDSvJDSjlfXE/Uvp80H9sHBQb8z3cYsM1mmEZI9zTi8fVYgbdO3T96C9BnPoQh1fZ+FQoR
ir+tuTjHKCS8mraxdSfJDleDaLZ2X6Mh+pirztqiJVXdtb3cvLr0X3PkzEf+fjTyvIY+C+SjWveq
wM6GWnwLH7arG53I+FF2Lx5/8DiqnobgO4yCwNGkQ9zDgdq1K3BavgPmjH8rO2HrIZvP5E+QW06U
lSpeZBW3D1Ao8aWPiFxZ2Hjdz7Nsid+Ymccgh+VxFTPuEmljWHdWvbMg+NzigOgV0/uhkuZNyUaD
ST0DVZOT0fxjvQybNmlzc2VVCjMXpl+c36p07Evt3s83oFzXs8r5rw0NHjMj9eJE6UPjhxCuOH65
r4NTYsbZsncJaQK/dGz/wgNTRwK9mXw6M/WcBdnkl1XpIXa2hLjngi0GKipQ40J9mbx/FiIAw2kl
Qz1Of1xOfeDHT2tJqfALgSaulvCgjpj5saZVsbOdypGRTW/s+PRbzQ9WxD5ZjEB7v6gf3CibopMM
EABD30CJoPUc8SyKWxGg/Z6wQXA6tF8wBU140cOBteiX5NKL8aM5+kYzhHfIjE548lGrwS03LsLX
HJ/rYl2mWO7yh8furtMoA45GtUNhyVONCnaIwZFy3dJehPvQi/T9srSfIH9lMjf7aYnkdHDhCed+
vEJmloeyts3q5phbebEYJ1/iW9m6ajka+7eCPN0otyvYcnq+1OkIGHIqGzT3WIx4SeKdNr7RqLRQ
2qhuxbaSwwuGW5wvQj8mRwoAsEW0lwrVFUBIyPgp/AituSfNlOPZFtt823slFFx7P2OBKEJ6RpoH
wWSQMyjBjSj5c+qVIuLO74J+JOyJPAPfR2PV9CM3g0bQBIBNMsL1q0s+Io/8FzyjzvPoMYwpLCiY
KnOAiShGirnl9qgloaUXIxWxJCv3e3HOWlpRcBKkW4EFM31f5xEQTHu4yIzBmnFAl4dwyrBNDiaa
aE2U2xFwT6jKReJPZPRqKeJ9WXpEGTR1R+kox8NUSAmXFKt3m6Fjo5eqEQjqM6nxbKiz1+b8Hbeq
ZLavE8A+QFiz1h7tdO6ZOCr//e+kLUF6hwbFBBJmx76qkDlyppqKVy08/oSnaIdWlJcRYF+TkIV3
4uMRb3bBsDbi93A+S0fRsLEbGqWc5El9zAbEvyHuqamt65o+aDoQHlV2Yh2xS+pngp5jHGW4w5NP
apryRr4v4FkxTKjRpW612/+FzIOhEUp976BbhKNhvfqBgePJPROTeLuImEMOgl+3VND4UiQgYsXr
FJD7nPq+NO3+ZV227OajwfRCkKYag+Mgs21tVAg52TQqrZJGPsYn5NsnriRuWZQGybwRKalCeFsh
aVA00bB3OjA4xtz0WHDt/Ha+2lyEestguPJYhtA94A/rLh8/cMqGnjh7E20tUlcajj75xOam2qii
TgKj5kWfquqFgsL3L6aExgmYJLih8SqHVroLxZHdopCsyFRj82L96SkbgtCG+dDlSfHAHmmg8VH4
lDPYi/nUzmFPvc1vmtS5boQx11H79zJs+jgsx9QJicISC9iTVaK2NfgXTTkr0pkb8HroDp4eG8dN
oswT7IK6A0bvgUVxB81qx7fY2cSJs/7+VuhkGdcFsSxLAyvbGxHi5Mc/lp9BYBYdLQFmdiiEWR7W
7kn+qHOuehxnxd/pj49cIo0gPRHGgh/4f3mXFrlpUyA4+Cf7u0+hEDBc+aLWe0p7knud7ZIgRK5D
BacVgLfxWRVsLubj7rkvjZm1HwC5pN25GX5Gn3QP0zPAcQw33WXK8ttIrROe7ef+bOhdHjcfUoax
8Wxwr0m9uSxab9cFH6P8tIAbNyT6VWszSIb5t2gTS83PcvS0vTR2RKIs04jlEZxuomHmE6Z3d+b2
PKR/vGSt6IOw2SPkRWcbxv7SZHSrafK7rJnJymrzZhpjKYmyOnmlF6P08WTzBVF+ZdHvJbRfIrkR
baDG1tOJYxMMD2vFXG+AsSDi9R5biUrAm6FSCUaGBOQyxk4ozZZiUshIWrPKzr5R5OtDw37Ijl5h
jJUHMbghrA3SFlb7P5hvLXXWAFNkILB51JmUaIdFF8MzUg+JHks2i39AdSwIU94Htms2gKNTPrxr
mSlplQwQj5xU/GZG/OxxzAb4psTwYzxpl6CgmcDjHKp29l4YOxxdHzUmIw516FsUsHtpr4lPHQj5
w8GdzJ4qT2cONKfOTg8w1SuCINSePGghiQDx1GR+mvff+Q4JVaoAznNACg+gbAfPIF/2d1ctvw0Q
GpZIOWraK59keozkFIoG3xmuNuzVpfPjJUyNVajFE10Om3epCs5NZ1ggyTeD77BxVP2MFrd8xDxF
6sG4OTBdEW9fBnNFR7FwDeMwKgeu9mSRXNmiCeV9YmYK/qECsLiiIqKMJ7bh08RKNResTniKei3r
s/D/oVdlI/Z6g3/14FmvdaR8cZa47Stxwqp9GdCiB7YAZtN9U2VKCbbyPxowgfG7D9dzhUXhvIey
8X0Hv4BM8kJaTHPhkmYnlCKzb7nAT+FMmuhaxDwD6qSyg0ODe3AhRd+nvZc0l7zZcphrt3IUckTx
SeJM3TjkGhiuUJnhgK2g97qrepHiTj8RANV3PdFnIu1vXCKXlzQa+cSjoBIGPwjJemWlEAWSug2e
c9wiJaEKsBjFB0DMuS3jxC9ZlRj5iuoeNBe4SJ7iOPnrlwTOvSs6ymb2ITXwNnm1aldBa0m8Fcmr
6jgkfZfwa+XxU0uNNTZ0kPLAjp5blxbjCvA0L3YA9qmx0HyW4XgRWUUSluMq5D+ilOMVcMd0SGt4
QTW8yJikxUC4iLy25EUQw8+I9ASKVN/8B1uVH9bH8I7X86WgBG4HJYvWRhNCN1MDTQNuwPQlO5rK
s6NMrWn2FCH+WcZKJJLzIGmQ4A47oGZo+S7mwOrpjpn3fDi76OsI0spKg31mMlk7iuu0BhcMlVgY
EFUHWzSsxuJA4Yi0ntPjYcZSbgwE27anp1tuHis8kYIJZJGACT2oQptcv/yoVMc5AtYR5eSQ8PzR
KjekazH8Ud0jy69FwcP9V6rFCeKjeQcwc2OeIGJwNCLHu0A7peoSPIQSkvNXJFWLmESjEqbmjj0L
adt6oatoXJrJrAYdnSfTnRb9/wltK1vmpr4pG2zTM/cAZ484nFqdMyJVZjGFxkujh1UMwESkFM7B
4c/4eOexx2xkBMvE2+vq5zD9odZW7VNbeql0TGgh+TvQ1Jywd2aT+ncpyR3d8QNugNdQdrX3oa6J
cZLmeXbbhZ9uuA5516Nn7I/WLjt2gCj14r5G+XdiDhXip90V2f4XOOgmDhmX6PQTtst+7WxQQBcG
nbJlHCszZ//IGZvwhxJ34DfXPRz4Yy79ai88NRQSEw5laYi9ghteKa6jmgAOmeqkHyvDrrCSbNh8
RJWtw5Gvt55uAeGgHq3Jc09ocUalcP82G6MmJg9wWWd82QBJH9xxQtnCXYz7YhRMBdgVEENmL37h
MWntcNVD/N0Lv++sMkzySoO2zIe6Zlwu72OtqF3a7sV29/UAp6cPn+87ZYcnWGTXgA2EuUgwcf+o
eMHOPEq4W4lLAZ8dDcLmg/RSEr00XbxlHkX0wH1AxsGCSzDyBEQz3jUhs2WlE7RPe90cz2lLsY1S
Y5zx+Y8klcE4EO0VemzlveD1x1e2JTFbz6ebsDzhD8HEvgM69cPDd2S0yUYOgCseagN+sVi5sKDG
bvIPkMDrkZClqRU7Rjh581valxgSTDftH+VBy8RofLi1n1YnTE23lkZDbhNrVzDhEg0kvXlnG/1j
YEl8K+z7kK2+WKjSAI9koun2iiR2dkKONcbOOXJP5u8OnPYvLU3M8+PNW3uSDFbzc1SwREedBYZj
eLsX4vH3FguvSiD/ydb5CVqui8aBv7XO66YSK0FdGNQCkZ+CKVswZk32GktsApyM19NkwmYa2maO
PpIPWxkH5t4SVob9NsKMjAKiYtlXrFOJNpzmiwPl3x2vCjfirJMJVO+xFSt+2ciLNT/3u5Bg3vby
MFsRFphXzM4R6Xq0HzpUcgV4f2fegGEQrmfz9itpJv831ovrQPOESyVHyPqeL97HKEz81xYBtiSG
LrOe/vERofODOy6FqsirwxlC6m6SPwGS/4/IKgEABMQrO/qSwQX501y5TxIR3AWMaUAa2r8BReuk
DBoXQUUq4YSPVEJ+bZsVrEEP3e9Pwhfa55VVWhTVewppSNbMLfBleqWh8RaqBec9dYb0hogyrk9B
vVViCBWj+rkk7JalA9hL5PZWiqxfxi3mDf7Wyg8UibATwOyyunoVMs9MjrKwnz2/GsjRAxwIcDCx
ZXgO8zXPzgHU0otVHMu3SlF3D3zTKpHR2tbb6a3Rg6RfvCD9I72wgizHkd2JkbX4vG6u94dJ0982
Fy6VGkhC4gPe9daivpg6cfQKz8F276tFdLesJK7ifpS7bx/hiOkJ/G5jHdVkgFNKXWRfPRfnpmg6
myiHor9UxQnXPt8UweJfHg7YOGkbSPH+OZAliwGE+CSUNPvaBEJHm8k3N2O1ioRsRUNWUgn7X3Ap
v0eSadqPD6sFHxeuqhopC2ZEaah421nPfpPExDx9QPJGLwTJKILpD/USSoB/24ojM2PAUFqNNkYQ
MrXRtOC0O+kE5T3X3g+RJOo7c2IYpRQWCD2ZxdPt+H1HK3y+iuzrgNMPlX8qlSTq1R0VQlu3bk5Y
RhEpkK/PmXlVaFNVjFPRow0yKxWJSbLHNuI64du/fQ9c+5U09TZXMlHqbcwxlxxViSL3v0tHoQ0y
HI65GNKGi7vnIRhUvqCPGWRbWdGn4+CkltzMYbcHCIfwXQkw5iTiTIlUO7u0wVnJeDnhy4XqyWVz
mqeDNhMiH7KprDV/Rbw0JPNtz2nK4sBTNu+Fs0qNvNCUxd5N7Z3Qqb8gHGru7d6++5MjyK5tw60Y
D/waZUq/aPmY5mF22/lX99Wh/Mu8Vp15PTl1IBHBiKTsHQWyDiWMsmxa3suynXiwJjQ+xzIpCSqI
oU2toVwr9UNwdI4Zv3IkjggXWpjYAvpsk4ZqoGGBG2oVIEDsf1xgaZputWNE3cceyP0+x8sLc32V
yuETjhCKjyq2vwp5F5QWeZQZtdAoIzJOoi1m2ppmSVHAliiXx85lqvpMY+P6jmu7Lc5j9PMCW/2f
TImZagEuLoGHOWJE2Vxx6sthWLkUVIZaOxNeMcIFOrx9eRdz7oG75bcuDs1eKPitxya0KiNd5P4B
VHhoBbslNq/7c5zFoynZgwo2UowzOOw+F+AJ8+VbhK0QIN+L8uduHPwSY4AXQHB3iOjUpEIRHrBr
PM+yubDyj4xC5LWgDEn98k2ptJBQlwwthOBpMvKUBwa7Xp+hSgTMs3ak/LUYPz6TL2A8j2s2UwIc
8zo4zGm4YVt08hlcZU+oFf8SWXgCnzC5qNsru9aN/ps1Jtp4Wc9D9Xwj2vzHMn7lE4XTkAN296ZZ
9csbIvyuFAxQWkqSKASpjP/XLIJ/Y3th4Npn3UtihaEulw+OiALlJinRYimEwZDW3gUsZQIOGMPT
sVhIs6lq1qqpYoC46jfz0O5mcUJSvfW1ISSyoVz+PMXbobhIY8lgQMy4J1lsDXvL0PmyiBmTM2sj
NtXwS+z4aML8qkWK1Jj4udzM9Cl16Zw4mkgpsXGJ07LL0Jm28AOzKEQb/O1AJBRTQUCgkXUk778z
ttImAizkKU+wkDz96Q71uvbN5Qyyps0FMAxe9AKbWwCm8FsPrW7HK2cY3xyHis1opxiVI1APC9EW
TPdfINEQ9YiOYBbXLFprao7jTwHFtTbuDPgXvLfiWCvP+2cPgSCx55Np7wIsbwVtyRT4F5GDS/D6
QZgyy+aklCvZEQXam0BleumN9y5ozciMoOHxlTxKD6fvwuhC0jO63hNykslZvpoMj18dNauemy+Y
jkhDWkK1aPYF5ec9QNDSx8MGmx6twwuZIK2atWpRG1/T+oyKikM5pifIkAHbPKjjJXMjeriNfrvh
kCKuM/WpQAzolQoqXKH1VJfHh6IIYqxbPfNsbAqCxfTiwpBSpFLIKUfxsVMwpd4KppEds6MSa9Z+
OAlLX/dcmrBXIGs71OggjGoMgSYdEgkCyCV8V5U33N6Y+ipxcHiDuZV+A5uiNCqlZNhVZPxusXNz
1KruO3tZ46k8DfNu6DbWFrdfkWQG7dtEAhez4bnHdzbQy4RCkHwY6QvVAb6qS9VUM4oO33q6LhDs
QpB9IldxzRh4+cC7ptRgnxJGiHjotE91lWAtR960CGRWWWHL3XAdathceiNEKDXDmkpsO55eXTW+
w65ckKQnuFp1YfQppoYgj2IgZgmbSWcEQdaRQXZrpWQAOb//gUziJMskHqQUseaa1JjeLNz8SSkA
xffr+gv3+cHhR1xO8i371Nv2PB3kvbb74WxEbv6P7vJ0NfbFmC7eq2qouEaEHbJaWmn/Sci5SsH0
9vkn0fUomDPFD+KI3e9MJ685yBCU4F0ufP+7j1SAhPhLd7BraMamhY+uZBh8bICRWAJyX2LSJ6gQ
y9LMLk+66Kch23YsR6FfAj0cQzGrh50mSZ+0jKw4UNTIxDG0zmGkaVvH8qtKMPd40L4LwFyTvVlb
qySSUPY6RY8GPG8qwsnLExL4Ey7FjUSFyRVYmQtdJfDCwUJhNoJ3tE6s7mRkKvRxy66db5YQFYuu
W2pj9ug5xBHa7TLCO5yRtz7n/LYpb9JQkknaSJRdJJ1FTeLSeysCTSzJoCvu0M+7KpyGtfvgCW+L
E4Qhr+cM1lsLExRN0Uq897l4a0zQozexbQ684xmmmPoQBbIIxt+2Hj7L4NGrmpMkAtnOVGsAnPmO
Nn5UyHTH+0rIvPGOVc8Uvst6Canr/Px5pPwuxR0big39g1h1O8AbNOSk/gv6UcH1hD+pBLxtc58W
vkrcvFUiGGyWwCYBpZ0E/qnpUCcqhJRoFS79KDam9eqsskSU6eiL/JHmOlijFKGT5/pvV2jxAXmq
SZDLoUdaGJIgKNEE+78Tm5hc0NEGSWKQlxZZ0J9+Lg7RSa8LJI8YdHcYYfh9iYfjnEGkwGmKj6AT
UhnONQEZLtMkolC4uVhrpR/PuW7FmQnb5tfr71BlSkJ5v3tEUCKMojldncwk/sI+2EqXWVh4wvid
Rfs5zIybH9vY21YaFjNNWI/qj9aMrxhJe52OjpXsyAw/89fipGzD9zhOnihNBo9gFs8g9VvPuUG5
zOxCzMm2NpuK2Rz1BFuNXPrG2w3fDnGGOtZjwdroA+Wa6dJuGNRykkUPRpk+E8IJNByqGOXYG6zC
/0c+HfLf6rX+uexw+x5GXwykwy40EK8YuZ54P4MJwpmE5V2Ie71DkcKYFV2ix8msDZy5C/AH2kSn
p5RjysGchsFmm07vl94ycvFR337ZdZz/UqDh8+35rgOYCv+bALb44GBe/2vsRrL0vld7KnWib3tW
anzFJ8R2IvieiEBeDAj7XAk/4wCJXRavq2N+eCBsv6shvr9afXo6iWl5iPK8fvjSDpnrEQ+ovhkz
knZ4lYcGjCWWUi1/ZSjaydBrKWe8aIxNyJ9GyXyAm+44hDaPbGDYMBGWIMqP6GH8u4+xaCw1XE+p
uJTrNJorlZXFQ6wq1pyQvJYhXjqaIQTe2qTKyfDsLlGrqU0x+os7FjIT3Xa/u4eJ0Il6rpXx1oDP
j2DLFr8u0jUK6ZP6mo7n2Cf2JakK4Xa1W34SqMyhAdqp52NFwgfPx8gv9PjTXLXIc1UUsZTzpkhV
KqOZDKRNv9Hsq8lGW3IIcRMk0iLb7IL2MZsRGCofPKx74+ihpU3N+PCuey4Ok2oqYE7AidoiCAzM
3yvVfDJVaKoGHaKABdghVnF01Ng1a9eFYxJhgzr/OmYyLtgSCc4t4PatjX0SbAoAq+N2bOr2plYH
1LLLEidM76ng9I5JRcNOQBkSYBxQp/Kr/ptdU8kEA75ES8iW3q9MRkKeHPgOmDwL3J+104uJwDxL
X+HLXiGMQOcST0SukSZZkH/HxqCJOF2FTouPJ8Ka4tTgR+QwLlqmSg9j9nQLkdrCya/d3dg0U4tY
nelArMfcUEUwQIJnjaOyqslBivnJpFLO675ZhcnG9EY0tohxIEfhMU/Oscs/a2t3jgCxD8eeh9af
+XOG8AU73QZLRfpB9t/Sp2wagTB8I3+xsPCt6df8gl1oDpXAdksxVK3X/Tc8QEzgXlexbq7m7Mnk
xEleBvrkq7kq+eL/yJLWXpahrbCM/SikOM3kPKMEfHUW9HjpDUj9MYoZFxcLTzjfN8slIsjy5zDq
tyu5x95Kg8cLocWKbg+QHYj4tg57oWWNWCtCTzZhQPKQhH0yuPEZ496gVm4xD6AP5TQC0nsEk5Rw
wv4fbYnxeu/8q/HDLUlyLUwLyvn57p5cWcYjCcwM4b2MpXzyLyksRGHf/V6Q48EJOpTWVIH4q+RD
K/l4riLVRswpzbmPoOVmEnGi+nROOl0XtVWoxZ65gb0mv1xPbwTX6i01OVxyWwLBUexNfYa2VYGF
cwi7YgpIFzJuzUtf/JOUvzsKMo/iFXSB9NJE94UL/+D0ffm4L90aFSzAxQL33rlLjqk6RYmGz7kI
M8cGB4NgWbljB0ub41n59xfdQelzZ0ZeWioCEnLsc5WsmOqtSzhjauPeMF5+TYyXD9asgTgDCd4l
Z0e3GNBG0BKFe9C5q+4xmU7Lkb7OxfGVpIJMdnus807faGmD/V+Vw320Duf5gCDkgP2j3d+SHmJw
776QKKk08F3jzQhaA4tTxRsU+AuAMfAEygxoBGl2/UdCrl7J4nXC/6RshTGxer9dQldw44CXP0Al
jq14I7j+25jyfGh5G+pLs/mDtLhNaW87D16ykdbicJDHBr2hlL4+X6yeK9LK9Wrd7qcpaNhDJEGX
2SwE7wQuGaAhlupDAX9iKKWY1fKpEwNXEBvppPX8Z7kXUQVzyV0Mv+eC1goCfw0RVLdgX2EfQx+G
aKOpTUTLUhuzJBWjtLAOTBl0ZvRb9nDSBxvW07+o0IXaciWPcUgsECPHdxOwXnLfYz3V1oUp/YzS
woNV5eYBYt4izZcBv1aYQDLw2jiHO32wFb/gRWW87Yn8LpE8KFGPduAHECdCyJ4Q+DHSPY8noafF
0ZPgjs8TjEx2sL9+ErciJHFyUpcoasK0op+gAfvQLQPvCGz1tyh2Lm3aKzup7yEkjnvNeY+YChNR
Zfe7/pNewnF6XF/6Q/B298O6KR90gcMeKe3WfIqJ5ajxwrYRRJ58pRZzNJH/BycIOqzdotqTc2+l
FqswirFw5kn/tO49nMlHSq5qjjCL4YP6F/lE09HVEUoCQd1MgEeSiSdAL2B9H8CvBTF9ceUfTO9Q
XXjvgx1j/6RQMuAfoJeOI8y05NnjeR9W4veElNiPtPqk3Z5cR+8pGb6ZxysNrGAi9uJYoRBeTBvv
9TTI1FsOdhOH2Y7qnWY7zMAFriC4oOeIOr17m+VO5gPqVFw0YSVdAtxoOXm5rOrcJQ3rM7HHf8AK
N2asdJlGGt9n/S2nxMEXlPO6hzbdPcx/YakfyAzV4n9dTgGtEOEAL2ct4Ug/vHWuyGgaexxAfnfO
5Ja2iQHTG7QABOfqZ69BDbl/PicGRwuezdVG5lBI0F6IKH6ryNGEFc2VqKJMhojxcfcbSFUE/OLy
kmXuRT3LydnqTUCJOY+8OBNawFt+KngZswZUn5rKflfOFIN8fzl8usOxbBnA0JTL0Gxof+CgqUjV
dJN7B1oJqJqzq7E/lmsz5YZ/avhBChBpEBfQf2ZpTq/x2UpiSjmd3De01U8ppdr8Nddj7s5Z5toL
E8uY4LrwDmB0yO3eakJ6/PXNEy4Ue4AAKXK2d/LG4cOACbTwaIPXgU/oo3177okmTVT/A8PfQ5MI
2pdUMLmP4XdtpI75Vm2jYTk2gm96v+dgnDPfwxFeh+dNxQ/hT+J1ieCCtQ7JsoH3UcQGHlOnfoWh
bWbZ3GnOloeUZag5DJ1hY1ysq9XjmF9HXE/zmjBpCBw37em/rPivNVSVpXsnbvAeTJCxHRaRJddw
FKEFZTQwGUhgC0I52E0z7LDdde8rXYkmT55Kx49pmcBrEXJgGiAa41w6HyUNLNnJk8X16bkN1HA1
yRmmiaRlqrs0FgbGW/J8s1mTwyuv38aMBHKeAvPAd2Q9mSFIzBZGPcRX/t34pUGhxYsP3FmjGnv8
+1M0Ilo0143/dprGFP8DEwScIhOW5GGymcsIJur8IA8DjtFswPLSj2VDl1jojEPsqLmpXj39b62L
I2XMC0imLNGBpqMl5ff/Q+Jz9jbP0FX5i5GaC3V1fttRDswrYyVeVKTCOq2lUx63uQ6pzkQ1lv6K
A3hiJwhkeBd0cAvKIeaJ8DRydTUUrDjvjwh1p1yzJry79lg+qYSEpAser/Cbi5VDPlkWcLgi9aZw
fc9JcQ3elnwic0wFkTP2KHpJ3sFJIeocGF4GsbPlRA6M4rx3l77zDcNBHYdoy+ACm+JOTCYHMVHs
FTQ3rQg1kVwtYlUlF5fDrqS+0iWlhyww2mqiIYzAg9qwxesFCsXRc2n0qradTWsX9gO5H3W59TkC
EwVYvtTFNttJKH9jmpDp06fI9Sx3zfimJyE+ic2KStKAj8c4oZsInjRvWjExqC0BS3vg/di7QRi7
ZPz/zZ/fkPMygju9gcMSYzwh+6pwVcCZM0vSIxTsfotWBpq6GOSgLvoaN8Y97mpMnuiW3eekb3yH
2CefpXUIK1AU+mj/8DL/h1RixX6+Pp9aBZaDmGoX8SpVeIcvGytsgwgiQ9n4Wtj5NLd+PfH8Z209
MKG50O0PRFOJbkH03WznKkMZUikeFA/9hkfmhfM7EqYqTQBR/9eFD8oSXTZBVU6XBS7kR1djgwia
ZIBjAC7J5Tiq6GX+XvpQwKeVvP9m/9qTVyywsvbB5lzDDpqMlNGIbH4B93h/wJQEiwHRBGbwV9v4
oBpqTFzW2DiDgWi5ZXs2kAkS9jYQeCbAhCWCCeDen65rX8bRVlxfMONlWKZT53r4k7/ZNSfdY3VP
o8QbT9q838GtCLCdwkR/Cy0zv+Ccg5bnnmQH9vP5xRlaGC+BKt7XulyObfTLxC2VCe8BcdUsSeki
RaETcn6+W/jePGIP9rGvZ5uBeFCv4+svqqgslDAy+TlLlmr165/XBHsHq/JQ6Yt0YTkY9f0tYTUd
dX2K8dFhYSvLBKv7PGYF9w3GDMPWAbWoV+Mb9gX68vgj7VM5HwkW3z+XLn1W9yM8NllSl13pYltB
rL77Zuk5uUtP+3FXuRFRousHKMDYOSVKm2vTclFqWCSEH4Osz2YQIC4j1A7qeUCiSW1ai3s0TYeI
L/Ig0XABtfINK+nqYBDMwvUdhPBCJqE9G4LN7vD45uQRXzQMXmSi0UodXDAOJb61Awo1jBkuKIuY
gywsNn1cl8pdH5fn6ffGVwFhwVmdFTP67chyqr7BLp7MdHBVfxWDkrBLC8x/lfgISCqCrgvilv7U
roxF16w8GwO+Fs3Oz2yfNa5crT7lKoaduQLnuLgsf8JdOc30DJqXehpLw5v7BY9v+ytQPC3YaRmk
zoMmBDMfN5nwwMnjcUpTa4h5Ckxv4RtI30d91OMfDJ0q1R+HyPiQWgu3nRUqmd5VzoGgwjpUSYFc
nKs/Rhk0XPiPhixu5LlhpXrjG/t8UQlfiFPO85UFHsj7S2tgP6knmGgggxeae736SH9qMvVaWX3d
XqM/PpwH/By2sMFZCk5NpoT2IJ0glPM/vbxMJEkCjM+DZlNS5IZNa5BC1O9FGi5exfLXU2P6mPMV
EQRlnXm/oHGVByv2r1BakZenNY/7mNE5UqQIGXpIQ+dEvsxssQAYNnbkxjSkLn3TDPsVAQU4B8Z6
P6wddy3tYfUunmxF7Uz7afF9SXi7NIUjddVfP6bkK31UVytE0drkq/J09VXe6yrZbY8hFVnQ19BY
iPcv0iw3qUQ6QQo3rDEVlEQtJuTJn/BpOelC8Cpb+Ddm3rTvIQyYmY8eUzI9bkWK0dAxXeMyHZ8y
T8ZxNlGDr9224XFhGnCDPCPGpxghKi4XAW7aiJOWcbbJXk/P9rFIK/XHDh1PsAduYoYAkoouTmcx
ofpQw985H5l2k3nQIgy1NDex8WO9qKoT3duK6KM06Hi2mLRJ66SL59zsTj+Lq6DssD+8TG3DZC9j
GLZKfeEc43KK7YQ8BWCSVONcFd70NeYXFDM7Z6pM7lk2NxMTunnQSn+9QhWOs/RPbt5yuu+vF727
S2dWfIj90qAK2ATc4BhNH6VqzzjmdoOBwqMyBgcoIdGaL6vKsYjy903gQHoW9Dl9Y/96LUeFJvqx
+BeJeUQPpn6OLEZp219S/j4pZfIbNCdZ7xKEVWa4zrJGFqibKg2DBU3mKfMgcZ6VzVT9q2wjy+Pe
dOtRZr/PRTOhY/yfg12RW34tGQaAgCBD3wSvR2f7iT7/7Dj1TsdXf8H1iiautdRPQmOzRGn9dAyP
cR2efGQrRTzB+NqXD30DK4zBc/nzD5PdozMTRVprhlQRCR9tOfZ1KMzYa/w4mIES45PNpIGZ2UOt
DQcbOjeGm+m3Ov40K1CwW3kbFVU/o0cZEZuestxK6jW+QRr7FkfWgH8nKMKbEtI9edGbvZY+urvG
AfePWFYiJ27Q7rVQjgVm+BJKjrpoSqdA2IdSqhwv5FU1/ul1Ixuu0pZELgYyjpCHtK7GOXD3yctH
nSBw3c5gxNkpS7YWpKdibYTM8hOfut1BXtUs627bv6m8IENGw3hX5sLIxLQxtzrc9x4ZF/ASSxvZ
uuralRIRDIuuIlEzJ/A9y5Y1WiE23MP3Q1w1E4hPLGy1MED1hQUhgwtXdFiZP/pNS7ZLftIgA5SJ
tAQynCx8hL0XfGFeE2b5ONKs8WifuxH6EgZCOv/Q+lDJ12IOTMe+X1Iyum71AEY7vTD7CLeEVrlN
Ct4BkK8B485Fgo0o61NW/KKpQI8Eyf6N0+GRuWsJSUoZkim5XIRMLUhnas/rQ+GxFwdBWgI6fYyL
vO0vXTilTpitZsRub6v7LJ2qQL9vOABwgOJH3dDHpyMy5AKnF/GaLlsvXTcV24uuKMKLNWmdK/CE
nxy8Ee45leIVUzdaoN6hGDa65MnIHkwV3OcBzEezEXtN1gJUz5wzAcHLoCqjFwSjPOFdYLLRG9nl
FRsnsuXgGC+ZPkJyBwl6WFhSB40WYzNcg/8pec2qM+e2xY9VPxxoBpREdgaVM3F2JNvrODpBLcRw
dRxsP8bMH2GZhIge936dWclXDaJHSJmDNdG/MhgcXBwx+GCGsCW9uUXOfQoPeO3womQIucFtqH6O
ebsx0ACAHDqhlrzsGSIbmt+QdDssVwLG5gy4ySBFn3oR8bchGW2wf1M2iZNjQ2w76hlKxRB8Kx2R
xhCrdwcbPNUlbb7wi3sYYd7MU8TkFyt1BecL9ftgmuq3iOq8GgMjMmZrivTEBfuLUVeSCRYLoY9x
xvHmlJFM7WIrND25kN3c/J1SZoG1LVL48DCUJpihWVbsY1c3tMqkD2bTOpOvopb54SA41bUwZ2S+
mIiDylgd/aMXC+8s0oyTec/jq55wKCmxljznWgeSC8hdlqmhlaDfGUERQXEAbQx3WrGiLSE4Yr5+
yv9DhhEg/z6GSPThZOoeIqa/faXdTkSrqJ1JCbLU4H/BhTzI45SOGE6d1IJ4ODGkSp9TIu67Ukco
inPpm375HUp1Ur8IA/63md8XFZBysmtEdmj12FEzgw6TGSjtaJg74O+SCAUykSZG0snAVmAOExhT
8oevNeB2EeIBWoMlzZOkmNfzm65i98hEyBnOXxxMEkyWFT0RLIC/CHKVcuCZJSNJVKJDBlr8wBL8
6NQXf6pLNh0kr8flrPVzhi0MwZiXLiaLXqpIkFYW0tTshdNhqWavZVJ1tkXxh3mVUxuHZZhgqdDc
/q+Htwcl2ig6RZzM94A3/xHRcJ3y/T8bMmqIGwWTPeKhb+btY+jDbKJvmX/7e6CO236kv6dxox93
Kg9hOQoQ5J9Hu11zphp3PmV//NiUEOIkWvqv/TsspQTzcNTd32G0X2EdN6zUkXS4H4sSOyBVeL1d
cxW63KKHnf13MqY4/f5EKkd5eAB+pGej2VSiTwS05r8RRw1wE37A7hPlW5kNtb8JYGtP8iafaU3y
OvuPWXYfu3CQ6ydsI4VHD7fqfyp7sE0xg/O1utmcuQdpseuAVseZL7ToGrtcsm+1pG6ZHixV5hE4
IzFhz7kCdp6R+xh3FcpoVGdD5nMtQR7WmxBbQbMc53m5D5N6NIH4+Vr3aRXxE2vy1QRjrwmDPjEs
UYaLg0buQOWS72PU3xT7jks0gj7661+Yt3yIHwSZ7wvGjH5n2p3JP9jzlBzRPBnN8PGndovkM94f
rKtAk5xo/E38+JDzHHkFF5TkWQ3PXCvdSs4zcZr9Ira7F7dFH67XszBYPGoFwhNqf8FXyBBt2xps
+DyNtlWJYX83dFRBqgapZnxnl+raIfw/qdi3q6LVcPs+SJDYeuftUnRsMhHEgXZD1kZbDNTM5tgd
d5J/BnvkdlcXz6i1HCHijySnjFOCbbghkLm3SKC/pjgib0hCNj00ABNASK2XazAfZgzKj5hK+fqW
cs+Z3vqldQkqDQtwEnLfGZMlf1EQlM7W2cIoopDBF0eDhOchK20CeLx7GCN0o2F5Jc8lz579sWSK
APaQw3/81Z2IEfwS3QM//w2HKSfCA9mCkDJDc85Wg69SHLiw34RsyQOkBCV6P1s8KsJ/8iijFX82
YqzkX2gvIL4WJQ2QQeD+FTx4zzjtjcG+SB3VNWMM74U84xqQ0sMZuxdsOWuJ5kIUqlSHc8xQXVzF
dtbYPyBDijNUwgAfPO5fOXDjU7zcvsOLXsk+/o22hOYrnFFvT6+pW8iT9GfpiWGF6Vih4Zg3rm7H
WXXmg260dDx/Ju0TcyITmbJqBWmmtAsbhwnv8ShTkaRWpjbvVZgmi8GhB7BHhotzazBxpKqDWE2S
lpeNW56k73QtZT00NDD7nECWrCAjT7TVIaHaHo8xTWYl0VS5Vx3rv4MvPDneE0Ira6PLlo01E1fp
SIu47zfXySG8jcgqL+VuQSj2Ps80opaEJI6yw/83jC4i3o5+6t2LrR98QqkHQmpplrGrSX2wtIP2
VIOWPPv0565PtjnqbAbNwKmFKdzBoiztxcb1J13u2ayJOHtd/fKuCqaBf5ZweetzDECEHT4gc41A
svK+PDYTru7sNYuxSj+LNyZnhLbkpp7g4s8Wgo+3KV/vMZyqaVEPo3Bfqo3RCLCgABzD05WlPzsL
rgeQVeJtwsh5TjCXL8D6C9NBCw+Kko2RBOF5CwuEKOltIMPt3oNJcN0owT4HNaUEcGCyY6fm29KS
GL0FF2IMnL23z8XP/fMgQZOV9k4dUQ9Z1/9109+50ESYTJ7aYA3qwHgSdXAhSY/rHPg0LEmXKk5s
1J6aqcrIIFOp5QRSLEz6TNx8/XTbQrXHlSa1PnP1bpN1GCwEVn4sIlQJKNLQJV6UvrjAZKdSohG4
4/eBbF5wivdvBf5UAILq7ijWN7SP4thkq+qR6cc/tDUVRH+Mlivxdrgf9Xsq8QkHpyIdRCh5YrSD
3qEbxfSdY0qQndiMskcuovKpirMIG8RRCViKh8eXp2n9SAV9JnZGDze72GcIujrpwf4PdTa/1B+G
mB1QYdpkUIpi5Ejsi+B5oFsMd1ga/+8Mrhz4b/YGYIvHoL4RLDH2UAiEF9C2IwX5eGec2lcrTzO9
SBS3wgcHp70DNfYawrQpIopw3NVi0mmeR7gZ+iLIhOrxJVKzkt3qE+jbB0dsJoSQERzuGiLamnj4
7HFs7iIggtoaDtaN0Af6W5wHkONIxVURuG690XJOt+uXqGahL1bLpDkGG9X6KIMU9kLY0rEDX0gI
RmjiIcqW70gXX7/uUjWebBZowEu1XdrQe800f3YUTi2DRwbyRV4M1zxQnaf2i/QfZ9Z2JXKzdCNH
IDz73XBr3R7uj2K7F/BtUVUdktf96y4rJkDb4uCEet8kVZ97zrTp3+nL3CRvXFGFhdTA3qUJpf70
lf4LDTFFspSyYtvFC/MdqhChHm5z+mXmKasaPbyhE2P5ii8bVsTUKDpC3T4vDWl7HaQ/HbbhXhBg
FlRepG3GY7tJqQFK2asD7h7VrfzUfmH+3p1KaQMQtEe1JU+HiVkrHrBxqc4V99ctCveElcC1UrkV
k/KZoBPKLi8epRzzZAxNO3hYDc5qcx9IbQGai0smIKQgng9ort5Z6lMKQQzR3lr69oBgrBSvzSWU
AqBxDm2xkD10lxVKbGphtoZGOpDqPeG5/kIv10Gr+N66ECDuEnNgOcY+j9WsVKkjYrYA1r3tOlCf
2x6xf8MaKTla3dRg9O3ZAqU/cAcMsp2xFJUAfnInZ+vGuIBQeM+WPFW+itYcEbswTRd4+CU7m1a9
vBKzxQD2FmOCGdM0XW2nobmgM9Fp0rg/5GdtU73xmIsrRAf3+vzXX/ALzwdf0x2+nPLESk3EX3cN
m77+D6oWj/0RLKlMdvodi8EQ3QKpOw4F17uAf5XWc9QdJ953TzbkbX0LuUTeW40GqdgLfVVOJqV9
/W7PevLG9broOVukIAduL3NQkpca5JrDYO063trc7xmkNhNtRvGNqb294KotCYu16oZo9EoXr7Wd
owbSW8/ivR4zJBKr04PC1yHpEcgLO7TPynqlVs3229LXP99ca7vrKSBB+awX/7WfIWqy9ySJO3ic
9JnZsaNyNCM96pF2Vhq8FoTbBdBPQ0+he3bIsDrgil98z7QiKMTzNW3InE/0iWPe4/T7Umltb9Ic
HjNnTgOZw3J/Cmv0lrlnFHlQq15XQs89je69RbHTGbF/aW84XWqpQrQzAlq2LXR6drfvZTvKJSSA
xRWeub7hqgo+EAczG53et+igY2GLivLvIUBagAaSQx5HhIWS/UGwNHDkcfTgSZqRDkqFDcpzBlBI
NjTBmOqy5pMx/kC/4PwNFba2n8GCwHFu4glJe+GE3/oTwN/2pGHG5+4cdfRkTKi/1YgTunNXAVV6
pNoDvpwaNsvZSa8ByhbsQZL4HpY75wrPj1Isv6z2zreG3F/8ja+oePtKyriDqF1C6HMr1ZNMgqkQ
NWqKohQqqbkzcVc9qsoxu0ZCJ0WOippR+HiZs2BnfzeKN4f9UTyq4it5FtxnDaIUT1Jz7N7PxVL4
gmflZKfbQLVJMwWzij7RGzmjwBqVkX78EhrZADgXWVIiJjfVFIMIfQcHBKCJZAU5QqT4M5uozyAb
U7W+46fANgLspvYlQNOrGZhQxHU9wuvv13Q244sp8DKRfCJ38mNit1/HJCCF91bLExWZEOtjWwDr
Xx0d8kwN/u6/ZviNWYxQmdUXNrB9XcFqq+8EUJBG9U64zh3U8vTehqxEBoAEEwbM/uv3BIKe/PLw
5qPYuYLAjSzyMI2ToeAjjrKzSbhB90I6jxOmVHgHGlF/xcL4T1YkWZimtWR55Wgex/cMrS6W4+f5
0wfS71wN/hmyk+1IzDArIa+vfOIQXLx+96v8tpmejfbAJKlCuLj6ueSdEtrQ26CigT8j2O378Cqg
3YdeW1NT/TL4e3GFg2+xFjk4eY1eVwVYNSJy3lHcKGT3hehNE5EDPIAhKh+gmLQ0/j1pt2sNOkgr
j7SXLGhrpNMFrBHWoTNdHYWYfuze/ZxafmMxTrHMjPGGBF9506B/yYyjfZzMNgPlqmKnTrizUbQl
UV3d08DbRpo65a1bn/wK/tdj+jCWfUbnjCiGn+FpItt89uEm+hjqMHDp/wFIx43szl4qAMyNA/jx
QCxKvp7sai5rysnCCpbSTtYN+g5Dj4p/PR5G2UOqmhP+zUUCS9wnu2JUbXbOPjWJASkj9A72cH0W
ByuP5MqmTXufgg0I5Us+lv9FLytkavAsoveDWpjbAdXN+fVKXOIoIpTm+OQyTTtBimTsX4T/4vC9
GKvuLwN6Zh34ku4KqPcYamKZtZwEQ1pSvNv8ct1ogmghpd6LiLSuAQZ3viY8FpH1HPCv5yiEqhdY
gnr1jAiQVIfZ+cjWJcJvL/MPswiGut2R/VISU79eTXcMaMhF1Ne5u5e1gV9y5Mv7QkNZ1R8I+i4N
m4OnsjSOAgTw0kIGE+AsPDWyISDosgsxPd9nV0dub4VPT+hx18Cskf0RpUo6QDwTwu7cVaV9aIfQ
9nLCVvU/kkYybYFM5222J492PjzPDRhzX2KyBGN2+M3PEqrI4C2mDbqTOX9YY/H6ELsaJnqf5vsD
WfxPzX4vOxj5iQFKhNwYmHK8eyiL59N2R7ok3dxrzyul6kqmPnuiVj1IpWIBMUlNrbkiUkzdpO+x
kPc8RE7WeZcTZ80ek5uTNFxqfwDLerwmXyPokR7y3DyKc0tSVOGImD35ec1DMonCidFnpv6vIH7+
4Gq5oJwXaXJZiDUnLI0ORRKTUPpLfTpXJ1NVyjDImahbyp+dKAdBK/W1gOUyzBWEW8Qhmj123ONR
NqC6+SNGcMrMr2nj8GiHjIqv5Cu4wedODTZvvbx3Qpd9t+O3ZqltFHQ8QQ7ESi/OVfSxWPZyLNwm
e7K2HWH3lBWbUaJJSXfLD1WomZj6G4tMAJx52z6CxoCjMF/zKXt5lOYZeKsosTj7SZ7F2S4re3Is
2SgJnInfgcSo2++qeUVlk/A8J9Vd96PdrghSArKGbnIEigMN1FoYwF305XUMRBPaQPDaqD4DRIkF
oORmMsKANLo5jaDPqjBjxRYuIAr0U/NUdQEuVWuLtux0hGrzD70TIERFTAVrTxRuMWuA1KPGl7Ys
+C9I2n9m/ptMDmPiEyAvLuYq3i+kOyPf2gHLIBcI3TYy0QkdOryqvkrikhd6yb70wfAjr/rsWR6I
dDMVio8wQtiUvG+mwOmDXDBL6yD9+lbFyalEbMzzNmMA6YzpXTezkVTkAPRA71qeKNd2lHGcHlZ4
DxIfZeVPg1qMT4yqWNQ6P2ZgPSryXleMm369gKqKCrMmCXOvzvsvLCz162lHbn2E+B/knnzTrzT3
n+nZveJgAJ/F1K09aS6IdaO18i3b4wGFDsWmiiqtrP4oCOc++FZ2qbTrgMbyhyb/rvCqiHbSza29
JpzEhOxPjPHzV6PmHQk2YJggwXP1l/sJHJ77qKZaMccn8XFSzd5DB9ro3ra4trR3ASma5e66eijj
D9ZVR6oE0I/UciTGiOdCfE8+E7xvUnYvfwG16UqoVpbaumox9uC9xs9aQ4a8TIjCcOA/sk1dgve4
XN+mhtYCZ4AXIssNwsnIyvI2Ack2gL2ItFTwytrIYkXyw3ru2uskqhL6kk8izv82yFLOKloxMVf/
xez0sPLP7axxq65m+d13/sA7uWwq+sUT7y2M/0yjrcTJIcwZcORbqZv3/KqzesntEuUGPp4J6xsP
yko9ML7Q4bYXMJz2CrdaEtYdoUjJaLln2LWgK5LT3cA/EuX+ioCi8Yj6ThbEus3Ecigyf9RPCAgR
otWibDQ/NoxIJIN1LHHd7FTX6ItkDf/5h/ui5KZzX9+Al+bA+lE61enTbm1FRIv4ic0OqERCpRgx
ZBToRoA1CUwS/eBDDla08M6mYwBJ+NFoRcdteR93wyGoN1F6HD3DdRwRl0uNLlJH6erSPCLatVAM
hDbUL+4FwYkuyrCISf5iRgnz8LFdrnn0jKB7uyYU53QFa+Y5JQ6WSmsjSPWEq0SWC4OzZ33V37lt
hIu/lO2lgKVB/Scv9+y9w+AUorLFhp2/NgtDsmEbNdIwqUO7/mBrsCF3FU/fGOgG53lPvSj/0M9G
nYJdDUmnh3DFwAhcvX+AOV+mK2D4yjo6iXjTkq+nhxT0E90icT+H5GDDH4L+qWit2lVfwn3lcPXd
ZKCAAIoB5xyos/uSCs1NML9y6yQ8CYL+RABbKM7pYQx3q80suwTHs453lwUeuUEsjwlpBF9clOA9
wuPV2Du75uaz3vA9ofCYGpjopNfYEBKYgfARdKXOrZkRJyY0kMaaFoIFshBQb86QMhWId2Oqzhb2
MYM75nYMK9Xxw7sAH65zmmamQ6JkC2hzAAZGI9O0KqC6G0yGyRvbpSilk24MYp1hcAp2Gd+A6K7c
YVmKsCxhnflhmmbfEzOb3yATFG80lKzo4qdlyK4d3Xx3NkQb79NVfZ6n/ZqA8+F3tGWSXgJI9rDE
f1yG8CG810GAMN1IOISIIjsYVXGTQD6Gya6NTXT0VvmB6+7f3nydty/Tj/8pgab5G5qtdj2gOM1x
2QhLx6Op3f/t8sXr66dq786rRevk13jzNIHq6eSP1xZ4e1Eno19I0t3fTOIzeJkjTa6EDvIo+Ldk
gz08XLQ040uXhEQBppwB0lsiagyRYDMtGixqsqdtexzqJ5Y7+PEI1nMssdz7nIR6hD1Kxdr66WWR
3VLTvBeyOKxn56mzO362lQQboTepmc/E/hfEo+klj1vi1fA6MONKwm2Fn4cQU9MikNJyy7VsRk8a
7elc3pn3lq1yDK1vOQQ7U8KRTe1pMYDvNeM7P03GQeEt1lYxWS9dLAS6hT6JJfieqE7IF+PLPdsP
myHQWPg/a/ENN/jPRd2zM7C5x4yQsHfE2YDkab2DLWYGMeaUQlU19cg8qDWk+2Omdi5PmrCWnJMB
cwJ6rBM0Ki8ekD2K7g0aQs8rum+63XqABw/BRWW7RQR4wLEcq6Z5NjFA/Dpy7zkLK89QC9UIRzdY
8W8ViQ3j4uLFOCbriRdl05E/uB67ZW2b5zV2prCgoUZukRu/r39KfpOeEr9nZErWmI4s5D99wnM4
21Y3venxLwMoY+3/n2jRkHroyl0XBZBPNVZbV5ZNg1Qz9k0FRlG9agBqSJJrB4uM8YxsHJI3y+FL
xesgfUtq9sErPLRtLIAxI1qT69lY8PjxgUOxyCBvY+t/9ZsJ4KWhIr5Qyp/mgQ5VY88uaKGU98/2
xX7lu1kaH4cKE2DOfurNeesH+pWv0SfN4JITvDae5kEX+h/wVeDBkYHviH6xPRnvMAJQBn69hFnK
gDszp48kHpBdgr/2r2kTBOZnfWX3w18qUvKNJNdBrWAfYUVbTaQZu4H3DSABEFrlComnHYI1NVQA
9wsEzBWwjnw98oeuscoV+eSwkJzRTF2RdoatqanARHzXNcfdu2mXSTSTnSOb6f34n1i49bniUlAc
r76DSwyRnG22whfAgAeYqcN4rlM456CzVAv7ITjlFscUiwqdUsnN/Hy+BGU/R201VOIo/br9gdah
GvFLgieES19/eONgkfrxr9zHAD4V6OZHStAhOX6rHOXqIT6SasfVaosEsUXVNrbhdYvtZgS7gh94
/2De5v4n+IKM9Wdn01AqeFCb3fwymoZ00uQgzwW8C20CClIUZfxvQwk0zWYvqD0EZAkD4LfkCgVW
H0Ihd+khwaMUp4YAG9wMwGr8Phua+yxd9awDblxaFIni66/QMeX7c5Pj3kVMUo++g++D3KJvDaDy
Q/tXie0Ri0FRn2RG/PRCJgdPykla3EzNLFts54GysYaqw1oYQJuSp42jgXSj/TUiAxhC8vf+Ygkd
8p39GXPIFrMDtIx/3zCgaBcvZLM53TJPiiruGQzpTDFG+dQKD/dTzYqaPUuxQByP3YrPSG6K7SJh
JRky/fXshfUNH40+YGOBIl56XjSHm/Hl1ne4bI2i8GS8ErJCkf35wzlHOwFGzPPbZoQAzSpsGDaI
51U6NzL6KyoT0pvpVdwhEWkv0Vj2BI1jylgqISz11ZdKBmNFPFHLPaZ9MS8hbQEFSipI08XgGOB5
dZxJqA6Fs29d2SyPhSOsB+/DLv+Rq17ZgQ309uaYZUNbolpNuyhVCfAgk1KPJXWag2lRXFTXzt00
+boeDhyich9UL+X8578EKqleeOGFmBbF10PX9/1YXPNj3JOt8qmZU2w0VMCjiy75MjBWyrk9BZDo
cTj1G7+TJCJtdt6BMYUjW6ZExyiHf2O0HMQN10b0BpgHg6w/0YhderpmiVm3Vac13+2syXvJv9uJ
VREzaS9LekXbWnG2xzkpyVqvQKJfOg7i/JWSzY/7GjX8c9Ry4uSysl8XtXNVAq5YeG/JJEryu2Eq
anxLykYxBvxzzrOHKTn+w1UqdzoH4CmiUu5oH522PavdhB4OH4T9COKPXWNHUeUDtGTsfsOA5iQf
FDvgRdSX1lR6qqzKi5YzZXTWD9VqxhY26lBUFzyC58zF2wBVaoYzITCsa0yAECIJ7IeA0Uvx0d7J
xkgxgUXVKD9VbiNDacwvc4g4MbK0SLNRz7nfuitWiS3IhKIBcEJphNi+HbdzTG9g/OFE+nx4gDEG
1BgOO1tH6VghrXads6gTdnHKseIMsDUbmog0Crf2XabdK5NAHyd0r/VI2y+A+hqRJcMJ6YmNkJLy
y7U9OToqr4NkhuxsR8kqFLGJHJuQr+6q3ULXE67oqoRRfulqToXHlLCluswa5O7c28smiwZcDEP3
uFoHOhpb313oiK2G4RkzjKqiZ58q7GOSiYqr8m/vUaUoYP6rEouKO+Rn2QSeLjyBTKqwJB182XDj
gvGvm9wQWtSTb7q0nP39pkJZpNyI9dyIRFfPP+ZlJzBIfSXoWiWyKSd2Ir5KNkUc6ftXQx58z3a9
ML4Ue42apt0QH7ZM4bxsCpBvkicvlrt9tSUdUi5d2IlvRgXZCwYYWxqkGlkFz9JL5L0yG0VnW2FH
wBK56eWGcPptDX9ITtPqb4BuFQp2laWtHwtXU71Cmmuirx+QXNsmx6cnXvh610piDfiwD1vyI7a8
GCnfpS4c9TWFhNytnXjQrDbveJLIjZUOrANaj+ItyoNGzFu/6tUbHDHNQOQ68dos2KXYJIvMd84V
D6xHS1AYghukPFNhyw9IyGKfuQCXKDTnSc/FJBbpgC2IphY0OLezqmqzatEnG+8CvPl4PpAFRpwi
ohmdXSfXbvvqKqZpzOqm/l2LgviV9GkITo/l7S215ZCmlFJMDlw2Ce9pZgv8sEQp2bjRpLI8vrzP
OevbNrjgzkP9irA+BKKiaxZKpunn+iH6+1fZaLpplcLAC0RVDQxonekK+d3RrdkhfjLAiyu6WNUg
QOwcdp5J0aZPpgJEV+d8qhwYgF9WhMesa3P8uvb5Dkx8dYA22rFZRjcyXkfbhE4XJmiUfQOCG77N
Rl/g7nW+SuPSlNyC+jzlEJF8pY/MbsaKTgBRCAAhFPbanAC5YfE9xtQA7eTlyrIaemTYMMOxOO+9
GY3RPzwKCEGqxrPUiTysmh3VO2DE+O1o4sI9o78wPOWHzhy2VipfImJ63geZOtaDxipk1+6Po81o
zscONH4Tv6Oc08p9iBAfncTH0/0hyAU3jKzN1JP1eN1kmDmUuV7SqWU+4OwMGlYqUQdAhrLiHUI/
VkEeIt9V0gVKIyHvpyTqX9idPZJPRdriAq0u9HiF2h5YC84C4uHNEnC3Xjd8j10jm6DlN00Md3Vm
LRrW43MnkRbLqvZWlVqY/7p3LHxFvQHIkwak4GLvFX30XzN+HefScobZO8ofxyupuUdM6Au7r7nQ
+oZZAPyH7nvPpEF8b5J8mt4ec9exp178ji281VWMYugZk/33q2h2tGeGK8bTafa4qJKbMpcQE91O
ECUtT5zLX8uTV0YdETLLtYzfFv07UAvUR3GKDdzp/8wpQMFQTNhmVIib8yEG3lumOOTGyO7HlXmm
vFGkkzidMfJWnMbMolzOSGiSijz0WO6LI2rNaRdtApGNghuwvM29OVylGEVnxJwxKztXye3f3bR8
QkjMhXdXldnShIf2sOGVCofx1vzuNMBXWaDoAfYt+B7pjHhiMyHTNvqEMw8wINBsBw4cngEe90qc
YIrq/t2OcWl2T8mBE8rr1zeJOuOAPHCSIN4iVpLflm6E9JncTeoHeV0sbWb7B98FaFd0FHTdFFhX
RCnrMqBnCwnLJ5UuHSk78mthMe5k5XPCV/2zmIvic4ohNirxh+FSmMHKBVZ7DbymINGNXhszPtU4
PEPz0uWX3WGxbjTqf+A1Wif0ofxw8THcfZ+T0Wlgz/tjCTn30e2h7PxS3ox6psbKtm1LUWTvoK6S
JF1K3nM7UFeXAhyymCvuDk0EWJW4RwwOvJEAmlKgM/NqltqDpwRBAf1tdqq763tKjZUedJaVO0Ze
2ZVzbKiUhvBH6rwTyEWOx+wDxS4mFYOOhMGuvNE4L850uENNm3YuLT9nWR/QFrLxWG4aCgptdUQA
SZiHXcj0pI2NWaZqATmEgniI5CghKF4nFmT8z/P4/vyY2An2KXzX8/VZseod5wJ9eOC5r9beYdkG
v/dLbYl1mJXEUssEF/9jmxZNtdWbhxgztUuyG+OWCPB/9Fpo+ozS6/4GketN3KE9XhYBTL0/Ql//
0BC/KwlwXTyO+eETFDG+gnD5+gL7SkYL9U1B3+3FjV8lgz0T/5GrM/TbjFemUeHcA5HmXsqGXLGq
wDVm51BiZwiwNRoTSvhQmrea7xX40Dyw8JaMZ2op5ja9Ccb9W1qrGnp7HlbkRuuTHCakh10FJOR7
KshoZl3+JfvwpcCSCPwhuu1G4lk8GTGdd0Es3iUggHnM5ogjPn5PnzEI79Zfc0q9zKPubfq6aNIW
AG0xzkh35rI7a604HkUcwHKlcD3grf/qM5IK7h5XSjl+7TpqZIOdHqCG4emN1vm3Bak3Qkc1ctf3
fbRhGfkk2kkRczN7kF9OyV/mFTlAyBpnxsGhp30yjAMLJFtkEaIzlu8Wja1rNwFci1C07Jo1ngnd
SseaTmPc/CxYhTbSXdAclDGYTSCYTv7m5PfDJz/U5NJIghDhiCtRchGvApik8TOzaRLR4eK2wwa4
qKOAUtqQoYDkF7q5MUqgFdonSUB+nmdS8z/TSNOopmF5lMJMTZtYgdU3S7EGUPkSggjLfX+itOml
dnmCHT81vr7lax53tLG62E+qddR/9KR7o8Mf7BOSV+kTNP+sRwnHmoekVpyXW5oj5OaYQmdvx9EL
/0GuPWyTJOBGNo6rJnsPYopV/2fom7yU53l9F7L/zGCZPeTYbVdCtYtutJqDwDkIS8/dR/j9RobY
0whwBsgnptgDvp7q5s4cn+jNLREVLVLfRE2rVUS/aj8aFl1/1cwN6faE0ygj+pQTpBQdghSn7Ryo
ecw9KF2B35mOwCbWxZXf2cCYlNS9Og9iVZ0Z72I5nZSRFnCIDH0oNejaiuTiWj+0d470R8FXQcWk
P44y4eN0w2UfQDXD6ECr/Yu936UxiCmvEK8bP5THg1PMSDFGesxqK9Y92hQqDAtztywSJdAoPe/p
Z7C54tiSKUAyXhuUvtvBRTKabTyu5gqDdkknejbrS2GGIK4NLagdpZ19otvBtYSRFSLJrSbg07lN
yWH5cC0Orfy6XPTlGB2yDcqu+SnUk389n/acl7hW111dM0oKGZ1eICsMVYGOKGK8HWV7cdY6705H
0LBhEpqyBBh21L/zt2EPxAm7HYjWVj0tZfLQnaeHeNODRZaCMSp0EulWGLm9VyhVBt4LhKmlb1J8
tTcpkN6/RnFvg8QfYuVHo2757Uva8W3pDCXVaFenzJKhO7PyEpcaVukpI4i9bcdPPaULBo6BTddv
GuMQFujqLJySnIW/KZLAaTmM5ufhpDjUCyrT2Mybjc/xQOtteIXaeKFaDt7j6C/vE8p39KLd1Fag
yszDosx2l4wRzx2e35X1wJnBXfhyygn8pdKryCO5H0zgK5TvXFH1vS6GFmFdVsT22Wfmp+fDXSV5
5IE0xHIaveJWbqTGTYaqhvn+LdC9aIxxza8R1eJ5Rj2frIW5haC/Pfah5Otnny0210WpJnMHOAYP
jwuLfSvU9bIby13/0lri3YIL/xbGjlscDZkl3tG7Z0gixZhhWu4Fx0TRKXvK3pnrAwsQ/uUO99uZ
ypGxz2ruYXboIV625+dlPhU1eB8NijuWwWSskegO7rix+QIflI//PVI3j3Fj659cMkv1nS3Mgm31
6MYn+TgaBRy7axybs6mrIKo4i9if9ma0l43i5cc9f2xYM5mUxuW79kpfY8v4+stHDGFUctJEpKku
oN2c2npNR+9orhugjjrn/jFyOg/W7yxxjPaKqPXIH+3l73CqmUhABiHMSfFS2kND4JCDHNubwkdv
wb8bToIBn32XrKfC6UaT+TAjh9KqqXhTtYL0HEKNx69Bw0fQ1LkqztsmH6nwmdC7wGBGuQcxZbvS
dDZQiQQYnNa4Yrclr4mT56EiRedaLvQFt++h3YczbUwbRlVwQO2wuSFS4V+9mg0Gzp6kfHaAWsqf
hljIrTqEOMqSq8tN175545V7eQQjYoIQZd9lALxSQkiwVNDiU7xCix+A3HN+eySNBZjeXExW+Zug
8gKHfVHXuH7sJyRC2OhPYrRSp9oWqIPB0EIeFONztFOW8sMx4NTzDOET43BMNC0caUbRfVG65ssA
akT3bBGvYpgltUQQf0eB/SB45sHGRRNXH69T6btopjxyMTfHqvSwgp5FCFnLk06H0O+D3/UYedb5
RKBJWty6BDLvkU3X9NGlf+usJ0fFzNdPoO/+xbyJMgQVatAl32WdILeUypXBp7SmawTe4akqmk+3
wA6eU3SoLlbQbBYDk3m3//adewJv/Q52j1zxE6dOwx+qkWl7FkyQquqpA1vrVSmNl21wE+CHhHSn
uwZbBa2LB+7/EIc0ln25LjZFWnQjGno8qQn5+gQssn5aY/BKOzT/xQy7vrfF+7Nu2wbKbTqxnH16
JGL/06+6flwC5qtLWgdjyl1zubj6NR2oZZSBbAz8lGUx+Vpd+lFhOW4wa7aNeP05Rv5DyPvX4hBD
AePXZMgc8y1ifI7jVYFPfXbsgbU7/1Vb0H3gwGOkodeMrLWnhyBJjYJqSMY5uUMggIW+WxMBvMz9
Luc1vuix3XU+5dMIEKD6E5Ri71Ea1O045xq5p4gO26sYmRWDdCOKlnElr0h/pa+ITM/RrGQSB3Pi
blvl9TPq70FlwYfDHzH8ghywAvlpjrirv9LOvZkRIB7/HBzx9ZXN51qswptKjqGalKljwaG7a/S5
KZAshCvqrRGX9g+w8E3Q/fXt6Rkev1TNAdiCT8RRTI/bBoptmxlhTEXh7VsdRdO8AOFhaGW08Hsd
eZqmRT7BYFd8geFUxN0wEzm3jNbDhzKgq4vKUJv1FMk7O1LkqGwpEzuMZu7mMxd4qtzlDXGqqOR3
vDy95HEMmMGxadncCHK6ksKcRDAf+B2BB0UibuxYZachcWqedSjb15FoVa84jvvaYyi0uoVYDHtG
k3uDvRBKgZyEG5z2b6v6iH1ouOSz1dbZP1geU+AaUSP1sHhlKLZ/PiOMSp2kACiY/Xg8VgZYtOad
E3kcY8nZRj4plCuCyfM0GqC1qdAp1xdVeiWvR6HQDX6xKE/LH1EABFFayTQGH94GXwWjVLhiNEZ9
LXTYvgKM0lyEOV57cZ6eHbLpgjXRL2sUwyNcFlpsJ/mtD2ff/Tuwc8I6w79Rfels7gLxQLwbJchO
SoHfOsZncSYRQ196PKyt6McBB3j/K/uYWVbF5oUKWzltk+A6499VIhNBhYjcomS7hd2L3py/LYZj
xTtOzqQsTpabTufxqasvhIvupiRaG0vEq7P5i2MjU2rCftwm/lqx9QarB806SDOPjZ1reLwEy2qz
rbPvBpMGJgLOXiqMDFgrOGz401OFSq4Zam7rv1tfBMKqTLygaggoJWFE5dHmmYU2SLbdLkz1WuMT
TZkTFC6YraMKqTmVOazimSH0hjdZ2e4H4wGxnLcGuoOutrxL9WJ1dzr/hX3jKU0njCizmwnPCczK
vBc45AsnMXKiVlwfIJMME66QgingiTXL5QchnJwZmN1EGkyGdeKj6QM0dDaKoKByFmopkYDTjr0E
IYD900TFrMzxJSf1cR/P2XqueV2vPCOsQz7SMOV7MMP1ttENWd/IBW3eu08e5rCP9aeoglEcqZd5
OdCYZ4LngxOt1WcJXWWhCCisdOPiIJ3cVv9vbdDsdXM4pDncxB4SV1scG8NBgOM3wmz8Wazgr34h
PJn49Rm6qjty3k7vFlCFiWUSCrVCvdigo8BWV3zr0QkE/bz7Lg3JrDa9zmnHlolhhaU37AFro///
eq2jShmqgbx9KgDdtC/j2oz1kHkMWbCgoyPjO4YA3uVD1NBquiYk0DmFg87XunIlaKRthRDwprKO
Wv9U5AD3w5wez2Zfj08u+hkHapGEaTxeL8OXn1Y/2FSQsKMnP72NKANZDyRyMuQBWdBNItNiKUy1
IEs9+n8t5pebuwjlVYlzQwBYgGC8q1MOvocFpbgTSbxss2MmJ2+byxPVZHq+O6N6Qi0DtE56qA8x
OfJihp42lY4ceG8Fv0V1EbiUkuI+58Hd4rW+KD2+HFpTGgg8/oXMANUtQvJ4IlWJaff/D61m7AaR
1gmmKVy2APBwvEgIWeJy7kMxQPZYQ9ZAcYRfWbj1K7ZbL+D2p8Wntc8ZmWhXaCvG3t03X29zmHY2
UfzROVlITOolaPdwxoQPVoeAL5ZbboGNBj7Vd+yYZy0BZZB8/Geo7qEbykW/c6HKD43SBXkSqo6S
Q1Sbd/PA0o+J/UYkUxTh/6S7S/Hqhwk5kTgborrR03/Ri8Md3fuLPw/gGlj2YzYGwoTfONQ/BUGa
v09uVZ/rei0nsxCwJyfHob1yKDj8hjAsWtS/enqccFKKa4ibcODaicFb8WCZZQIKcQPWgKbvVJTO
jIaIaN4HERDlpTUUelqJ8Gdj7X6L1ydlK+mcPkdCCNbkqDuU3m2UBgJm95N5QFIxEtXSxUGhoRU8
2z6YjjQ8lnGMP2CWlaCHO4bLFqSveQjSRpajbDQhh3SYXoYfCyzJo6zxjAN6eSxy212EnYOs8J1P
qqpCNsdAFGRBSphmzJZsdyURRf3V0L88PILW9wqnkJGppsVzinIQS0C7d+MnG2JFlEIz0dEGEwGy
VDTvzhod6UNOdlj+Zqo5gigiI0OnXmNimnMoBfoicaC+VyKq52IJWMXw9B4mr7rtNNIDKT4QCbTN
1BvO30vXj4Xxa1j1JEdOAOIrDN8d4wUYN+pNwZ2nqAsKkTP/xkj0yUzXH5C3oNfF0ZIVizkRDRic
b9fxq/eAcw5y1QWVxMwGiWqUVkxz3RNgEXvKyRR6fsZx1g3LrOjaW/3Kc63hSyCcloPB3KX8W822
dP1XVI7bzUDkJe5egQkYyGlTPBj3VkKMYzzJJXEeR1dkkZtQag5zQlYBTUiWt9/H2y32h2YPdhm6
xLfmVPOEqP3dEeIc/xmbkSIC+5ryINIJu7xSGLgF51mqRtke765c23SCueIGjaPAg9Pum6ZStT+0
ILbiqqJWXBm1aJKnvq/+wL0l0un1PQY4keVAG2QQZklawqm3Vnq79/5Oj8QLGzoohVYXXI6ulxCR
8bKja1muaJTGxmofXMZR3Xu3YOW7LC+OxXmF740RXJXuqNj+d7/CLvI0Kxat5vN8FEeVjnHNWcy+
Zt4Bd1ICySSx2sgsbl0ttCA3Q9xnpqUmPy7Il+ybiJ7sznDyRSus6CSe9VdBISJk/f6agh31meU+
MjSmhmeRuaeWDKeEGkiM6pcqmuQPLKOc5zzv1n2Zu2QxEZYaPJMF+davdoMJcBF4LT1eBYiWxNDw
Ccd5t16g7ay73m0cPC9x2lLsP96/xtSO+Xd66vsZ15+gBKCDFwLz02RN8GG0CRvI+sBhPg6rKQad
Qo5WUgjEDL6z3keDAt41Psq0IbQ+raUiTUMCm2WpHl93H67KPSGhHQAfTaCBwCCFxY5z5Ho+FXiE
z6oO8Ixw1Wni1y7SZItFapCU29GdXisg9PDUW/XL7INJGFnPbjrzj02UJt8cY3mCnttyig2HDIh7
isaBPjASvHIL1SjnN8Bos6aRrhj+wCIwQvdsud0qbCqnaeYTnmpEj8ubxLLjgTbifYGFfbR+C0+x
08tCmReEXrXHFVzl+4zRxKmGcf8z6zisrNokLVlAnHFe0T6S8HuNtRAYsawc2KS8Q+fVX1evq1g8
lXP5nvaBa7NOVnCkkITfWnmq1pRY5KSh14TOX+z9jej0fejnrotbOwyKlo5UWWBcjOMROubS3+U1
kqtd/M5/Mw22nqkHPlTOOtDd1+bxz3qQ7H8qzkXUrAnuNsxgbZ1BdtCCPU7ejpJgCCPAbZWzGioj
pb7EfLczH18T82nWzyNdp4Loig7LkE3XVHYQ7+gieW5CV7hQXJy/q5uQUMGg20ZVERDYtHwlfUCJ
4B6dLgYv7kGQbefiS/QvthFRigxi7R33q4S6hkYnIW/uR9teXSNhKBsDpcLAliHSixy/HXJOXLKM
9cpHZEjHGrRuGTGM42UM7eHQN4ttEjviDi+47kTgQSwgi2iUhcs3Oq23oJk+w7xjH39vbTsWZKHJ
NDo8odpp/bleNeXmHdTxJvW5NR2WzaHAI51w/nM5hn1fHTnoLk73f1yJjFwCCWst9ThjpCZ4iJmW
id5adCQpTvGeIoL8IdRL+bK87JTtCRatS/9J95LCTQ1xekNgLlWSCN2q40KjXbC2pvUWBJHQqycz
3YmcxcC5t538sEZDPlwwlDpnh84mqf857+5rFywuDvli38KyQo7kJUyGKoYXZ1nePkhgCwnjDvk5
p8ubmhSzUV8EdlyxtMu9WZInCPPtBMDQzgYkkkqrYM58FwGEg/TfTkNqj07+rcDnBC5QeYxpbjOo
6OPoRBJVfoO09T53WBwB9hQTpwH6Gpv/5+T3Ov2jzNxt+QK3IqSFPp8Fvzd2CiN1x6nsXeILLgmO
XvF7JKN5P8+xk3geR6oMwawu/Y+dQGJUJu6QqonZkZAlckg5oM7Tg24sYaOX5uktn9426wXxP/J2
ZqUerPHCh7L4B7jAEGdyrgezmiT7uZ8UKZhpekHNl5mVdlhxR9ieTN2TF8hdCWFPlkL/aMPg9TG4
2PuxpLbvHw6Z2v6WckLsPWHLE8qYtOgB4zZSJ6Om5ocfG7SZ+BJDj/dL0H0Xssn5n/ztfXM2TqXg
toFQIWAt37VqhVVSoRoXtkVCxRyTLvbxD7aWj7YqfRlwbj+wJ+2QUiRyOnVI4axraa35z6L5BN1j
497E2Uz/lgVfTYTyomfoYFJooP2Zn5LjBi5IhdDe9pqu2nGkYDD7VTxy5tCbaFgUm/AQ9wfZ2VLp
tJenaT9GLKohJIYVzRm+A1VOek8Nr1aGdiNGX23hlLImKq4t15K0d9uFzFR8mdl69ouT2nRNu5d+
gftMnc5jIkcUHDRoQFfvKuMzmlt8IQw6BCdrvpOYNry1SPKLj4IS37IEV5VVhTVMKHFhf0ihwVmM
+wjKZvzpjX9Y6CfSYUtdsbDgVghrZc4v0sp8Z1jo9eZHx0bFALoN5mA4EOdF/b880JGE2S1AcF+m
4HgETaBJF9LKvjK4jayPwyxKWRR3oibbVe9BZPg4XIh0l0/61eF12vgDCp77gsVlXM4syJNvkWtz
pm6lmy9fPDSQeD2Uwx3wkDxtiJrQx5k8ap5gviwuM1AwsTdTqK4ELq0svOGUI3ng8CY/O7z1I/q3
SERIMN1OQ8kJxnpNQAWb2Bj0QUi5Omw1yHiamN1A8lHJd0DDwQ2p7CiDNpqpzZzjN2tD6qRBtnhE
tml4TG1CFv9dshi5XskKQltNC5EzgDDxm1QAAY/fgi5AwqtQaZlvNA+7BHcr7V9fdT3xLOtS1IvP
YZD4WZHX8yWCR+Wjj3YiPj4Dw2lIAOT0KNBbs1CjBOcPOHjniVS4Qkqw4beky7rOtzlHWeIWk1ya
duxv6HTm1CvfSVXsifGUS0LlixJu1hjw9wj+2OJ95s9vCTGA7rc0k6MVc/IY0ecGi6IwikghqtZJ
vH2IMElVIj5lkuhcHhESZTbWFnFR0Mj9S3TUUaFsxELmxRC1pZmriorbg7rOFDvaZlR8+k3JmYeS
lvTgA68FF2qDxADqihWbOgp/1MxMYWP2AtAxqQw2eujLB6EoGKWdyufnwQqRdoT9ESc54XGgkX4W
wD8g9Me5LcPFMdYMYmXI0F3tJEIebsxmebrL1+BWw64FzkM6V9roZ8J04kuqeBV/eCkxj71FNnKS
4VR2oWYvnujwF9JMzGHVqDIoNXpgzfdOMD9BPKB7IVHgyK+YQ6eJDV7aH4ziBqbSijGmcV0NQbbH
Jc51PXSWqan47Iqh87xbSyPAuNv0ykf7bD+FwJz4ESHziI58peb/q7cxBO1TQTSRwDsmZzcqw/vH
W9PDZz1z9QOqqSsTvyQYmlMBhOhojIiH7hKyoRfYsqeNxoVggRFikYc384RZqqH4YkdULKrLoPgY
uiaAN5fLe+J1czP1j4RG+r+R4NZWPW1J2l6q9t2IHv7xg5Bh7yc5ri6owg/mxGsDYrLT9jMV6k1O
DpQ76VezfbrYws4DpyEbaSACMAC6tyIMjEmenRyDOQNffeEh5GuEKVNFT/GmEfAs95/xTxXigqwd
fLtg0EVD+pBsPWfKx86WYg5DSiX+iwoSTgr9j/VGLW9vQw72Op0FaV5rnwfPLH0YZeaHNm9fsg45
KD8RdOesyWomYsgsO7ZRCqxo8/cKJwHCVs3KgwQHG/wM+ESI4bhD/mpoBNx/3jsF5lHA+p2pKGZh
8oFZ+nx8zXDH5EQUpl16NCjhb6huZJZFLU2IDyFT5h7+w9VOW407DbhrnpS8YhIsJsBFHsATA3q3
sQ3Nh4nf2JrAd2pbN6IOr5SO8dx6Zok827rJGNMtd1PqVK+OBfdeT33hvyT2AH+Pkae0bgRb+cxy
w0Ix9RqJVAHXe73CJsTHkWJt4IHOsyvr+u9At61/hdpsLFhizTsYZ1x/I77CfqnUaZQCStZ3KC1b
j8AvAybI0KsJ4EJs+kUd0uWUqAO9tCy0JC1xUFo8O4aecAE1ZBIPNKiLmVpi9ln5lFdQPBBlQi4B
CSoVlRNXmoxJRVqMWf+b4DBQ4ecnwuMtsJOJaKJABupjgXBmpEWkSpWQzK7jtrxEoTERxZ180JzX
7/gSS6bjq8iJwSWuxXZ4vSg+6a7W9WarovqY1iu+fDAS8M93vR0jW56ZqzbTJK+Os+sXevP4i5TR
wokRXcgYjy9BGC4GpDT0mkzmYtlFjcQjKm8UGriZlnd1S3zr4lihA+VtX7bNkEsASl6HNksfBSdO
x+NYPxi3Pz+lNzbeXbZzqpiQ6M75LtnVDcqNlkwgl+T6SIkhTSpdzLPJCPV2vXJ/G27WUSlPcPPA
Qefr2NpAycp8eTNy8wAPEdLqD9Fmk3JkaVG4P876Z3tQGpDsVjpXY2a9gqECyvG8/yxm2mAmo8F0
ta+AYN3ZmjaWMPenQ7Y0WyejoxtzN5WbpjfBJxkdqnQqlXvavn7itsxYTx6mvC/IqPOL0AAbya+e
6aoavOxOHFNOxs2sovAK85UJiEYY3y7q7+K7BDzbI4KRIZNkCpESmHT5Rg9n94vucILFH3b8vUAk
pTWFt3miWBbS6FHXDARGH21QRwSFYQLYnNI5N8Jzu3X8W3HLZkNoBwB5L+ldjG26EitveJYmn3p3
l8Oe+fzTCR6jFr/PDoPnj0K84N/9MK9sNWOq7w00Zj4DyzpDlCHZsLIRh9FKGUBrdAE+5DrenVYV
um0xV4k4GX5Zf9+Wx6nGVLmL3t8eIxdolcKLu7WuHOx54FPjO9OPcmCIphQR0/1p/Q3F4eoxuYVv
VSBIS3UDF9rhY5eNy50NNZUXqdBAt9B7v/kY/beDnHvHZ0Tp7cOkgQ78AshXoHhi4ZYM150t7QGS
0Y1cExj8TSxj8uz4ZZOoik3WAdAara5w82Z8/GgXJhqHrxdOHzwTLfuQdFGIUigsfjBnosP/IpuZ
ohOLtGTcAHMlNQZh/T96lbtX3fwa6jR90dC6S732q0udVTB4JZywGo36MaP5ml+yfqrlHaXGaANo
t1NIOC4p7VjqCV2QR04Kq8VWD7hD9fABjVDxVqsePnQRPRv4m12/i1p90ZxNdJ4Byp9onSrJwiqx
YdC6CcqnAPcNrFiEAGoIGUMIC3EDIxfplO0ZMprWKaAXXtGlfc7omhuNGXulbp2Z1SpFKzUIMbik
JvLjv2xMY0txRRmh5UHoatKm3bQz8Tb3DYrFm0FRCn+qpfiD+kw8MwAYnmCisXssGoCaBDgLZXGS
k9rVrgk8u3jmd0xL1OeUuSsLL71icx+pOdZ+CFVTFmnADptk+MZWdeeJROb+521++17vxiQO6xKK
4jaj2cCypgaERgjDbi3dasXBFZ6LWKNqqtpS8O86pbHK8g8TShNdtGMw+ZVS0hQfcJmtrOXplz3a
qg/uj6SO15wEnjSmvHG7ZUV0hVnzjz5/pBt21QHq9t4WkfVYfLW8XEYejaZMyFH66YD5glSkgoBp
u97lVnXsIiurvvS7UAKsYqzVmbRwAJxU7eMbQ6V/xwEcAdP3iWjJFzEyqBEwQs/7RwdcxPmQSe82
62RMoyG5Qk62r02sq2QYya1adZf755uLKmiFlu5YLlZh+hb/6YzjBSf1ps3Hvv8LKulzKYf+/jbc
5xLyo4In59b5tli0UWZgTJfYhIZOTmZprcoTYm9IcCCAZP8UH6p3OnwnwDnXiuhPSlSpi41Gvtxm
YRUTbj5NP1S3KNKO40av9C18HxWww8fcaYATb9cdTZSiJpNDc8mvxyVFw3H3/cC0knOcunHpIbuN
hk78SLuIfiMCd0BZhNQmoaUbgTxVuwRhLjlGQphXDqSPRKxpU12tFWsV3M4KPmaweerGfn8jZeBU
ICl6kEkKEkhYUq+Y9IkF/jonVuXLdS+KprFeLnvdKlSc6SbWrQx6cjBk/QSSwrw8Oxwda6TGv/Bd
vIuc3oceoZPsKEOA7OqP0/655Onbhsxlq1ZyRWfi6RmyaOPFeOzdpx3XfuGN32eYvHqNvuNWoJan
ToenXqLXGTXvTxoKVgUicdmioZkxysp4cIvj92fXOhKjPcGD7x5lEUwDK9ZTWDpFetwG8TiNFANL
pPf+sO57v71rVm7Ak0LKkuHPRFq4at1LFzWNcsAi2Vo+Im7RfOMeXSLJlZppJk3mATIGjuLVjg4z
qbA8s1AK82fgWtftE9gFpIvGnFhmjew00xJRqopTW5r/cDcKjYlKRMdCA5bwjw2t4qya2kisH1/s
N04SqhXX28WvmETX5ya0tcGW9fIiaPnAoYsLxPSVdI2n6p6tIIBfudKdXqV7Ch1zQ/ia+0xE/iAA
YCQ7bhhvvl5VV7W5UI03n8pQbedkyfo4JT/QPWYvh/ICjk0svAJUOXK9L/aAhztPy1PERLFKeM6e
JZxq0FgZ3s2SwISXnVGWjjCUW3VWZU7e4noKxrBVg9ZhQFipQ/WRld7sEa1wexP6PVA5DNhVBJsC
nR43sMrigWtAi+Gokt4OrRnQ7B2pliybB/z2DTX/swP4n/BtWK4lSOXj70ym8jGNQlaXeCPW6pbd
5PN9KiqS9RFutwQLqPr9BCtgSavwTyX6dJrRqazyEyipO4rkEOY6/B/TfipBKwv6DJCZGB31Md6K
XsKTFbojWJh/oKS4a6ssdo0FqFVhkw+tT07nHnuXWyiy86i3vIMtBz0vlYzDgmPcpm/QJLiMVmbU
eDo+r4CO42XtZEFmeQDZoBAffu63wRU6J47WOb9khAHA2Pbk+JEbiqFCZAPy/gbHe71Nm8Uwvxeq
qhU073IBPyREBVbcZLwQ9YDV0KjBS8XFfQ1eij6ONvNIwzALvcZoog9onu65K2pDFQK27uoBR5Ph
TMAhJZxy/bCZ40QU/ermMa26gr0WK0VAqiU49HmjvfH5pWYXJKt08C7BoLkgztl4FyNt5UCPnpqD
La5tBEQKRaBNcp76Ylxc26eiC20OubHCxq/r5vkJpiGAL3XyX0dP+A0QcgbhCEAQkWFI4XVoJ/4X
PWv3Ut2gSSCv/JqwoJzpBLP7PhlK56Trpu5n9+P9yIGRx/x+OfkBLPBBwaFwIbhEQ1hyU4cW1lEt
tJXKyvhVPWP7oPP5LiL6AJYEumQbKccxeyYLaiVo8pk4Fp4oUWUmIEM/slax2Q7YmOMNuRmfoAdV
He6yvQBIa7mqRxXGruXQCG1T+CPwVc2RC6TvaLkF2DHSKXSoQ3G4vMFrtPaju9+aJoOg4eTzJD22
AZzfDKoqzSzwxyaW6Sq62lfxIUpE/BDUQPQsOlNJuBraww/NK8x0z3/rydpaGb7BSrf4r31gx+TV
ljmk0XefKyA77qr3G5BcEf4Z+pNLF8QDjjjox2OJpSkv4EbnY1Dx8edvn5M+SicqtVCnyVH+RDTy
3w73yLqD9QVvSoTZ7c4ghfs0liNTXalTEAP+9LFjnl/ZFsNXq7rS7Pm5PWz7Oo4cqRWbd5Y7N1Gh
XxqmZDWfuqJQIN6umiqorspTxgI1Q8RBrtPrzd0EbQUxrgBwIs4wuVDObgWnGeJNj3gtEa0hWw+d
GC2lIQWGApNimQbtSg3BT0OqrOh7U5+yaQGuGBc/TiCQskbqDlM6BD5zgxrf/gv/asGGSescCdl7
qIggzTFcRqv0NWWbb5Bj9Wlx4h2NF4cZ3NHt0k16p7Ny7R8kYSf11lAJIpBw8aAO0PB/kVSIrH8S
69W0RlrXVYVUlal8+we8NuNGGSQS2BwXNgDy72Dfhr5EDQF3vPWavt2idUFMWFKqBGZ+gFUNm2fV
s8dQS7E05kzqDTTLOeZfpz7Ntx4FbhvU1fXQ+W/MEaIi8eSzGs9uM87kKOHoPCEWtUYkv7i24bTu
zd/2aPr0E0AGjwZBk3aW7K6Kbm5DeOcLwpKppfZ1nz4kBaIw4MOVm/WL79p1SfMeU6mJE60ifAV9
8+nkmJlLhXV1H3jGWkyZ86rAg92j1CXPLsCyNw6xIdCMcUmYSdh11fiEB2pEXZeG00l7qknfcHCh
hTqusDDoQP8d8ANkZmcWvmwFeFTSXhh59pkV7PlhAzn4Fnv5elG/RSGAWkE1+zX8RCQjQdXuZlh6
mjpm0gIp4wnvUCLVaICMZ4qZk6D2FQNfu8x9jJOuGH09lZrJWDCxYxKQOIGXJeftH7T1/CRbOX0X
WOXLkjK7m7e8FyG7AuoBjuqmcYE70GpbRay80yxoD/RkGBQQB+i9K+W/rdau2jwxEpqsdaWD46uT
MXWiIBXkPw8dDmZ7+S1VPAWsqjk44+oAQZGBYzHJlTA+7d3dZ0PFqpLghrg+ALTJTftkJ8A6t6Qw
ddfFKxDjy6ZKSBdhW+smy4HVP2/ng8IdfGTlVgr9jKbcUqwE+0GNawgRJxKbqvhYs6dbXgs6yLcD
i73wJIgpnpIzNMpVu1cXU4hQ8JoOQvd5ozdzSG540UcqFpelFkED5uSqyQqMzEl6s7MrcaHP63zG
BhpP7BAXyIsD/vRTC8hpZy04fkHv9jDOWcuQUW35ULAL2FN0eYmxAP8XbC1V8Y0bnT/4GzaGy5dn
cpUyFGXAZqxceBdq/VVZM/oVu55X71IPbs75+PNkm+uCPaGDp010liyjGHRDWE5BBx1MpN+V20WL
+fN3nTfuSpwct8h6KrKQPBpK3j6GQcNMyK3pbW0FeOg19B0KEeuRUX7pKn7nf8JLFwxPWUeQxbzJ
y7j+k+1NWoKtepPuKGVS93weLjwoIBDjozu6kcKSNfR1gtQBeFdsaIna0+eTJoto2MDEm7qcgHwu
Ql+FMR0tcPTgFeGM2la/RZ1/j5bZS3ikybZqcyRaoo8mfAiTtdi4nRa9/bTv4zSuIrpzDg2Ee/ru
5nKgoOFVZBe5nPU7xb+9U8ybadmm0ecRbh6v3j/OSD+F5JNNOwLVlrdZaiYDcYwM8IuwrshLkjmw
/L0OKUjcGg2Q9KjN+j9Z1op+vrztlMv8uQN/wZf9CipyY1ROe0mcxLe0eXpFCJiFDQSuMQnR+CMN
74reluBoswJjJpL9IDPAFges/cGnmFcXkU1S1NEkHm0AKZ9vMRt0coDu18wtnsZ10HYclyQb7ePw
NKMZYjsKMH9ALD/600+CPBs8utSeuGL9WBuf0Xd9vGsC4qU1Xcibmm4NhYn/v/LQoNrsSIUy7uU7
TtEK7JUWKlhkm/0f0aGjSTKID3Q6T8DqZZxPNn3AwC3dEdUttXkfI/9fJupqcuWuVG8qUnRpGOSH
q53Dp8+bvxFJQCgvHqurfcWaYOdNv2sW+KSa/Uj3/BCrvKFsYE0h2EPorM13NQvPD4wDNUls1k8d
Be33y+gUUAFN7+bOOUCZSqfIVBWonwUpCoBYuZNb6Zd13S2kFSLsM2M8kw/aXcDdFUzb8IS2cJ9J
FhGM1Nq5Dd844XMzu1GtOOGBpObRhPhVI/huXh4kzFbTElCL1crZ37gnIGnQJkcjx0DE1FABnv5d
BT083gmnL9de1bGC8u8dMmLDmcSFvVxFy9d24oei8qFwMirmVIBLtfoTRaHDJ8wHijDGSTtbH5IY
e05++ZE6qGQaWWrxOr9c6/jlZOAWlGnoIQvOpKEL4CFTlYalSPZVA5WNSWWRT5Fpyb59JNT3weK5
QkTJLmKV3yBQgF7b6QOA1HJTFQL+sPAdZES+G+IDIFcN89argApmRvdJzH69e4LnIQRUSbImGQX/
8UvtWOwlcmu9MsM9WtBBt18de/KvdrCDJLrnPaS0fChhKBcAoqrE8STKUMTY5HHZbLT29KO9++pY
HOKQ6mxWljKP1Xf38C8X+qichnOp/IFkO72X1RR1iUj27JThxd0zjN3vplzWAosJYsdv0pstMZkK
igsy2z5fQlxzKH4+SGv2YaoB0xuTRkQ+WTau+l0i1WzEnXw2G1UCyiRCLxISDqIMgatpmhY/n+dn
L7KC0fdxRIOJ2aLqcMoYhqRBgRGe6VT3ju6i0wbluLNUCnHgIRHMFMyZKAZEeZl5yjc1uM6kerft
rTaZwzbdAkIiRj1EqZ422zPcPb04e6Evwq9IZVOH8yOrHVljJ2UdYqI8bVGHwk5Dp/0bTx20huy7
u7b5wkdvbUc/Jnko27yA8NcfRPZ0OcAQznwq17yhLlxs+ERIhistDBdfIjbeqaiu50OfYtaZ+WZX
p8JRRQHfrwFWbF30vHYmIRjX4pVFxJsQdIOP47gPqDwW9EiogguY0FL/xQbfhSROoEqiErh1nb/O
d7qUB8BnbWIZvhl9iMkkjM1r9Iw/yKVcq2kq80W4x3jWI1+gbG6bAANCvsc9h21MEgRtouFRFLSA
FLLOyKwYO2G7P0QMzazT5+SyKESsQ0rNw1CB/E35j9otyHyEo6UyoX5Qon6DniVC7kiEJosRYqe1
AdMRnvyRPCBDma18wXFCgk6sKWvj08f7tiyYUcRVvdiMy+P80HusVMJrXlyl+MogoRPmfb0shunb
87Ds3Zx9hJP+sri7bJ654v/4vqXFsI4HQE+5UnzmDuiUt+IYjc1ocFaEFUIHIdDnjgvrtXj4czZY
UD8+FGMrTwqBNnGrgjEGYGtdYQjEW9ulM8BpqGCeT/57L9z0maJRQPdwyWIn1Aa61JI7CBSOvjqB
CXGBwjhuVs0S3J9CI3Z70/9lMl2w9veqk52TzhnyqoloVdqhKE26UtWGp3xAXwx9vt6yszxLEoDZ
UhrUqN95OXIQXjHwb0Wt651wt5SIUyfaGOGP89kxEh8WD8qoAsXD+yCsSz34dCQfpOJu5M0+WcCa
flpiZJlgsTW4gdNQyD8c+wBrSR5DzjXUqHiRKaVM86pMsC3HUATh1FujefFp377t48RsZ2DI9fnf
9HYFqsLKZeJToIFIB4y2cy3VflM090L/V2/VISNbm+OzgKfq22b6hOoQax5myzVw2ULjY/hXgOWp
VZDNOQ2jfiLW9jIsSn1G79SCz8caHa+faRzkUmCzUGpII8PZk49BSAVBsGvhuY/d3gJUKoSZE1Jp
v23zJfoF2jhNlUWEx+JRX8JSaT1nAmRz5KsL7tloBacFahKS0mlWYbjNffQy3/CgqvoJfs0H/pcv
xQPMRUkF0SvDSWSy+arNhc3FQelNdlzRue0NZ+fDzcRBXGlpM3H/1mNHb9PJQrcCn2BAxYcSo4f6
/zxPsTnyHIJPWV0cHI1fAjrBf0Wl7eRz/S34LzZ3OOpv0kLBAXFH21CNSv95eyqD4t2XBDK9Nzpr
1/SLuSsuevcyg8GxNj1facfwCszfo0pglop+agUyZ7el6CHbUUZsVHBrMPrZI+0DbWhOe92EKHBS
RCyZwtnyYRsroKSY8kHhU4OmIjNFlZ4wDUYAHzxQeoFbGBBpwOaxNt8gglwTJQCMcOpGZzwOOUIJ
ZA6MxErzjKE34BdvkJm8kPcSO2Ua5G1zb0ZYty+kyVx7VBowdDnX+Bg6Zrs/hyMQI3GEkhl/mr1/
R1qMMghovfRTf3nIpDHuRZVB7cm7VAnMwsEvZWvvy3lSVGnXOhXbkNK6QsZ/TXFviP6b4UYFRP7J
kIGT6TymS71WLaK/o9NQmdHvAvptVkO7ecNYd+LSrufdMHLyqVBw/nx9Cn6hD5/Y3Z4Js/UTCacU
jnn7WiYWCR3CFmYn4hrRSufJ0FGJSEfelvFHyYlExxuTbTHEK8uQ/oRp2JhTlXr0I72dckbzfx5T
igJ+KZ/S1xOWOqNtaMIPuNVimPurllu41T9rg76b8miD1DLiOQw5Z47D0ugndR5FLVdih8cdhQIn
WwQOQNPgZIS928KbS2+1Wl4n1gXbj3QokqUvxDwv/I9TQm1j2zcn5yryE1bQfc+bGAbVMANHuZLc
NWGqJIVOMsfx4k1KCg7MV/nCNDbuueHNuBAKO3nS1Hv+9DAFuaEJc7YY98psW/AMaHoKu2J0PE5J
zmiNZnb6C580Cm/Aosow4RT3bvKmPZKMH1kWfSoVOLDwUz01C31eoaGwjXy6zXeTW731r3a2sJTF
Eb7rnn86moRoYN/FEXQ/psL9y+D0xnR9/smdF014dBKd0A+egalG/ALnqeH+AI4EfyVUWRCbxjqw
mf2jIM4AJJpnwUrvk2BJGXxstfIn+6v4UsEEmPC5h6xo58cCAGnW3Az/UDNCnSd6bfa7m6iHs+8S
wOxvfu8lJ4tMny5pY21FrfpCpA5MoQaQfFgEMSiURYE7e6mvafXoHinJOQrQxn8vxQ24mqTnTg5V
Sn3ZmCMIbq/X6H0l0PXrAMQpzkIocK97Eoe3HPxQOxaR4EqMGGFUodisQTnXDPIDLAi2oGrBYNeI
4eXH6Lpox2jUX2QZwdnS0DEWGZrAJtEJSs9NDdPAeiGQxW+T9keMBAtcJ24Aj+PqkA0zRzCKQieu
xp+BExZsLpVnTedvuUb0ggj61C1hBH9Q9F0cTQ0e/9AXcK+y1nrCyx9oifT9XooqX77KsuBjY6Rs
/mIfDsHE3P3bYIcCOr8tTg4gQq8VjmIRfzsa+2vP7hSp7CawSh21dZyZJ3NTu86uR+Dh8nIHoqqg
yzydjnOF7Dcoq7OFoJxhoXJX4LyAfGg6oPo9n/wSH7g9vp0UfMa5SFv2/uLjDcRcA4G6iCqs07Yg
gZtLKoHYLjo8JC57fkik71j993kZe65YSCb606v8Jq5SG3PFs3oaeGvw1AOSD+WJoc1I61U1q4p2
vMdQeLD1G2DRgFuwvXduTbsZKLJmiUnbyOOTHaJ5/aAbq5cbeWRpPbHz6amEU3Frvbn8QkxRRMOl
LT7GWKl2nXXPlf7rnFK9+c/IJ0mW0ghHov8PnS9EZm1l3Jn5H3HBQ+48J+MG+a0BTlTcODtQQ0Z1
qfz+0d/oKyAJJ3+Q/7xBCiiFIL+DMua8i+T6XO7tvIyh95hpKefD9zvFbTzctBUL4PjdMbVkr6Uw
IF4vOb/1BBtI2qfeYqUMJIlnaCOrGE4XjtQnE2jfYRsbPD32JpENq9t3B9UHvio3v/idTlk1uClu
D7C2jKhyz3mZPtv4NKMyd71s6b4y6o2p5F8cpb/GZklyUf3Pwhmw5smPcfnDv3mPaGPtAWlUMHVh
L+902i8V4uCmWn1eekdG+OI5myAUorh7RMe9Iz38ifAgqNnwV6+bdXZquw4M+My9Cbtpna7gxs0o
N7m00/AtlClUpRCYN0wRCG/tLOAW0WmdZ0W88jyFv+U5IiIUiY93dU/JLf9uyBmIkv+LRXyWjP6Q
w9qS3kVDma+rgO5EBrMusqU7EzC43hL5pr4hDBMIosU1xVWplu5XAz18/j70SGjzagO4ewXctjuU
l2nPZUOaDi7RVgd/EtG5ib8xiCyPZYzH4F4SsEHqvzhfmnuN3ylD6b9DYFb5IHECOqDTr/i8gaiX
fZywQ3TZ4G++koClki54TxLdkM9F1qVj8zDn4Z9HRzHPvcVqyJFt1NdGF5WFWWgw4GoBsN2SCk+7
5nNGee8jdIBNeODljIKpG0v7lfEeO64OvqrpgJAP5vyqxdphh6lXrlrlVSx2qPVkpPSDbjh+og5p
3NPoLvXWJ92bOj2kfG309TkGnalLGoJkEbMTcuBP4emuwTvqs+sVUedGxltsgBsmLGQpc94fzwi4
RC/h+OQmo+AaaDKpox1NsrIesiWc/6n7NNovF/z5ZtOP1iVtUJvVnFyJ4vviy/VdjxjtTKlYwknw
1IGNkc/+pXb8HhwUN1654R+P78mldwGeYi4XY0AHuB3RWMZB+pwUFeThipgIBxKOnFKHTtBzLFjj
cluAi4bv/4d5+7RUHOdZdyRf1DfVZG/+mi/1/S8whsAnpIdL5cIv6G0w4rDM/IFRSviKU/pn30zB
I2yIVhc4yGtHY3L9BdHtyaUAU7XyoshHvLsN3WyoVLfLxM1Ft+Qx9kL2wZFXxJ7CboUrRFwCLauB
Sn7AVBbV113et8c8rfl9M46rD9BxjvLV6/boEjMiIbWBJo5279qxcYFjzEibGAMAHicvDfEPv6oi
a6x5QyOWfFC6mP8JA9fHdD7qfgeLKmDPqtn81iETShR+h0qNRJ9b6UFtj8dA7ykv20A4C2662DA2
5XX5fTgmd6vsyDlYDLnfgRYbpwzIHmp1+Oqea/MWB/tRCpwxP3IG9VQQTIAfl/ut/hMiysJI5eWp
6Jx3+P5JeckJ3olG8QDic4Yx6RoHr7ne93pqAqayCJdnUKx3H4anIRiX2IychbvQ1qdJ8LPfZey1
ErVGkK8xOyGsWKkQyloP2aYQIHcWTFIdtuLzZPikjxYSoXetl1wv5wmf4Go7cp6ceixRMQw88+C2
LDPsKdIegpCUak2HLtmarpMwVSSLDyOp/zT5y30WTtfx9NLqOnPQyuhEvTKGWs7yQF3yZXBxi1d3
619XWGLRMhNFqQsIRA5wuulDO0eETnXvqc8/4IUenkuG0p29VGw4IrahTezNDteKSzwzFQ+d7tcw
/U8gwLJfgh+VlN0YG9sFKDbzuPPkCOJPQSWgVDKtoM3FQtNUvcmoXs+KP2XCmG8fFUGPBRJnoWdd
8QHM3Q5wwRECxO39Zl9OhyIGtZj8qwL+ypImnc+V32F1i6xXhf8FEbASUYzwp/06N+GFspaM3cx3
rv9AsniTxnhEMnIx8Ggdj6e/0539o+cLnqLbjjedIf0sPMBUHumjnmSey1QZUbVfE02ZXGH9iwaw
zsNvwmEiTNOK64BZf8a4t4r82NWX9qPfPWrOXeBz2XMxqY4w9OOx39igjLmdtDEZSZ2EoNc9Lwim
qBDXhvTqZShWsYY1HviHXwgqf1+UgaqBh9+nzfagYYpVLU5mYrer2c95PevK8XIiRmcdMBb0SVk4
wopVtLTsxX7RnxJDlsIjdaU7oKj4kT2JZ79UkK5BGcIHS4iRaq3sbKKipftfV2XbessHgLhpaSpz
tUIp1yeAofBkjscqpM6jBTAGJ6jTRgC9dyyEeEfGLRM/fAxJJya5fcAXHWApeDwSqyGB0U+R7o7X
K/AyRckDZym3VepaMjsgX+k83cgqZi9rgK/ka8eP5nWdLa7k56Bytt9FUEabU1osMQ+ed4z9csOz
2ODXbsxbG6pI7KYJRKFXgDuQj2nvZKwGqMXiVOrer1bxUK5QNQX0ai/LPmgWgAPwO7swNgl6hK5a
qy8RwOKf29txYOwF3eN9GRSYbHARh/NUZsLNXytcQshjM8umnbKrAzhHvJ8Z6qh0B5rR0At5LupR
QRFvC/p13AivDpZbKGtfynO4rgbuvjDoPHcrAbW86vRoO2iBpNA1GnpXQKuz28k8xbsxqdSOZTMZ
VbWfQKCUIjMzXcHPtgSQtSntZSxRpDfhc/HYfvcy7Dmn0L5ZQjn4UI+TPzchO+0c6+8wlZrqMhQW
IDQ6pDFzlgXVu4NTiuG8mvDRCRffbvQWxp+DgvIFXQp4x4X4eqbdCr+AyXVxsPB+4GD9L8AzjZBO
tN9ypOJkbAMeUEesbjBoNbOKrxIRFTVReHTXLaRGyiCG7SEg5E8qJ4X0CiIXSNaGLUK6wbyw00Dc
pffLlSXlMXm3AmT4lAZPIto7orjxYReuMq6dSezIOL1OEZwnBcwLX+9d/+mIyGZwPmj9h8v6mrLn
IlLJUdv+iMZUPldxutFdqVEmemDuGq+pNwB6L6XASG7VYZdgcfuZJKpvqHogf979EsqTMhN2Xrwu
8/YvSvU02N9ShCG/LotNdV4qOZD5Onb5D32T/KxxkXqU7OWqdcHoDUAVFMKtj3lELzN/nw0a/AKI
57oGilwKH1r9i3udbeP912C8xfNe4Q6wpLvnFHlSwBH1JSKxrCGhxL3GSVleOR1yMd46j6akUq5N
E3JanZOyUT1t0OGWxAxw6NFtfTdf90p4m1Lpo5rSjFsbUcZPGOfzGBQ0xxeTo7HmYpCoxpaQzEOx
fw+zfVK42I/DVclTxvGUXB7fOg62NeiWDdJkq0RXwygEQuvFZCK82dxQiZhYX9lBJBbrpI2eMRZV
srjUeSYpWgiWNqIBHGsaEZec/Fl3uKVWnJS/Y/6IXp3wANl/SLzoq3Bg+QvyB9/9hRgO6jVBp1IL
G5dvh6MtA+qWgkH2LmYopBaQ9SoZHKA8kbRX+bYdXrFzjbDP06J9Bu58QtvlQ1DYcUVi1gG5WgKX
gozskg7E2msVXY6CYG8OOAY1KV4/dzgvEhsr1t63J7ahSvnePZ6OTilMD8Efhzx+/a0TKYZ1hmIS
K6oGpVaHEmbEi1DAO+e9VPkg79JRHxiACGS3LBKqVwlGGm9uil9MIuuQvSXQ6NqtJJmwQssz/FGw
W6AGj+BUn6HHhk94lIU5IWTpGzVYOKseOo3T0xXtgiOnvd9sF34gj9UULq88ekjg4PwcScSu8oyJ
ArYY0AHaMkE8VRkhR84KN9qSoQJjyscKpZX2cghjxClmfLX2s7YtHoHxcCir2ALO+djBYDiyK16e
T8wT5tAw/2U8t5f5P9cWP6QxYZDNDoStIAhvUzSYoYhXi9aDsua7xuKyoHMpm0RbmU0fRousuvuV
TG8GX6UiJyff5LD1B5w0+LtS8a6DAbI3SD44mlxTH+IrxGqdBztpeUHBK2JNflqICJMsqZAkyywK
DRAShL35BjzIOvPT8VZzZbWJ/gjV0QLnmB7EbGYw0kOz0EpAsNJr0/30N8EuR1RvM8myxWhepLfj
UKtHOsuUbCFX8V39DRhrdyWx0IEkG7oAoMY23JN4fE2iFBkActU2brlJG5p3hQbNxCoVISqjUiIL
ejqBcyyYEnDMovS5yUwyNWj2/CQrklyT+MLQESkDVk2eoaGMlJeaJ8i4l4PB2x+C2TIxkAFHPuYc
AYddSFMQcTWdekMaM3beGdlN0qcqzb1+DcGTQp8gMKBLXdGzjJQ1F6JzLw3j9gCqn3/gQcw87mpw
2gijvGNXAX316sqz37dOGrYy9cpdM/0OIDoP+Ry0IDlBgWH8coAQUnwDkjHYxXsk1kezHWstJgbA
amr+uF1/YgqZtCMYvDevEIzJaFaEWkoMB78tk0lb85GD/SmTgknjS0PRAEALER3Tkh4x7b+pubpn
kJVYt4fg1wibCPM3xj/kbbiCT+jb2I94+PoYUd9mwKM0hlMHeHrSMQ8FLv7PZWnqBAPnJS2zX2oV
vtvNPcJOUYYLi8knfiVVibxotFHgAdzg4sfDv7k4NlvyOjfUZpNyIZKnzCc8UXxsXOX7iMhX+RCV
TGAf29b+o2gVYCAXEUeJ+evEhET6HIdfTcLVoL71+Z3jYnwFwKONCTF7EcAGPoAEiucmbRvokQrd
hYzZb0pPenNoiWRbDYrw4w/J5UYglb2H6ABz6qQaQ90C9DCmUuCKyEkkxwQzOAhdt/X2TDkaSrEF
53VqfwpxYZQuPSgteUrO+bJKrgEAkSY9h2TwFRn6syMf6BNKet4uMuZDIz3me6Q0h4UBgu/PZMFT
DhETSvduAWRfQ3pwrFv90bYdonqPAZho76Suz+xUg2/C97ujscicB6Nu/UgtaD0vUTx1Gp/p9swq
ygKFfpvPG0gPajBrC8E/jeGc4xKWdjmJMo7eXSYq1RGpbmo3wu4U172l4kZNsvJm9TQJZXRdwkrj
2rvgYkT67ziZMi8YU5hBdCwzoCCuQUPTHM+tQBmLFiulOg5wGZVrKUGfq5Ci0q631VYLm0P7eTur
qX7VPmRNBgWU+QQWMHayl0thiqCJK9gM6AY0UFhTa8zPTyexLD9FxqRGDfEa+GOCw6wlKVQTnuGB
2kXMjPOHlDrkAG2r+vZlEiSL5IRLeaHefhqutbU+9yq/uXp7vgYJHCCqTKYq6YBhKBnzVJaQN6+c
5fdjVXnxqcyg/ePAnG/wNw4ptT2sPKlnZ+NYDOFMMVuuVwl2A/UC10F824eDed7iz/RBtM2GvPtR
BKm0PCHdxC9o4q7WKuyo44AcG+NNufy6718NG3tkxetrNDpyZ2afB6ZjluDEhS4FuE2pmee1Zgf6
aM/1X+qt28OYWeS/7QlJc+0YP5W2DJZZ6rfv3hiRKGB18QR1jCXe6SyJ8uIHsxUD0iHSe+l5B6wa
JdvYIuj/QdIYEpa5ouKCwuDIsxLo3kx6SmJM776YKDQsmO36WXF1ggYRJKWNDLb5oF99Q2BY0O2g
7Esm9SWPqzRXnLnmpiT2pGrj4jmaYlHliwr8FbZiA9w60Jbb+lpVPm2Boy0vJHRH+qPhBmFzUgwk
no/pnbPRw9FzhWqhiJOZ2x33+bQ34d/Ad4plg/qHHabTIvUg5yo6JHuVwsb04X6J1jVb6aS7mhEi
09qIyk36R0X7uAbpzIQD+TdyCEPFykjObEt2pzM5blFpF6jkMtlmWYu1GkSwXs3WqPT7GLTnnKpm
Xax4V4GQtGEcLwC269YiNMxUAEWjRQ4IG9pFql3v7li5ZjFrMB3Wbtv8eehMV3ZQiRr3hNILCAiT
kwaK/Y0MUiKFKGqvKxM5URvCzEnPC49dGFgMqb89PHHTC+8KFwfwoPh1sZr99JLyAN7uGnxeM/MU
o3MzRH23cMUaN3tj2UaqQwMP4zKE9FSqNoZ3SHSNjvtoUSE2LgYZIZpf5h5rdooABGiNpst8vtmC
8JN5u6813d7Tje62LlYyVxHhrzVctaSfzXwCdNDuj7L/g2AaYFqDMZ9C05XFhT/D/CUFqLBRxu7B
LjZnD97atZcAmkXkJ75+ecrkdutA+l+yT+v66s06sp7q+3YVUlfdbjXH7xgCIBX7mCvm/cc7Hha4
P6bKaGMR0xyLgMldsREIs6IHJvCRIwNJPNLfPuGV+/SUxD0xBZykN3WdQHUajQfa3WBQdteABhEb
ZtT4I471QUwgcpsqK/G7gkePGbgbBZ7Qy0QAUGnJ56qhs4KFWRTi7gMLIi+KK2RJh+Id/8UefBuN
GcAny3a7shZxmbvjFiimLH+tuSTUsBDAKSmCPzGHpEFlTfbECTT0ul3qsm8lDMPtCN88W61Sza+2
V9dtmaREj7vAh5P8kNvNbb/hBBSrqDaH50GKiZ5GrpRbSc64DP/jeIpkks3YK+SzBQGzAK6GXQUG
A9OYbwsC+jBfeLAMdAhXWeSNaBAKeS7EgoYdeZP2iE/WjmYs2uC/s5w5QnQ6RHDThY8fDpBpNzwG
ZCV5SntIlRD9FLHfi4cRrl3Ierw3RCQ/+ph+wdhG2ibxnAkvh7VRp5k2uuhz2RiI5x5+sgOGrsFW
/GdNrJbf+NkAQ5bNOZxUUNZKT/wPlvp2ejB2bDK/IxOcRNU1/beBlp5tW+LXG9wqxYnIT0MNb+34
fX0Jl+x/JX790A0ad3cQWYwdMidcPxAuM6w4hGGMzcz8kypLdM1WeAlDf4sQEy9wxxCSL5Zcj9nz
O/VdpG0Jv9rhpNSGCpbo3CKCaxlFNayW6HfoKu2y0XSKRfu1v/m1bC/HJEEUeb5seG26n3JTj+Kh
TIwuRMZjMkx3W6y3BxGYYHB0Xq8kYCPk+zvCjICjlTtGWAz/fVIC1CXCcY0hru/jWvuylpFQttGR
FGmXP0rbdnupzwD4nFIucxnOQ2xECqeZBgsJciGQtgoG5Bp4hR0NPVj0fIS+P6WMI0oIRqCmFp6J
rUXSebSkMKLuatHzPpG6xaTrIJS3A7QG4RlYrsDF/chhgq91qggqqAbtV0hOrnz0dX+6OYoN5dpZ
+50eFenb6cWc6def79DhUJF4oJY7+ixWr8boSQuen6mPejyBigYhIor5O38LEYshEtoep3mpGTUp
WHlv8/gyh0aBz592zLxVf9NfDXtgl/Gn1RBG+KW8YuWNRU15c7iSQpJxUG0OV3qgw4j8VEZ26kEo
XZFFEfAgJQLZVzgQ+HBonSfNsxXEyGUXCR22KLLh+EzCU74CG9hHb6aK8CRNnq1krkcwiqlwbN8B
4XINBGsijUukSYhzwvjpbzUXBKs7eKtnB3vDXwL8g6/1N+8ZYkxmcaI4T88CwCpv/tBQRkw9BMUQ
SIBsNihKBQuoa4jyyTPmslmu6JR08rkcxLg/ltP7yLkRvD0Vo6J2fvcTnjTlxyOhIZ2cPUDXIGV1
Kvml8Nwr3islsmVyaoDRinvfRRiMeHK3j9ZeSUauQrs1cZ7NEy4PLcqnwKlgnA3/urV5BAmcJ78l
dPxcb50wtQsTSjNN2FUzrNIVJc/oszLPuUK1ChGxKmLVVfLVoN6mFR1xtwCzVlhDEuxN97vwJO6O
bgGdJJvx+EATkYOGUBl3ypNOLd4ORbi3X/0/4Y5aO8OI0kZNhLN+YnzyWbFLS6NskUbDicWb2EMd
dG5Q7ri8CMrknRSYEoOuHH9UCr5BvhWTIS9T+Q2ho7/PtGGrLxFYFUFESdns6ie6yr2HQdrdP9CH
KJOr/DcN0bzzFkFNiTGGTD0pzTyF/7jAkndcF1YiyRbULuL4qLKuIQVsbLFp2hGJbDnOGmtsx+KN
oDlb4ff7/PQWib9sJmO1UI0SzJ4nGhIrf9NQemN/jxHlyeumIizP195UnWx72qHfHM3sPIle/yXJ
TjMOg0iIDarWTlvnfh6XTZfPw3Gm3fFXNAcgWbLpEnlcVJqJGitiDWwL7GvTl9mrlP0oZaGYRm3M
QPgrmiDbhFvMFXtHniGjklzB4rsqDjEfwyB4xhQOxWhpF2Jqg76vFmS8IVnENr2tiRqTB4C7C4wG
i0C9JVGxrpzIdQ6L06fm8P/ZnTHIWZqNUdmHYDIjxZzIJcV9+AweaeGbsEUJhXMxxIozv7ZBLFsS
+omKJ26vkXGTihyKo5qrViamtiJA1s8VH68sn4+4M7GCwk/nxetMoh/+YcdADLP8UV0/9Fm1XqQS
PpQ/iRR+AyDRbSvr4QAVpYE84PazG8Wpj6AOgaOGg66/AdasTXJhbYYf56Sm9o2aGBuI2hVGTDgH
KummMteeM5WN3cWPrZS6TZagb1Uts1Jk+pjHaI9EQ+tqqurKgk4sReXm5pVHEukJ5ohvWipUz6Y5
6X7V63o2MAbqBBcJQv+D2z8xSR58fGq72PWDk70p/PHnqGVYdQ6SJ9i+x8ifSf7wjRAZD6v/2wbp
LR248asYdxmcM+N71WoM+4AzLAqwxAn1DoOSqk6xwPEaGfmRUEh3XgAH+yXaH+mW7hGmeU1NySWZ
TPhtuWvPVY9jCGqTXlCGZWTU39LDHwH8UYavp0jhoxTCtUE5i49c/M1V85oV5TmckCx80gbYqTm4
sjilbS/pGbJjv30uMt2mPsvphtR8hEpdu7KBp7VLnjtsJeBtdEgHVzoma8JAap3Rji127xAGz1ks
MvZ6e3AOejvCpTzdVHycpgyhrFpU/lvYDGfm6qhrW/pmQBXI6hHWP+m7/o2XyI+yJzjFieJkyjsJ
aSuQqlEEdoe1YN/o/UkAszBUzovXALVm1BBycaBScNAlAkDioOe4cMbxhwmkLbkxl521c2SopAot
EqAg+DjUDURY0PBqUdkPjZ6FX5JZpr0Oo++3xoDFp6/EzWWkNXxjC2k2AEpFz6rCa/WWkeZfy3Tq
AhcOT9nsqTQUmEWh34RxNpL1Gi3JcjOHUEDccPuzyIZluQKhg5pYQhOZ6r8cw+T3hd+lx9nAV5hE
mzvMoyQnU0KYI1xE1ycY8QFNSCymoTmndKfpNAWHQQ2H3GbXCp41vufZshGF9lFwhdaF7EFKsogC
Eb3Flb1Euu6dWe1FaQtdPgHs6WkUu62ugeMwvKbmcKVxyHsD2bqEmYtg0ir3/QmDJ9T0DUKfjYSg
Ox9cOKuJgyD4NGvH0kQy0dQH/5J7A38puxAGnvVZwqSD3kDuWm7Tn89Gv4IWXCfwD2BiSsIMJOrZ
kiI6LrQna+3ohf5rJcKxeF0p0HEnsNWgANJOgisN1t6127Q9d/wsrbeDw1wYDB9BJe+ouUKKi5YK
zgQP0M43FOnPbIG2tDpsBMONL/9GIMxJI+bvqoTRVg+dJ+4Ij8QBmZcpHWpK2JuMW/Ir9JPBmpTx
LpqOBoOmaXnNz9nw1LEZouxJ6h5K0dx0VAdFxcg02661zMFV0oP0df2Fedq3U+Kq2m1bR7vYcvzG
sv1FVt4YnDxaumpNXwYYJ99UL+vn24kaaNVOrwnbSouF7VqgyUzsgOfw98rqKOqSsArTTHtSSRNd
m0WonIskjZDCm6jDPkiHq7PbCUI0i/cA09IYSKFeXQ0WvlT0Ri2Gt9frxfyWpVukg+GHX7xe/t00
aazrxDBeVnJjtAP7HUAbcWpfosnJVt3tAvBL7djFti/ODHeQwxX3xPuShbzw6OUHBPJMQYNmrPIP
jy8NMX/1NOSxYXyQDQhKkUQ9zxqFiby01aTND8fctG6ueUkkY74axVKBWbrrqyYIPn8Gr2SuNVjh
OWZ8v0689Nb2m8da1G0tGVsFeby+Vadh38dZmmjD4ZHaUEuFLWkj8kqX9xfJlhtPLWwf34g3Uqu9
N5rWG/Yrq/UfOcoOlSU6tgsC604p9zjoGi7cOv8p0M7KXa6VjObPPp0ImWpHyIZIItSC6hZN3w8j
ikokNhzgJrVitOKgz8mVCRrkfU+HgaBE57s8hdXAc28r+EW+KWQHutieCdDVOs7hCj6ac++HqM9V
KF8PhOCRFy4Jxgqr01kRdTSXjfHqDmrAYMS7TPGChKH1noZ6xqVeeVoVPMm9h9lBvNFlxz1+dDl4
IThUUFaInUgbDEACNPayu96wO4+5bkOqRMlGe9lfvsXokCFmeXLSenGWeREYfpd4Xwxv4g87mzSm
lGjBKyZ9wTVrMBHb7AI2mbJUASL4Z6+2gv/SbjTdweQlXo+a4cxt5IdRsDcKmHbx5KAL+MV3te1G
Ud5h+pNZrZ8HKomaqRlv0ZwEWRHCUkP/1BcHHM3NGMeLUqPx0CeQFUZ1W4qlzmHh0+k04NUAPy0d
YOvGVgpnFiPXIWtXE2KS5xVedS6K4kshYKRci55L3uz1kcgacuDByUukgSIwJ6wjHpYSp2uvVcaT
oZ8CNxHn12bsF4wIxxlU4o1U5Ie9tdZjO6zdAmZLxB0+ntuyEHmC0R+saJnKoaUsJIbz+UZohFM4
QqNORDGJWEFWJnWX8oGqrFH0QBhGJZJAbLamwem4nSpvXGiUAGTBByz6FghCzhIurra0FoUZZTQI
Xv15ofcHaOGxCkq650AER8eubaUzwEpvvx7xvP9JsRAQ4qt0XngNlhuFapzYupVvBSQABIPTflQu
vbIrPyWz1Emg3jAFhlI/JmyhCoZ8t4G1C8Cl3b5oivceX9bLOgrC4rUtCo+FdPSDhI/hfYkKGxBP
Krl09iOyDuNTdU2MHz7cHdWiQCxNikMh6GT59sebTzS3EBFgOi6t/vkz6l9QjHjdJgldRYjpydiw
uM7mX+OpLUe1GFyeSKyDOucuShijZAGTnd3y8ItzTay+GW95K2iMa+qzSYf7cBsBUfGlUN50fC/4
zeDlRkpBMVan24B2uki7tWrJY17ZciXuZO9R0c4hqo57aKZ2iEW4G1CCNi+Yhw3BPgFVHAVoG6Pf
t6glFJzZ5c/o1rt+GT+O3sSZuJ6QD+6rF/IiBIc+vm6YjTjJchJTWo5Hz3VUx9zVSOcceDAm6DlO
8hxIIT1wGsXTEkFTt3HKVMwnoID460OcWHxurW/9BpFPqZMUYn8x+fwUc20vlcI2VolzfnjRvyKW
3bMqL16QYHUXTXhKy+P6NE+mYQQMaLoVApFRD504W8v+TjsoBi28FNK1xENqGfr+3IkYzQU9vT+Q
w+l4gA/5ePgOWpQjsck9l83IMWMZ9DR3Tm3PfnVvHvQiS6Vt8YyvJ/Y6IB+DU2nRLpIDmPK/WB4t
tysZ+OyRdV3WWbfuEoHoCCbOO4LBtYocO7CT9p65PqtEUGaCxLeJkK49pQ/h0eCmrtCf3ZnJDnCO
lHherQi+BHHmoUcYl/j8V61v2c6HRd0PlULEjmH15SNq+RHA6FOPLZJlqnVgwDi9HD8UBlIOHuE9
9NYl/Ay7rAr0DdA7MZpXnNjJ9htb/QM17SwUiKM1LM7GSVDkOXfULB6wrYra9/AkDyO8bvcc12hG
hR/jQuyYpKDInXRyeXQamZbImcL+QBNwUwAsRBXAxip/lztN82rJEzUCDMoLOsmmdKeKKyj6+vd4
uW5vBY5JwOIiY0RvPpN99kUgiQoZBvxDFx8HQd9jfTvc+fS1a7iCed8cpKN4/kSP+gjeahy6eAUk
t6BcbAfyhqmXMeddIhAc1tURda+GcqmhefJHkId0HZKd2AiOyuEp11Akl1LdZ+wkFg1+PX57btzK
NeXpLJ65V58ihbHzRSXvH3oTib4NhDr/AceVl05pN10tTphQ5VyyKJwfK1bHsgHeNzD+9NuAoJat
jOs2qM3Ioysap9uxPIlcpbHJWtEc6O6qQxlAQqWKXwSimLl6pjize3aTU/iTiEKnoH/Z4/acVdWh
qZG/oeG0C3Lao51S8sssXY/PdbgkSrolWkF9u8cQ0Hw2b4z5Tbj4GyyrtKLUXS23NSXBkVWRrTQx
IJnPSNGnhhEYAVcfQO64xCEn1DMeAPqM13GGRT4grYP/f7RiITjUE9hoZL/Ea/XYqpKSjQFVsTtB
3I7nV04aAaUZmEyGyFwqrrou6wWkZHnsiCEAhtSMBwEybv180lAoWNh+pInCiWgTS7jcxe0/Ay0c
e/1RS4obHvdreWql6en31nDXBXiwpmB+/fnM9YEKPL7hJmgarg6/uJMGqbGioziUfofv9w668lH4
ZAg8yUAq1GhQvDMERHoKwcEu/a7nM7evNHG8QB9+QWHllwMKzgFpUAVYdkphu1nqsyxRprP3x72Y
3NjkEVzsbk13cPxSxFme1cgkNDEHLf9SKkAl+KQ71QkfFV7rEYDY2beHyNHbOBfDXDTppQ/ULdd5
SCSIBvXUElqVnb/xTtNw0TLSS+niztlCUhMPBHKqUZJdV7WxiyBWLaXF1YVc5ZdzSwrgSBX8g7w9
TIOGYBwoOJw/k/BkEpeHRyMWKYlHDFPMOaORHBZmdcq56lZgBe/Mf/N/15h691GVnSNHL3mEguCa
uSkVMgH/oUO/Tm6r5hRMTc1nweyayoI5X9kDkOvlUVsAEeox20/6LrVJ55Rv8BlJzS0Vqc2Lzc9W
ijPamIRkzE70WOrE1C2C1rkBmOe8Zibexp63tuPBKAubTWdnNG/diSI9Mf1wiwNkRCCVAYVF/rPY
8eVa9XtdiPJVQNM4iNQq0n5xGDdydJoWm/dt6Vy3oo1mCc6D13hTUnH7Ewgc15LyJna+DTuM15mW
TsCUv8Dp8RQxsrjimqUNwcPl792jujxgdrfF9+IWthhCOzKlUxpcjLKQIiTxlQ/7hE+7cLkpQBtC
JMsuzNY9TT9jwmIx/j7RGeBQWVdSQDE5D6VLc3o35+vG40SA59Tandah5W0EXeS87O6iJY/A4REx
GtehinProlmTiAkTwZ2KW3pUmgybbKeCvIURVcfAkTrvpL/wcx8sXku00s4HjjxoeLCa12SrProW
5VDpqQOwrswH7GjwSFeKRRnaJ5+a+cjl8SEOA1PJifBXjwmPfidm5lEzPLJNwcRQuRAisTUCI1yi
Hrwvvp//7bIdXuaE830uvq7MTmXw5zgiMOv2eYzZQkTUdZA2SQ/sKs72wLtJ8q0+zS4H+YHrSJye
mslWSVRSNMBPoIa5OIbrrD7AzMBPouLu6GOQUht8MfG/SbRqvlJDOwxYBZspDN0X64iinmLR7p0V
KSFqYwwscig/CJytWjA2TMsqv1q7lor0RoOHJLlSNqKeCV+Jc/5SxrSNrFeouy1Syuw2fWBaoAeK
Rl4B5JHQkCzjg6ehCZjaUk5tP3WH4JNoBwYE2VhQfrus4wZ0K/e9PidlOW7zASDr8HuWR7Frwo6s
C8cFtwRqNJ3/tdlwwbDMLtrssiBhlDglIugxkcbxDPLOXjZmnbm7m8XxmPKBtKUSC87UxqJckHMb
OyModnBPYhJdaE2Tu43YUH8M9fnu7JANLHB7ZSptadiAqakNMaRJSixDsZSmua3hni/ZwJAeykPK
YqvngNCChEPSCEcJkNrctEJqJ5OE/k7+UfuBTURHOGxxeGaK0K0xN5UK1ClrJ5TO8atXTaK830mU
kZ3J9/VeVVPJ7voA8PHl6L70+fPnXVoW8UvIqMdYykYJXDxO4Djk1w9HvSLiEUizLQ/lrsDKnqwz
7ZrK6pKLMKOGrSvdj+gzRWSW1i4AsZqqJITuCyQytdbuxi/f4Ryov0rD3LyevIcS4cKAuMU4VU1q
ZKVy9zXZUONRDqyVybo+u+rZT4JSHenfLbFZxytMzU7XZyRGaCeGwo+5mKk+QnByJEhq91MGloBh
4Tnlmhpzk7vn+/JJlQu13L8x+pOeduSyTSoch7ilddZgHl+LcSuzEG7Bev8MPjuBD8ZGQr3sGS0f
nPmqKow9SnaO1zg5Z6ayfUOYuHP6f5nbTEIEF/luUyxBtazSzV0iu5P6ju3cfeWjBOUOCT8XG0sd
AEX4Xlp+TRtfvozU1lOrjCpVBXS9fok90XIV8cQ6EclvFHptjCpvKVT75NEY1vuJqKaV9pE+MBa9
i7WmjMx2YbypXcORpd6ZdiXPDRVHWTiesS61dItGdMML6E2DTFxoopBa6JCPPw085+ora+GZmDig
Ln02jzEnaX4M8p6QdRG0ll/z+YP8jSIW6AJKm1NW+BicLjmEPZKKL8Dgw4r2vGxFTTMnCcRsLOHl
klB67XdMVvde51RwEhWbfQWze1SpCzFx4LwxAmUjkBCTj1VvM+CIp0ktaUzNdW0LZuQMvYuJRPO7
A3mHStJk2j5OC47Yr9bP6q2FcwKGK5auCl9ZVYyIaCKeInPSSLbdnP80dNkDm0mFIU+wgr/O41Ik
6kmS9Nj1aqS0vt/NQVac5bKQZxr4SJlIgkC4zI9wQft2DAnGUx0ZYw0kODzziu8q96QCt5g5/816
0QWxvihP3PTF8rBR4LKq7yMDKUaY+W8LlcBAuq6DFDq697uoUAPMOhD052RDgpPM5z+0/a11JYKc
l+pbx21YOmTHGwnZtfmvVNP0VAwXt8Ng5dXnIhiQieTuJupGtpqiYXSsuqE+QM2Vd6VINty6sehI
uTKz0xBJZVKeFVE54icXYskRgqfUgT0+KmEN4qKHkNtrVbHQbkA4B7Ht0WZURC4r7LaOMY4/ZJBc
9vT23AyOt1RIuNMwR0hsM3yJCXC4ythWns270lCieFpaR1RCmwoHiO4+HjgFzGJg2xLIlexuhDmG
Pq2gZbOV4n+BfDrOwE2Lv6++CCVQ0YTiaznYXyA06PmScbq09DzKiJDLDDJXfw67eYrnKNaWanbH
QLDtyDlm8M+QrawFJnLJKFGIebQxFaD6WW8ycAogMUb8Ftqd6DKIXpslAnr8/FRbO5T40CjF7NOl
WdJ06v5+V/ujBqDm97+6IDQAeaZqNpbCMaBeOKSaV/sPuUgXRDo53GQ+uHkoc1J7qoOuDvTwiaFu
CSC1Y6Y/39tr5oIpjV6enSLgPnyrzXb6kZ6prL4njLO8sppc0+QnS5gfj1RgWTS+te1LGu3Iurqk
U9y0nVL2+y8hOorh3woCBzFbmWXxszK+fwsX/LrpaDCZHKpxGXviKHT/f3WwxL57yblrFKy/7cRs
gfxmyLjaaXgieotghiXYVSiWpI44e+Vu3SYBupv5DFI8eZMHqmMJVs4NX2ik/Gr77Cbvi+Sp5gj4
CiCrRMCNXcFauTn3ifDZ9ovV2pVPBQGCYy4EREuLgxNOKMJKz5R+ilpfqfcYEE2oZHgZ+SjFSVhe
DhbSmgQ9XNpzaX5YaCwi+aQv6L2cUVp/R+cwLKuYPHJRsaExjab2c0/9TQA3pxGeJYMqrsN5HKg0
N4v852BEf4MuarDestDNSCVFNwc5/JQsWIl//AZUUYzib2MTQXuxo77cUMJQUu9SIk0CHS5XX4pF
V+v22WblWCBF+Jl/6vo5XntCsqL84koObwCciLPqAvLAitsWPHwIHtrsOpQGeIwfw1+dKRT4In52
whqs9d7tUV9YbvcrHECf32XJrM0p+gV61LZI3C3h4Fq4+8HcC9k61RIKWkJx+qy37/6Hs3xWlZHK
VbhDLDaGdbXdrphskV+GII/sCXpcHN713mw1oGEjvhbXUFA6uiGVbEriHtYMTiDTq8RT4VR8AyV8
yKer8BMq4h/tOlJ/sZZNyIn8ZO3oS12EYKAYLvxWmgZewbJOxSvClo5rHwPWuNcTdcqBQGPO0rwi
cl1ox8m/SuRdJu3C9D4kW3aSqvX7IDicepyFm5NEYHibBFzX0YRWiaF1OijiiT08i10gHU9JYwFV
dWS5yvk9tDHJEdClfaxBl5EcRUl4mR34rODyFAmuve5ek959DaI/Xqt7/bJBOduPNA1YvN0OdmyL
TA7pLy8WQ7hfurXbJQNt8S9JfrmoaUiMxmwVmK5S/h8R41bWiQNOd/svg0kv6RUClwVGWVLXFVne
zLGM/nML6/osO+ngolgEheTvGJUY9YT/AnLE1ur8yTXUnMpohkc6f6jQ+qMO7jJq/VZwOlOgCHTJ
OIZ9SwFufZo84ZcNClvDveQ1IUhSjlSjakPkCeP0kYRmq0bTyApvVQK2LEHfBNqypMiYZXrVxJ6h
CTJP57xTVZ19DbYogqkgXfzzzrRTwh2DrVmgHR3cOI/RYkTyz1WEOVY482rmw6IdrgXxQKdVadie
+KLVm10j9eNcTp+ceHGj2ehJDaFxWWBqhHBFkhXHWb9+rwnBK3CPYMg57vgBudZcV6/2OxlnKhL8
fRuK0rZg+wGwF0LaXhMR6qZNdPdxSsacG3yacYqaFo8hXV7Ebf3k8yMmKTHj8yj6qbdVMcuKCgVm
MaFkxuWLa5pEnVyshvLKCLSxdFMVpn4nwPGhloXPLYAVSL8tegSZCQfacoF2wSZtU130zWlunl1A
/c92fas9OBXViLhQpDx+mtyjnzG/0aSKUBpVEgQLoRIlXvY3rOW//k2yQz2sPd5LJuFJYBvFdWjA
nzGyKnXA2nFAJipGCwIFzZA3D9AORy1+hODttlLMz9kU11LqLHk8f/5hfhFbkSIdpdfcKw4WEH0N
W1h+i9VzbvYggFEgt9k8ykKWetqfgisdWoZkeWljmM4lhzIpXBbx2iCBN3TJwBiK96/1cH43YlMW
lIQjj+Bofszjxlrrolg4Z94B99i1/4HVeuNz3EbVdfM8EyU3tyPEU86tgzC+5afDrwKRtwVdCR0l
NdWkBwZqsnpGgr8LtyXDtLV4QLwLAsd5hkSl92kOnnowgCz7TB0/bWNKvfqMUaDBFkwGJxSrHwJa
Z3EKETrubh8enXSP3jVA9IeDOV29B3KHV9aDYUkzRVW2CDpQZ+WY59WCYttYcOFtixc8qOYnZkEe
Wo4ec5ow+SDJDmq4Hf1mC/c/NmxDKqfLUbMdxOuTHn8ZAidXimGwRudhC3MuqWer0A9s6Mz1EdDq
92pnyYScSAa5NCqW38nzMtuJz0GdEtZi/b56vJ01mPZhDfkDETo2OUlW2yqK8bZ9hJWWBSl809gx
3vSonKBFlXujABX4PqMCoBGvgzk1nU+4DQgN7hLzWUfB8wPOjVee2UzdeJGvqD9drixzseMC51Go
i1X4fxpBpyaMnxm+f2Z6vWkb8Bu2lfbmceaWFnlIQUS7LBTgsRItpaVgw3JCiU6orZDr/Gr+r8ta
zhta1OlkSPmzEJgeI7ixB3HIg0S1FdirruurnB058uU2ild1pCD1li/XGvu20aTLAPqSqXZHypEe
5kTRsKHPbWG+hUss4lyo8IUT7n1J8Beo7LFUc+T4Js84rCKwWete8zp6XxMOZVE6DfKqeCF61qhT
4wzqC0qFN5ytLbeAFGUnmExOzbpDcHvmY6aBCvkt2qDE8ksdMM1NAjNj0ofmoPWwajuMgv3i/6BU
jCvhZVaxOjjEpgkx1sAnO42+5rVjlKCcWlxuXHEKYuqd1gs9lvCnd4mEpEBxBTzik0jPSouPvP3x
nj/CeUmtAxURSLQK4sWMMb0ZWmgn+eEPnBfQC7uXnBbnQfCo6anPMwvS/hLtZCQf8RiVPJgPubRO
sR2ckNwx+MNKTR1jJzuED38esez3EPNz381srMly3FH308cxJrlbpeoKhztEhWGJmR/pA+p83uaz
yKXsZff50zGQxC5aG2FwoTiiUIMhs+HYZdQvkDzx4Xh6l7sc6ur/jNnsMTfzBglwGGh2feHPVelL
ez+xOLsqQmnG+Yg1hizsHFVSPV+GomoMCBRtwQhMz3BelmvRpgfQyKHJrq3GKbjN5j8xuoIEiJTg
9BS61Ym7yFJM36J3HhRUee0YpCTjRhmphUFyEKOoWqHoJJMyy5NvMmJ1kNEs2Vy1sQjYd2mdCWhy
gGccK8Qt8M6sge084DuhaAceCVFVddVSZZZE8ikZQEg7fm4sH47UwNZHk56T/bLdYgFzlgOtEqGS
vDC59oi6oBKwX63XDMuuy7S4AimW5QTC8acQYdn7h5GsRK5lrvwJ4mysyJqitQkEOR//nisNUdsk
aYGOxExGBC0Lqu2jGQNm1Hi2kwxf/c0DG0+IuN2CgwGYTj/pOP0Zv8J8+mVnd1bLEg0gSJC7WJC1
RuBxibd50ds02Ld8DutjNZXmkXTBgxrD2BX1gbEsVuAPtDhreAaP3G90W8WJXkFF2ilh3W9lbv6l
baj/LcjVeP/rgiTJLy1HMcq6DVpG898ZdSGAOMuUNnCqID8bbRPfZRNkTcGXXBdEUueZ/ZPdHbar
g5ANOnEsZPdntf15BYUT4s+MAJ+AEAFMBxIdRsSsVCoJDw9ISsfmn63BfRYJa3XGa9+62qIq3Mmr
DQItwPB9MN04dEiIlsG7uTG9yyQDh9Ddb8shU2Lalag0LXDAUnt7XuZPpxtPSbcx6MqqiIx2WcXT
P5MiT2M6jxscPXaL5xkOo1dHzX1Suyytd1R9VmIwdMoIDHw9YVjeZyPCj+AjpazGmPH6dXLiDu1J
xRD7RDacGz2Oo0MpK6Pm28futFzNc2wbj9wVFISzOGbH7TiEG/+YlQlJt6+XOIKxSi68PszkmjU4
VrfFtGxt2PNqC6rLnh/MsjmhhgC4cbxtm3Qfwo/ki/1gtcNbnkifEj/Ba2K543u52WOrS1BETjQ8
dSPB7fHzGYAMCWNVVIkZgNa/SaStyfixKGeSNHLSneDFRsXw2r7fvkC8ekBJOoD1FkbxGhNrb2e1
D8Cix2erjwf0VXJLiMou3Qvd0isR3ToB76S0tmnPdvEzusXHMgFHClCrRu8XZfgCS5hOf6ItfKzD
9KlLbQWEdBKVBnHRrXlfROsH87BGDnrgD67v4RJ8YFF6/f5bcxYvoRLiR2H1plgJljGJ8CSmt3cA
9JbSYGDMHGhe3Z6G2bpKY/vfkRwquOBiLN2zHJQ+UGze+5sB8ONPTSagIlrE8DtdH079P/G6ugZc
equy8Fzh+gn3gR5pogGvY8/txf8D0vUiDiT0SowxvCS1EaI7WaquUb6a3oTYKcuoWDG37DSHfp8x
UnBEex0JThVi9GJALejBF+nWbQ0bjyvyBdIKiNJ9zeqRUweuwkj178bucF7sbwSRKQf3IkTwA/x9
Pw6cmGgvZESG3MXX2pdB05vQ/kxthcoqvoWwYEjSC1XSvVgs9rtVlCdZ1Szjk34T9VCxstFQSHzq
bRMGs3AOrQnZj3e/1d/DX8i2srYWxMWIHTGvigB75qMeRSEbZG5saWyPn52/GBKILFqEAtJku7YZ
r5Bb7zdeEHNcNC0MYInaScRsNIx4Aw6XGhnoyVTfZXhrH5DBOjsFr0Lipg1NsV5B9wwXFmV77rDg
BhuxW72Lk9SEj/j06EirYPARpB+5lPF8G3MpPOGRVv+XuVSIMPIVNalfkzncxiUh8NNHhZEdomYA
2s7GEoA1pxeAnszi6qgpoO0Vzf9dwOxTvIKIMSHt+nuu5vXb3i05kK4Bu5MEkP4dj7Aavy2jR435
Hd+N+l0XbTrmKYKU5HvA9QKrrRl2pgU5RuwhaiSEFF6cEzjZiME4Ve8a0u1GToAZNDSC4ANuf0Of
Yo1KIZGqFwV4nuhEKLP1SJSXrqMYqYQ8ekm5QVj+53xb/MYZivXdyb5eaG9g9RVQbI2+12jsDg43
whGGKkzvTbuuThca4p2ZkwM44wTC9hYXAS4GIBsksMoHBld1uN9fFNb0KbyiLwUpnUiSjFCOqhMI
5t3b/aF/pFESsdBDYPs2JcNV7SEowCmmd7X7WOcvjgA+kpVv5YH8FIEmB2q8XHPaI87R470MDps8
xZhu1/5dt0GMGoGjW3GodQXi7AvG7SrXMFUdib/8rY47QPFSq9DO+Ku2ZYv8rd8Z18VC75eiYYeo
h0ZYKDZaS8qSoRd4FeXxROMa4jFZXrLu0tyYzpdm5x1PQ4/7QpCe2tIM8qQ9aBq5J9M4Rv/2uuN7
PPvWWXMMzzNvDO2xyo6C6YnZ3oVT/mINDv2GThvohx4XHRaSMfabQO+NRUv72mpwOZImPO4eaJnM
TpeEG5uTggrhyseTUJLbS1VKghJcinIYZRRNGhMAZpggJfsw0XQbse1DKzZYANnweEW2HE2Y3xUO
sKksgOghPo+xg53mGNfnjTxBfgMlbUvnvsxIZBemorUHXawMTASje0vufKaH+xtEUtKM7v3IPzH5
YNC12mpVWF8EZSq4GVkp/erXm5oTaO2Ysd4vUa0GpbKKlVUWs8id4cXUqj6w/DxgB+RZcKTvHt2p
mL4QOB3vaP67q2S8gS2Ke6ABx+1OZ62Ii0THs5xNGe4OUcBLiyUeEzIYtCRXR2TJjtyA2fAf3lbO
5ffRlFiH6zbZLtJsNWEl0UlZX6/buU8FYwLt4IT2RosfE0PiMIfcTVCjoWz5kWO1kAw1BlZK9cNj
9CguPKhvUDO08+mf0eYQyCAlefM/Up2IusKuTZg8volfrhydUkA8CmFZZa+mUwOTPoo77nGBhB4X
E2r31lhrfLD8cgQINsFaT+g6sUYJ5/rDZqZdsPcXdeb46530Rw1yZaGNgWx819sId63/4xJnxeFz
znNSYBZqlaNadR6gHlhhmpn2N7nFe1c7zc2Gd93cUiul5h5L1JT8W1AhRKE/1udzvuCl25j7qX4l
FrQ+rM4pLzJfaNSYVRRkuesYp9MWJ+CpnHCXX7yj0hBRNKAh25aAtx/mM8nfCcp1IUp5cWB5fElw
mP5jZviDyz1kmknz4V9rv1tOaokkag3XHvse0vhN9NVsZHHtZlcpHBeQObziV4I35rOJir9S5og+
XcMGOx66XRIGJBhrOYs6lEUx+4N1y/AQadO2SJkXngMpjD0l+WzfYnIRQj1nGgSVGdhFL95Z+yGu
TgPHN+ERJ2K4P2syO90la43vvP9QoZKEdwW83gDq+NCJY43N2WbEI7fy0nzfgDqNeWQfm1CAwqyh
X1xoMzo8SfQYmCjRkYVLFqV3QpyZCxyayOXTsMBKZCIhBh+EfsaX3Qh1TmeKroTEir7MSmnX+qdw
0ErH8EWhoo6dtW6HKmVQ8FNc/MUCg0Aq8lcZ2jFryyHAEo0JyjSuvZ9sz1kHMvYHKY87yhyG5RA6
okane/H9MtBI/LPLOq6Bcw9bRpGpWPr3Dlqkor1MX4NUd3rgfF9Hvs0RFFgXI9LAtVwizuOwcRAi
GLM+rHUQ7i7PyuOMMlmtaHdOyvITjButNWOnTbcN+aJihV3VmMFKQCdLdWGm+V5wgYOcrLZzkwed
orhJ3vXgLKrpKvln9E6CGWE1KJn9P2brZCTRKWXZjq+I8rVVVIXZkcs7K68Q8XNggK3JBevqe5Uk
pKQoFJ5pG1mo76cTOP/JNs1+DzNsijciSGftGfaOYdOi1loOA0TlrVySA/i0MfRpCIluRyrqiDgr
x6qURdMCT3CabfAEQ94yku5BVCC9qzBNh4engTlzAwuoVuZ3ZV6h8OkCDpOZqCrXRYcllPb1A91t
NQeTh+GCKEbeoFWgsp7bopLhXc276pJ6xLGt+m0PGPRhHkTqQlDxsQ6WX909K4fV8RjT+ywrEmz7
/am5Xw06c8zH1pErb+WUxNSFXe7Tq3/tfAK3UPKo7ELUwYzbE3qFtR0rT2q2S/ej38ENHyOiqQnB
6nYDGD17GPhVSW6UCDViIXvPjlf8Gxx6YxygnFuO6/XdcnFLHdVEMD8uHTe/So4yHAwYm67L99ej
87A6HCg767mUYNc/Tv3zCpGScXt680kFNX1cPlo0N31SIbueUCeN+QzOAHTxNF7xl3ADP7am3/kS
l4FU5pDHLOwppN31OzlXiUX9zMfV8HRavfcrHKUDtltDWXi5uQMUrZS+/MAU1yEfrDZAeXhvsRIj
4/Flcn9ddc4brKvCBvXSRKeUW4K1jvc24y64rRP+DJNaAuoMJUrFdrpfZzDvBiSpvZCG/wja4VeG
hU4fL5p2xg2imUSz8osHCz2GvDvOvvYrbBTO29zLA8rXv4chEh8vFGlyxIiWpSDNiO5e5rD/R0xj
dh/nHzQG9R+VRd2AAfSxgLer9TLLesCElv980HPvgVqJ1WhsUkXz0Mgn3dd0/yDxiQpNu3ySkLWN
J8gfGxF/aEKuv1Bcat+zSSHbrvcjwTl9FNHwqYYXsYeOdLEPqQfuCPCyF2uIU5Ke+WVnmMhvgq+q
oHiNlcEUIEeuu7r4m0+q6Lbhx8Tm0ASb2yaLkop87b+q5HIDkQdxfzE1lgzFB05EKyinBtcsiZR8
ONi6dHn5NeYuWz1NmBNxwkRDU/fbXI6LVGFaf6a4tzIgd720AdFW5fq94huXsFg2vKZTx1CODOOl
SEz2ttxglVatEcIUpsjSacczNOpFimKH9AZvoTzG3QOmNIx9hIdXLfVU9lUXe8tChK/6+PZVrS4y
NWNnnR/SGHCG6Cm5nI8MkQY9Rdti03tlKMl/Y4MIBXuGqYby8JyQTg1qbo4M/ujMf23QxyFXvpWn
drlhmQj5clKn3F3cRLPJU5M+nuGvIGo8eJ6lKsfH2xe6OVNhIkZnzE1e+M50UFWS4wjKwjNYxoTJ
9WdHeUrsNdGi1rZjPLGA9s7KQEjODPDjpSut9dxPLsez8I01sTzBP1nYZe0kvSkhUTQXQIOL7egZ
55iGDfe2psJXMPMebc8eFQbZRmdGz4/56dRnzKSdsFHiWXbpqz2lW8z7bHjM4b7wt5h/WSLejONN
MPsb3/5rwqWgFR9HLYJXMQQoR5oVKm1MX8Xhh5QhRwO3u6XqopX0nvxzuuMaXh42yawawfT777U3
A74mtC7XWoeagwECh3V1NS1g+oAX9WaK2D8vVf/nCkPevDDuhzBc0552O4d63Xr0HblisYjICjFt
+juclp1KwjnEO1ElOIqqWb3VUg9CrbMaqztKfNghFhOTsna9H8+sXZvZ8fO7x7G3SQd7EA68c2pN
1Vm3TaFaxY4zUSbvH05YS2Emh5uQ9IAR//2D7zAWoH0kXkBVE0u+7mEB0Y1S9BYSP6kIHY3NEqZ0
ICCiIG/1tOps5kdaf7zd2w8XI3l3+rWHYU0rUuq5X825EWowwYi39a/Ky823gl6W143GBgxs4KN5
dVZS/81oX4vqrGU/SyyNwHwPs5oPneBsIUzhHNYfsgFtJ/PCJG4Ul1qb8l57EW4lRv8PKH/5kkXD
2Bdonjcd6ctcD67S1r7Z2A/V1TctzkGuCi8G3JGuavo6fhPuJFFMSvHiShK/xwHy/Iay2qZWbEkw
yDTu3NqeAf9e2mvf8h/bBxLLG2CATfugVwEPrqvEjxZdhecXlQR9wRpzTIh7Z3xk0of19sgtGPKb
Afzwy19gqB4oqO8x0arl1RGXadrJG1vmL7tQy2CjH+/AlGxO2kJlaCweGJLRziC2y/Cxfn+5Iwrp
UVDjZU8+WpmSg7yJyF6ZB6nNalY8TQAdH8F2wFVwauHMOwv/leE9JO50CaXkGGAqBVHlxaqL9w0t
nr+pISCbybeEkGsdpBgXWJDY14nJL/nozaCa+vV2sot3dMrL3Xznj/tcBqr1jWUajh6Nph+KkhDB
25z0faPVJab2YSyFvBHwgc4rADO41EMHPnXceU1brh20rhYITDBq5f4Gg6XTUKq1dwfPLurDVVFI
4ZTQ5cyLAwo9VwalWCpPSZV6P2UqG7/S3ghA7C4bMgOPow/iWN83uInUjfRshGy/dZPa+F6torws
jVmQy9xHcPxg3QyluyN8FpYjKdX3olfPR/SEHmdnB/TuvshJvkvkMDM/o4mmjJFpVus5Pjieyyi4
LHuTjdyX6RmHzOuNZfYvYyudMQw/xTg+uuh9RFF0di/4ZYvAmEPnph6P0HEzIKg/dA6HnvCyV0RW
U6MXxpIyVZHdYXFn9yOHq0aUwavf/ozQkccA4dDFPF5xwXZrWUy4wloNX7IwWS8Exi0UzF2LA89/
8Rx1EmaXjEMxqP2aPmREnAuhobwK3OwNKYBQFoDBtS54thbSYr0J5GY+1TdKfAJol5yDIa8JOflz
3oBVdsdGIladh7arJwAY7O7bBKZ4wYYXcbHqG9wZPm9kGtW7/ZgoJ+gA8A/qFECQBj15t4gAAuWa
NO0G7mHj/6rnkg9k+vLJuVgRHpsi26eN2qbh8MSpe1mPr6vTMSNSvkZNV/l0rf5cobXbJNyPi0xl
i4MGMLl3SOI61B3FWWOMGMlIabFEr7COWiJ61oGFEkf/i6yu9zdc4BdANgpj4zIQ/llyECmnuTEl
+edRwCWYhbD0xR1YggBEXDcmsfCya3C9xkEOan0UEzjiNpyGXmGOnGa+FQebQif8VJtW7BfBy0po
tjZzuchdCQaKZKblqC8RV58bV3ZJe9Aj8qx+9GbjqrTyByUk1FMyp7Qs7NTeBi6LqkeTNklX2qOM
C+tqRriIKlKC+/HFdumAXw9g7I/tPr1z/+zov2c76Ft1ke+XqfGC3MEAjR2QwvmWGfXEshV3nSpn
l9G+twmDAtySjcfjAns2KjaXqJrUlVNSPmGJTqaVgoAMjuCvY19hYpqWQZ70ZTnVdaUhWLrsUPCM
cytwdcC6ScnHsKGe1gTVeO+pdw9XOfMY6zuGsKWwr2MIY/j9S+/aYVlvJ+03+q/Cqw+3RUvvBChe
ICwv+9FhAM+hAHAEcy2AnH94H7FLiZIb+UMk29QpMwaQFqNT3Q1MGh0CtZBbs7BeoYwtJsCTmIh7
j71RUflP7OsG2l+0HZW+bpIRkGPUkiW6uiYwh1bVrgme9oR54CDxMhiXWy2K89gh8shmvbsZObk8
1gg50zJQjGfaHc4MO4hEq02boLNsz0JnJFpdBmxmJz9GdpBfyinOtx6yKBixzgb19PsawEez+oqg
EDN7CZOrzumHga0w6yYxigYPdfnoxq5U1QCRNsILThmvcqEuXejiS8TEmM6WnlFgM9Rz+TjiF9QG
w8RB4j3rY29fCGoxST3xi7Lz0eIauMsMqysMGzjoW/Qzw/jHmtcqTm8z9vbxFqiOBdRdOorMoe+C
eU4Z+h/3I7T6xsGz8X9j7Ct/EBArgPVi6vKXob3mVtoQ7uivG455DLJ05RFUpwcSXKGu/hlLNa44
I1XIFtCmg9YmtScpO84gh853gVv6DuUG0dQEh2mQ8+H6R/C4vfc1S45Q76DPGNbW2aD/1KLANfxN
KFBwqAiJHSDF1SjXIskP4M6ZjbekUQsmDiykjEWdzKiNKCT4EfGplsX8GFZESGwIHvWP5KMtkEDc
1C8oV6QYjOAuQEq3GNoVqvpVKnRfW0Z9Vk1iPXWHk4MeYdNylv06PoDn4FTP2JfvV1eM3VxMqCao
im4gSxVAgYpiW4q4RLQcIURgLapMl0goje+TtugPXyWhc8K3LJtVlAP7U6ArpNR0YsQpCPHhcaOi
g6p2YIRHunhxH4GQx0m9waOXNcUt/M3nZacbJjzhaDo79HETcYmbTjLFOGd3p6r8woRS6nEispEF
DoT57tmcs+KBDWqOgqmLpLjU96r8bdkvJN8oAne8VFoxb3R3VUosjfkp5f8OozjgrCUBee5MOnxs
jRx4w6a6tA8GPMLExx05Rd4+Sog4LeGFpyVSmNfNtazwh1q4koRSFtnRT4nYaMxq+jqgq53VDAsP
br4fmPOy96Ts6jgyEr7keqqe0Cb4tcNyZC1rr0be5cizu95hLpnSE2UZzCb/+/mWY+RbWdgcA9oU
f69bE4lnDtgWsnEVsCJ73yX1a5QBV9Tu4n7hgKrwuP/xc+4u/q280iMEZBkyfpMmaY8wrVd2IqMZ
8sd5fi59701FEIfN1hh8yTCPFhV+KsA5ej23Ytz2Wgb3drhfy/gDifZrNZFPmAq6sQ67x9rmf7n7
ljgCXsAjUXAIJsTy0p7VBxZ8VW+oo6pbEa9GZTL0/3QafBjLEfajOWK6paWqIsaKFB8lDI0o+iJ/
Hd5ADHcbxvVL325Ni9Kk9fdzK2YaZWwuUNajEMVUhAX+kO4anT6t1N/Qs9K2W0lzQE8W5G0zjLqn
eAgrWtB+BpUDVbWNNsL6++0gTAj62SHE+ZZgJPPAhE2yuyuntSUPVNtMqHXpnkm/MqyOhfqgy9rC
LQ4f/TAlzsuS/x+maeDaUoncmgwMHBJYZtzwv+joMwUqMajCGa0ehmTjaD2eYuv68acd3pPxuqMG
QhIr6HUi4mdrkDD3rs2zuJYk5VNGJRLlIEQPFAYWtKnH7YaH0T4jEAhjhOwqUNgE2z4h7QXomF8B
rJSIPcIoAgnkuRFN/aiJco6FKJ9ZJ4oNgHuVR6LhyvbVt36CSyp3LOfDmAS0WiJpExd2yrQDLorN
xMLjAJN3e0JbaVtNUdgLSYXhCDML6EASaMAruPGsP5ng5r3v2fIheJW6xBqvww8jIwFoS7HWaEWX
iIaghl9pMc0iZFRmgkxMTdsYwHNqZDhdEcgsJFSEXmhS9UfrQgO8hsvDQGeWSk1Ae67vslp04Sd9
j/pquVIiIWjCe9cU9iKkREx9hv0MSrXH4YbK+1o0I2KcNax0dMk/+EQiuP6NKs4zAClTFOMkJspu
dZYO1Lse9CVsIDLdPNrX6NkFu5pGb8jdq7Nz2EllUaCk6AeqGTmvSEJ82Ash3f1EVv906IeTkMvR
6ZfEkfiey4FcRoL/bcES62mV4feVmCQKg8qKjFd7IYWKu78C535EExUL7rnlM1Uxca82MMyH291Y
l+1HSZY2ejGis4EHuP98QRzE5vYm4J43AVoo18YAweEwXoyH+qTgwKMfTRDNAINqrT69yjFCd/Zf
LWlu3eL3XX0DKXCkuJVx2SJWawNfxrxj2LDI/6ZaEH3mSaTZwmo3Go2HsWFPi7T9+8Q3zE+RAm1i
Gy+LTKUzCqlbyoJqPHG9of0YhZTfyUv/VrbmcGIirsuSqyrkkOM7zWrgjxVvS1ecctubI32RzMgU
+z6dDrn9XEGOMZH2tAnHCINVlXplxiUyyjpfndP0/CtbHyhTFVKOBMzTfdWkg7QPjMtMF6lkBR1o
XYff1KaQrsLOviKoZ42YDFsnbVXF9xT62VYb/sq9bQM1RfGZ1A0IuEqg2qtD4yQWQKkjTQvScCBw
cTyLkI0T3+AahyCMC+2fCRonsg+5A0AsulcEPRS71g5EUOi4jHmoTjCzbBkTX3WqhAuJN1KLFr3H
C5U1RxfixQ2pDCxcFXTyB4M9vYI4ZfhA5+RJSHfK/5nBgfEVGevXUUYi4ZG0kofduNcOXEfzwF+W
HgxgrdMtA611rzQZyEcGahVZoO3OdG36eNi1s2IbeR25a/GnmQHneBczjN/ivO29gbzXSbckR/5G
ofpXA0DvcL3GCRJSeF4QiHtxiXyZywh2luB1GpyMYClEOMLF1FRTMeinQ8kXsx72TOSzNE6g6X5h
dxlnUCIq54QRvDusPhMZjX/923lMrWAfkmlPzabUd36+EEwD/um8ww/clKGApMWGzCVyoRSEqbkH
iKWiyIrfnbSMXs8JNpyiEko/pnO6bnyFbzpYhBX69BDmo+5t11qXEjwiMvTp5K4YyAXx7No4lc8O
UY3QJl6RPsU5YeR9rFjoPTKKOJFsCLZOOZrt0QsgGTyXXvRTQoQqSPeQDkCXUETFKcNAlFCSUrdW
4HrK0q6kR8x+Zx2L67mOXFne95Ir5d01xO8QIp9/aWaePzHSrrO3TkAP+VLZhrhhCWqd4YiD2f9V
SIMTieBe4I736HCysl7G17xQHqEQg5ayQgIsWBU48gEaL2l2mgb65qSVKp5oV92RvSb6lvVYnlq5
+6YPNUAXl3sFtZnpeNMDKiIOUPiHR06ix/3IXZcSL4d0ibImNYwe+/2uBoOWtpPqmi1KxD7ImXjd
VBjJme2H21OiaIVvvtguBqS8LErL1wzh/HcF3GKTcLSfy/hXp7ZBtmTlyyPHVQXisFZ0yBJdSamR
Ek/lOGLziC7dfqPJUImv4E02J+eFXipANpfGQcsc6LbPEZFgu+yEy1xdGyhaZB1ErxFcvpSsSzGX
OUzhCX4dWmUFky5oKotnbsUvpK+GloKM6ER98e/bNj+tbu2jXRJpN/4ZGLeVPYdaa4byKKIQUhFP
hqU0Bz8iQHPckSbbJiYD1LwK4iRBz3zRGxTWAx1cbPNIXFVGXNLq7fy3H6ytKdlEbcpR0DJUODyy
7Qt0wuBq5DB4OF/+kgZAcPaLerRrhZ6NM7s2eOtNC4guLKGly/FKlA9V9K1enz6seT4u88sXl1D1
cDAnuwrWNgBVoDRAMa6+EEcp/hfQ6XKTem3nAo8I1wQMsXeA09kZPchw7pkVD4eagWIze6nF5zm2
jpQwUbMWJ973ypgp66lW09fg6z1j29orh6T7pJJsN5EbKwEnQ7NprzC1UjzvmpMyhwP0D13k7QGA
r2VmNztbX8Int/P5rhzO5eaNU0qGRSp5VcskdO+Vy76gFonZOpw4VNu7ZhoRiDpX3Yjn3ZaMEFDP
gzPvvIYZBdjOjroU5tMmnXFHGHf20dLuqAx96Mqp+HLTB/7hsoPg6woL+emVDOzmHnFJH9ylW6hN
m0XLnKR1uQd3KgdebSWjZ73DIEJhMhXD8E8zaW1QqALVEuZSqNJgXCsjip2cyJiLTDeA9hSU1vxv
JgUpz8B7kzq4/HU+jAAhKt5heu4mYuRcy+SVtscap1CPDi4YWrSxZNTyrt0wwoz52u9uGqeE63GO
ZQsLilWBZb9nyOjzU6UZQk7tvd2nsCwEpH8SpyFkxMww5mxD0FZETaxQNiRHu807h+H1xVzdDEzd
Ya1HrZXvMSfTf4Hzoc8CYo6uLNW5w2Bu1wC1NRcQvZ28wCRXU7e+BwY/0ofQQvP4pd0Qd3dm/G4m
jagV8FB/id+YnIvtih2lRsdHQOcEnU3YOfKtgqGidn9eCSLmTbRXG6bmVYbqZdntDg1chY9BVg03
uo401sIP0hax5YOmbLovSPcLg0LGCJIxgFKCzAWw3RsgF9JEbhj4d1px4Vuj8IcwdY/pIz80+zg8
vNfjG6zKMbB3FS79TQIgBD1cowCiaKugGZRMSm5UyujjW0gQ0+ilB4QyFu+bfIb/krPUHo6tz/TD
AcAjfJxROhyXqQ1/VenMLqSxlXuNr3ytMhyrdUFzx0szibvWeB4erp7WGEufji/D4ogxiEdfN0RZ
33hKzH/IikzDu11D5lJ/Jc0gXcSBBWTsYbzQMyDsfX8iXUpxcw3i9Xax17J5+I0l0okCZrHqtwCP
Xv2WGiByas447ZjPhCx53ghWPZcpKOfsdUZQqUPvFhTU911UuJetM48zy/4Cm/dyDnFh/VILBWKG
h0RoV+tJOsVfq5ifUahXZaK/1gupyWz/kxp0+HtTOfBvg3N8JikUAz7xuH2cJHvpGVrzCOrpPy3x
SgW7aRajVxFc6XZJRQs3OuLEgskTAlKNl6b7ed8dHk/3m/I4l0Ir2TPH95P2WPC9C+6i2Mum2+Df
v9EEWqyTBHSfsJpid1uYguDn/PRGxGj3tpuGgRh5bWH+QZgYDDtlfOTXGC7TuNfsPjRwElrxumtV
+xmkOLTeXml3R4PjtxHwjRd8U8D5vlxhSOq0OJypaTe96UKb/pR7gh2d0KRUNCtNpt1aUHLalTI8
UqcV1MTmi7JD3yp/lGjey2Ohh6G9r2B3R8n78JVPXDvKmp8i9Oh/OfNH+Sn2Ebh6igOXTjU9yIYE
K+8S0OCxukH27xalQBFINdbM/kQdMbh/VVddybRJK+h+J6pvRSX6GMUeTHZM5jDvGyhqs0yPTk/r
2gZllP+BXH/ffkFFLwzLEPRfXbeZGtdjgD+rSw71jfqcTK/djn0RBP4ahoNy6kp9vjlMBSYFpbl9
/6UlfdE7vcep4n+r8DAkOC9ko3ggOkt2xrjYrOXMZ7P+aOx+NvwsMfeNte/n5P9PzHxkY0w4Ak92
3Bg1J7YYQNmwqiZqM4ycENoOol1ke/WodWKYwF6bt+AXdz76NurYgH/nvx4nHFpD8B8NSl12fVUa
ZMxGu82KrINKYh5gaFxOetXT44nq9zWyv/58lZE5zbkkLgTDEkpOCzdNji+IUDY9heEq0Ecnbj2/
kWDDwgP2WsNa1QhG0BYGX71ZcG2mCTg26CBLsrTl6pPo3qwpcgEXoiXaqFJoga6qk5GPkHopOIAO
6SRlyL8HpGtLAwuaUKRvpgI4S8POFJKadh2gs3RAgFT9bPirzYTlPKafYB2GIUnQ1qrMzS69gs0I
2rGXsrFJN8U0EscPCu33If9Vmy/LETAt5x7EzZxOUbjmc25KmkSbp1mluhDG0m/WALvPGIR2PeBK
HlkTMEG7M3IkUGBMMpS8evk3PVDxmko5YEl5O/lmdLC2v6fMZdp6biStmdY4NNB26lZk+3EVSX1m
uowMwQpSZDRsRSmaKQq7hSzscMdltUQo82+6ld5nE0OrdkqF3YJzbPwij7/hcC5++04vyRz0BH6N
cx5uvija0lNTgxmgv5elr78FHv/sQANYvjUzh+J1/ZD0H04NiQ0aqsTTlTjgIcXagmgiQT3Ybl8Q
rvXPXy+2tJBU8HKojwfrjEj8mUahObrqKRCSMOS/JoCRu9bYe81gSnZWLqMkS0xEADZk2B7z9Kna
yJCu2kEWNfpmqb8E/tiYDL+rC75zFKwoX0N9wPXYmwX2ysCHGuGBz6UNXYr63lTedAjqoh+ybnjs
K6/CRN2wf2EdCC75ODv23/oQBg9OJlyo5LLpbkpmLvR8t1ZVS/cgWtR/xlG4PElYQVah3qF4pH9S
7Pn3E2MzjT6+Ehw2RQQCWxnLipLi6Ebvv9Sq6w7erK3oxYrJfWymfuyypeb9oUaowyEVT5RIP3Fo
iUuIkQtBo5bnG+Clb1Zjc5vCfGlXEdm0mlDnh/1JZL8DX3qy4F70WU7pyoRPyMfKE2lXj4U37u9T
59yeyw6OdSxSVIY97cws0L5wsX+B1t1fOY9z3DlbMcJtssBk3ZD4yXgAEs4W8JJUuzFF5pPF3uS6
Hn7q0l7UsNu0LqVLNGtiW2Tyf+sTTrmPxdn8fgZLmTp7FOIYlqHIJu2WL2zuBdYR5x1dsjO3Hg6o
dvmMstoQl6Fnu5vRiFUJ6njJC5Pj0qHpYUdlKc9aAYrXdpbUWw1DjFqKuUgTbBPzGLg7/mZMTAFV
lAWIGaeu6GmxaOHi6OyNFTv8JSvJ+xJswp+Z953Z6vkIbMTpBJ/gHF9ByEYAFnoL8J8ML27RrsDj
ojWt8Z/b9vUenWeVEoJG+eh/QqMh2CwPk683GuH34OiPlphA4dQVxZjnj8vLew75q0ahwH8WfXWi
HdfKaVzuq3AjKut9xP8dn7qKvlVmWqa2xYsG2p4fSQ2uL6Uw9G3jxjQ1uOPT9oTWn6G3R1ridsfk
y4RG7cwroDn/lJBj2n5ooNF4HmpP6SaL4UwuXUM8l8YXziTEb0Z8XbhRCM5PF15uEMlne6dL0KBp
PNgcnlkHMmORGU4aUzJShlkMYKC2wSqXtYVYuPyRJokIauwfJb/hiNN+qtnqxoQHIeyOS+vHUL7y
JsK4R056oEtaoU1QSsyUXd8h70h1lM51rxC1OMwbR3m69qfzHg4mmLOY+8eUd4BEMSq1tl16bxMi
873ug0M5VO036UIWWZKPseq7qcFBRMWLeRU8BfiL4OzciZj7V5hwB3zrspftOGTby1gYw9m1c+rM
mucFzibXj9KK6CXUKa74jr+vVf+SResF6hLptbDowPve0EzKFL4yfO4EY45bHMHebavxmWHGr5In
Glxw7h5yE3QpvoqAWkTCjF5f28kQhgJ2d5ESFcwgvUGQd+rylWkpg6dMqviFysmJJhc17w2PdCuc
ZyfQns++CGrHnYJK8Lzw11jSOxcfXdFhUHm2yO+IfR332p68nno/sOy/iDy/sFCWV+Itj/I427Ax
eqicFkfR6Udn+jnK5DatmpyVFs6Cwm/nVVtLo+KO37U49b7tVjiyphWuUiv6SJ9XKdZy/UciNBeV
o0JgzQkI5xkk8JQjXaKexenvRxS/4/nI1W4veNbnqkrBiLh4LxutuwwcJdE4zozo2NDpGz6j/1FC
jLY8kTUkzlBFiJfkAJg9Bl4Am5cQf/wjWOCOs6FmQoy74M7ZvLWGhqZ+74P8DXjYqQeORcvdVD4l
GVRVLhajrG99ACdn0QJM+pThTpygCUczGIDdaSU1GuTlFVtjFchCegOWM9yKGk3Xwp8SjGUwC8bq
ffR4HgyAO3ewVpzYAUtAmtRDMHl2pC1NPq6N9pHmsaTKpXeC3F+ABbL2oJ9+Y4zCp3HtLWAm3NE1
IU4uPuAaibc7r+5W9p6fjpg4MkrCpasmSqYzd6FFjK8E1y3lmFEtUuVwbVNveoj+viErt0xLuQYN
+UuBYSqoDjVzhH8y0Umpg3OZijMQVPZP8ObOeGsAQl+hrhe34WZtxAZ61FZFDvi/hfQ0PIMIJ4UR
uUex3StRk9+Wd18JrY8wOe1AXXWgIzxaRAIJU4Ut0RR88tS6uf3fzO0aDWMS0s9K1WBcENCjC4mR
aQBwtIpjT5f/ARaJgHpY/IBfK0uOSugtXhZNO/fZXzE5GfBeCEWUhYZkK2z+ehUHU6JISxkkjXoK
n8uKHFwkmHoPaqPZ0ao876U+/i+3yZH697F07+xDvWwGJjqNP8vJeVTuFxzGB+PwpHo0ict8VGjA
dotQqzSmgQZ+1awmcH8Gh0zS6Ktpba3fRYNmXuCZK+HWm3xfPn9wI/gjHQyk9nq2VCzkrxignYSs
3q2OeI9D66NUHL/5d2DcOO4VLybHNGGJJHCRvZDMscT0+j/LOO62Bnm8nm8ISGRbJFlXHP8vTAeF
neKhpjVey7ByzjCrw+wOPbMayLEUI+X+v0HhcP3AoBBAzvAVYU4GKn/BxZ6DE8w9Lgt8pleSLKCd
EPUQSiHoiwRXbr4KAYuxDU+IcLxoXlo2b4jCXbTFLB9RDZ3QC+2Sph4Ni4gbnYxSWuU3Q3Gm0MbF
sk4+XwkXakGOb6ob2vjiTVujANqkC5/iF+iEVoFEnzG6HM8Bttq6eYG8zmMaB7X7IgOawMK/TA49
hUHWFQ9yhlS2CaRBLdn2T28f2cmTSVtaZ+d5yKauoKpIfDegk/iyIPHb0G27O2gBIYUjfeAIxEsH
z/IYiy/pVIrIkndeqD74p/mJbAY0RDr7HkYLnAywERz4SJ/tLShsQ/scQGy4omunK3Gg/+HstSHw
WklS0jbnLYFG4PsBEXkElZeLMSeXlS3ACrOTkEnG5b0xJE68L75QVmYHgC3XC+VM2SvvfUCyqCLT
A9ySWjqzKzmg6DC+v8CwgrZDshkpE3Lu4/L9px1LxvzV1IbIcP9J6oiTyhOLPkPU3Abbwj/kAQG6
5LGQe9RjyUg7vvQUr/V/7Nz2WBIZ3ptPaGL+9u3qPMA6sTJwPlm9Sd+MxYjrzDHsYTsAZnUHaMRF
8WbPoKqr4eRGw4sALTMAPgePc1udFCk0W/vkZ0PCozjRy1SXmz9eS8jXKhgzgy5CwxeaUHk2tl4h
hBkbfGOZT48NmUKZ+lG7Neg24REuCxOH31M/ggaSOi5DyjjhT42Pt4DDtrYxh1kN+jDGyl30TJ26
YRQh4+fYPL2dtkQAIR/qDbVsTYiGY8Lz3AJrlUKsyIb3F1mj9Y9dbn6pAUDqXBnKba4SHaUwrCPS
CY0C4qgQwMEKqeza2CtaFSy79MqUsC0gyQzzqqks4yqvgyDqeWwpA6ZX3BNhADl5Z2TI7mk7U03R
qxceeKwOpI99OPkniYO1wsboNI4IZtnwDSOaAotBHSZGFs6ASztpMcPOBhVHXiLcNyHnwl70o+o5
pccoepd6v63obrZDTYw82xL3IQGoSZ7CsAl2g+65434U9JvBrJHuN12anQJZyjq/3hps4P0qOilZ
BM0Q0Da0MTQs4UPPhhJPl/43YfNhKl7eNWim8CSI/6nrrVJx6nttC0wf4CcpKTSHU7Bffzl+fMzU
hlvRifVl0vineDxCqs1Lmf4ImpwxRVKgekSE1Aj7hFDPtqJDKlZd9hZaHiARw4joyXsQVlrlT9GS
kHBszNNqtfDbt+w/N6oKyKsj2JvCW9uF/p+DlZqkX9lQCMIgaFLPSxt6OU1oJ18LIpUGkJQpuQah
PCblhDHDqn6IB+DtDo1eUucM+TpHH/XULvLB6heUqgbsNc4H0nkiWsF6MOGf3kpZw4OcdEcAQS33
gcqRK+rUlh+/yZzJTdoE3mC033VY1tnPm7tvFAfLVEp7AZVT/R6rGvVnsl+47T274XBLFLly1TbY
L19rIo8PmHWqMbOoGenUYrHNgeh06TlidaprsFugw2iLEkWx9Py1AaG5TPfikxo44f+Tt/UZFlfW
FoJsYKHnloWxoJU0/fSyNQNWFQGmArWaKHHGgQToM5mZgrScIkpzfDerrf70UamtYyXM3JHDQQ3M
rQGbzlq3PcOh3nfjPsLE8tGrV/5/BkL39LSQXkP1n05nVcqFPNCLIjOiA4fOzHzTFdvvKOazZsr2
NOLRoqAoy7V2weF35XQ3UBmnKbBZuJ+jirra/Uu2sCprmvlxDE2jj/o514fjUiGMmlfbLhGcijAB
fOmG/qUk4o0T/cFi1/83E/mXASHmBRVjwUhevNnO10E9uMLgWjApRvAgw1rm7jQVFjglha6meWtF
0srsKYhuOPHJVzOuBK4EH3z3YAiTKzcuUyExOQapytJCnXjTJKmAVzSwi0lcMWghNRD44QDR+brb
oqAwB9GPBAoZAgkYYfwnRvZ1lBNvvPXFYZdKmuBhfylQANQctY1qfPe4+uSMWYz4Kdb1r8nLU3GE
4eyUbRcHI5ZBLLtAWSANuaiPSvMLZMHzvYzwqt3FWWzlpAF2GUBbiXKHG6RvOMey71S7kSSqoOhD
+4tFsTEaiIpAcLghi9HvAd43ZwMQpWHhsAdz3oikibD8AwuyxeVPqjt/5DNa77CBwZO5sd7zqQCs
lsa3a1QY+t5nj4nLCNUak688t4Y/O9RM9TS49oQ7lNu6yj3LNAyKlHBlwf4aynFdxT1ynmBFBIbe
NL8jFVX2F5l3pRzZXWslBcVm4xzgGI8J4Xz0KJg7R4dXKqyb1zHAOnpgIAcLYf2zouu+fgWUUtd9
V9QlOeeBN0mWJNzcoVWioFStOvwQ9BBajS7Up+BSzHRAwC9zLpjehPynAPZHEYjOOVK3Z/PAnQAv
IHpHg3ZrQa1D51MX5ss+LhLKdA1T8gym3Gk/jy6SZqgWJ7n/6uB89QSWtRZCCeQfmxOnM4Q18mp2
XpAzKp4IyK5HwyEYKSGMZ6suGcQ7YFLJqbMdqsHvAQuvXo8ReU9ygzdLCsjL9YY3FlYSyYanhcwR
QLzGIc+Ecvcpy68L8tZLOMW5ajynDnsfHHjwMy8y3TBUngO50n4lPesXntFU+8TPZOINNlfJZGsd
XuoaET0AyhTmAAYPTowwFqgsGKY26XEwmvwYzg/TK88GT3K2KlRhrHa9aNkNWur6s0/yjagKOmLE
QXo6k6c5oivo7rgZ4kb89ahhaRx7vMO5OO98GJ6nL3iKSBdAkrA8/3s8zU6bqM8dArHdaQ4YgPM+
dFO2XkSRrz6FT3bmlaBVxfx0+4xGVus3Y76PzoPIP9TDicWCdDXyJ9AQT95n+8G4RPWAfPfpumnP
OGdCOzVBqQLvnmyQVCa7z93lUowwZeEIr0IxDw00xn/zbVcyFTe1Mlhu8TTqj/qoPgMhrwPo3O7T
iVWegt5O9ETSnYn8MvYWDbcnMRmCWRCoCbza09OtWtK8B4WQM43AEQQhJkeg+j0RZa6DaQiA8nFQ
KnkM+AT0GCj46w+OcSflXYB5zgZx7w4gHOr0Vruirz9dnktFd+XBCEVxnMHeeZ/fLzrDgfyJJZ+y
DN6O/I5m3yyzff3SmXnp4VA6mDyGEU0Kf01HoO7xyTsQxeoY2c39y39sigj8hq5/HkLlB3FHi4Fa
Kqdbk19+2lEry6xZgrHtg0kM+OaPCUUSG0GrYs767RPutrB/wfYTqOhvlH8foAPYVS+J+IFO3sfZ
3bBYmOVlYM4jNwpowIrxNHK1PSOvhZFnxy/vcQ8SNgr83EXhEw8ndCit+Qr2An3JBFdIpK9k6Tk2
mQGdk7tzKrYRfPGqy3AYvkqnPkS2XwzHKZpfsTJ+e0fyTFbIsVXpD3IvJuDkx5CZP0/1HGxJZNR3
mPRqLD0Hnj5EA7mET4KjUXBmYbHhfyBdtKVqk/9yhSKm0dxWcN04UjQy/f3Wlv38VzliN/Nntwue
dWTvgxMirEJqYj2j4KUFFdvCJClhZU/4FcU46wTL0HSlQ33RZOYS4r+ua3m8gGXu5Y+T3/XJg6qP
s4LjmMC+xF1kVRVJiJrMintjySvlpnYBfLDVxGlHbCCswlsl9Z34DlstWzORzlQO5FoQOWQEfVS8
gmZh6Dka/PgTFDLesQhoHXQQh6EN8oUO6/ONhad2xbMQDXy8l4PGp77GfpfRRvc8x1vXWYM3mIUg
1vT92q/DGtKg6GVBjuaLQFTveeYMDTKScRMLAF1VE0A/X/4LZvWV/Pcq/iAR29eeYXX9BB0ek4FI
rHk6uqHf7N3JLeDOSvP624Ur6te7eLlYjn0n7DOFSyrNo2gKWgzwsY7FqDj5/3okg9ISXTF++B7I
2SszqYrJBdUHL6K+UUmGOjja9o3zELAMi+wFE7mcuby+D7X1s9eIkIVrVn7YeQYmS/eIgzjeDwqL
RK2ylnkBwCLtT4uzz2BRq7d3xyefYmtuFkMObKRVuXomoHyo/hbaK/5HNRi1eg/H7E/OEXGxGdbE
jgrSOC1XxhYA0dC6o0ndkstx9hDqUNVY0LoeK2s0fKjXcQkBsVnu1kZ3lbxIRSOgVWx/ievBYFnl
M38XXt8adaJ5u2LL9OL0rWoJonlf7jHghb0LgYeN9L6/5x9JPvk6+eK1fbyqbRkiVUIb69bl/z34
Yle/MRb3j/qT2c6N9CHBqhbOsFjSV5R5Df+VhnY4YzYT9Vl6RQyNbOOFnAsR3fNSWue2FNT29WUI
ZYD8ZfjJU3MUiHC3dbvv93fjQfmpVhr9OpQZBix8jJr8cGLHyetThlDGhioij+JxJUKGKno3xvEc
YTKB5Ytlp4mDaa0+HZ3So9yL9XJa8pejp2ktkGZly1eYVWRmK9fsb0Y5wcxgOXov8cbPTy5i5T//
bFcxi8R+qk/Gi0johbN3Q/RyVF1s0s5k6WsHf+E6TWtPileK/cPDFnzSs+8S8YjHT3n7LNWmW2eX
oVUaOQM3HnrEIrQ+7vqJT7aJ/8sVLNDvBlC8XmvrU0ZQUUmKsiJJQTRxet8hpz0re2jWYdeDFi5t
n+2CZmP+fUKKpXWzBFsXdXbB+76WP08vbk6JGVi1XGatadAcGne+KHV4BD+rzD8PDxBK8sqUtTZ1
v3t3sdQzGtnz5SmSjb5woA96ixJgrjRJlbWBiho3mqQ0IdRktLYNgsBank2GrkC9isGuGCw8DufG
IPjn3YWiwnL63n3rZtKBbYZrJpb1YTGp7cGPea+iI95cef0IBKihAOO50bWQjbmSmxOJB3xKnRZI
I5ZF0GXklOmIdkbsx8mnRBOng6Ps92FM2FVjdLtC+nyMjc29HFkawTvsE0oZoFxHmxKYnz6tixY+
I7g/lNdgKlusUXBdHumInuKnUqE6NyqGwAFT+1s63QN2zPVB4M0E160Zzy/IYet8TMXbr4UnaDPS
7+fLi6YmPy9lSYCCgKbMmN06xNX5Z2nE6nztMc0DQXO2yAiFjkvMSXyinAOHYIIkvfps2vTnxnEs
916o+HyuGJrfES67FFMo2C5jZq9KdC18tg9WKkD8WD9fM0CF3Fht696D1P9TraIc7PlavL4K6OcQ
PF/52HWJS2sDghNf9e402ZdXuAUyOibgbbaymVSfCrzCwP/iO1OyK9mCSeppcCpLev7VrU7Py4By
ANO29RP/7njuDMFLAxVyseJNpDOlls5u/xPX0AjVMP98arkPSwpnFyM2zSncJ9KMuZreNW2nhIVz
8GHOdIGlPY34OY+b8PgMAOo/Nn1wEFBzBFB8/iOgFm+EWlAvdVjAyu0muwIvpmm6mAy8bwxByYVm
bBGdnL60M7I6coTJgjUA4GMapjj6Zzz52/jJCDDVPVW979LexM/FAwt3QxRFrrxejKIw4VOFMXPu
8V3onkB130wBsUF/Eg73Wz4+R6QCwWcAk4dEPx80VE67HTcxfkffDSUoZIE+sLOXLgYaB6U0NEA6
2R5cfXBwFT/QuKvXqsjbJTfoVf69rKVJfKAagksJyJRnlUvo5l0PtPsvAGoB0/2rMVgrv3dtdc1z
38+Mz5niCI/KPlc3imOjIROSBVrCDrrevHHcm+iwViNFc6wqKJV1+A5FmLmpizIphAIFno4C9I6A
F0+dDevn22SI3y/59nw2oPCegB9ULZHbrZkWh4iMKumSKrHdaNZa8MojZdk4a5SpsTewnWKZYMYL
EqbXwMU73B90IdxKYebV+Q5TbKM27KJBCLFnGnc5iCSSaajT89pwG9lEsVmypo8o3/aU6unFr4Kv
zeZrP/36+8E0iJa+i2TpNgrbs19wzsEnDUhYwgHj0HYz1/TBNWCbUtFliqjm76yS5M2y2/01+EYh
k06TqWiCDUUVbuG0uGDouix+Ia9HqtFdwwGn6iCvG1M7+obhmDr7GweMujwAM9kzZ7194MufR6mg
H9fJHKTUhoNAOf0FQXtiJ6lGFs8e2qk3Y5f4EIUQXHVnZF+kVOTUAzFHCLgLR2wXgk6cmwwntIRh
isBXgzsjLsyQGpQhoGKwPY1ZRLaROS5dzjNigP4mWLtVbyTtygwR5+dieku/0FpULa5JqDwhhDcT
TF5TgU4OpjjDi8tKDTg6lhZ/XHNok4ijBddnXhRF0yPMWskF7zf5A4Ca7l/7V65tpwyIa/cIzLEU
WsskbMYFyiB5BEf4v9jO0S5PYamymaRPbgAwfTZ7Aai/zB24bO/grBB6tH8JvyOTSsbj5Pp/pQ9m
R4AXCSY2rbW6dt3f/DcdvpHn8TZYhICrtIm+mloUjNqb7TeIZqdTMjOntuObzb4mtR89lr6OKuGI
bXs3kX+018bludCUZM0GnYtZsPy9HfzlDdchKp/wWqPlFiL+ieS3yiJf9hM6G/OOdxFaB7BdJKbb
C0NtUXO/xp33it9G7HyiGouA9rQ9AhLLN3rH6HcE6qy7866pUzcNvE7sAswXd3Mqrl/simEnSvnB
LEYLQtcYacbpJx/7CJfrC0BXbORrjMpuernMeM6qYQekaaFfHPHoI47f7oPrdNiXewiYakvmyJtL
Bgtgy58O+c/Ec4CEJczUo9DyWrCjULgDByWLiIjkTmTRWLBbDhmYzlZSOcsbwIOB/vNTUvCbvJbm
PloLdcW9xf70T4AvED+glnh9FTPWIWz1/EKGArFJ91UTlsSPKgvzFRasJQqr/AQC3FSnlPeXBJz2
MQxOQDkJGXQc9lOeJ35C75l1EAF0Ee1/02Kn3EqWDiRqUnoOBd+J34F5Q0ZYg819wf+dw/Viq+cj
blvQ1rUdUfABxiTp7B96hPiJHHpRGw67AzZF5Z2diUKGF7jifPDYmeiEdchsCRUBz+KDdNtDQ+dU
Je7XQK5aPQuyd1TRiiqeKW57Nl4SNRsFSQjsM5xKbxYW7kSfXJHqebEh9zTcrjNAdChqa1KqEp/8
R1BF9LS73M+6ANCvLi74nhglN8kvxGjYpFCk1KGCoDqoLdIer57lp4MJLm+UEHfYvtIQ7Hubo0u3
Ozlzy7t4cHJ76vriIj7CqTZk1eHNk3imewkbvHDNTEXAwyOXVaOGowUkzLGtBM0wCo6eKrMmvlEw
/iyGDbtS4PxWmosAQijjz0uJDuWpVqYgCejdiByIjbmwu9vcfpkhgWIz3B/IlnbbQC11r8NjIYDG
6pqYwcv642LiBVGqLbbYBi2PKClLxB3QEMb4njrTqin7tEofYaR9xQdDVg9lCbIp0Ns+tnabP6zU
rYqPWv8ZsnPMErhjpOvDM5o1v7kyph+w5iMwcbVb3UEvjuummlcp/IhXBtnUgv2HOWcS32vlHVvz
EkXjAqaZoFWwVQW5JpO903DlAgzcTye1HgfGqw29V4xKft4iUudO4dtdG6pmTgzAJZpFgEofJbds
elGauP01yU/amFYYV2f1QXG/K00Y5OzHrJ1CpMxi91KOHPhoKPbapvdL0vvrjEJJpiPU2BuWzgLO
CSJm1gc+k2B2qcMFOkWGw0pSF7W9E/VLG0xDvsb0QfIAY60nWXafllWZu7TrlwrVW+htMWMSwtzy
ERB6z8iKx5zgXbOKb1a2ut92zlVNI5xejgFuIvSUlZX2UMW+e5dUYCaksHra2dImcvAl+fjORRRl
Bu831zR6iJNkEygB/Oh3Esq/j2GYOSWrmu3hUwUGY3YujZ8n1cSbLKR38BSeN+Owk6dhhp0fdS3L
4fTuXocUn34/NyRipmkYyUKahoQbAhDy/XOydL3tqGNMxshvRvZ4aqxcA99orlrHA7tc2kka700z
4XxeZm3jd23yHaU+ZkP8uAxN9GNlWoeEFCWxaRH68FJOCxe64zb6LbO5aUBcrE2lzey461vhKE7J
ljoukeWir9jbKl7+B5+zjgYPaB7kRiPfQZ6bGdL+MWdeacxxnTPUPgkFKXh795dl9YRb69RkO53y
IB2ds9J7fU71+/5FNboXa2Y7LcHHNdRzkzOB4Hd3Kvo9zN4tlLpQGPVMShKVVBJv6amGu9e7+Kfc
Hw9jfPSrvuHfejM54ggfV3+wvKMDdwfW7GxEQWga+ilPaLPFEQHorFdfMd571I4elbJbZp4+gWrw
b4i9S7wRbedfqnh3b0TX7LM6NWib0xKad9n6J9Pq8vEOlpQlgnO9be0NPgmbitBRdBxBqLW45vgD
OZC7B/KZAwi3D61YaGANsGiJz2jukPg7r+aViYDSNRMsjktgY7RSIeX2S+/DSRlw7M8QKy2NIvT/
jMvltPNXK+x1ADPPIVMhYRyAVonu7xJ2hoMMSiNOQnZiqyO+m+/eyLdsra34ac03Z5+PV/ToTUYb
q7C6l5yGD2v/3X7xYSNldOBrB1jOUMplo9ny+MUbob/jd6UknavJH81EqdN+BuJcgs6VP2wsigEr
ERJ5cR3p1j/uTUEAWsSv/pGd8NgSdLbfe45L5J+nvzvF20WJh1sN0fNVVgdxkDq/AQXEwEBnKymD
DpPlxULjiKMn2z3U+M7lSEYcCsJTEtd9+ByOM1Nv4eabG91tVP6H8+vYLRq/7UIc9q84OFf3T8OY
VP71NUz9jdfN/Rvg2SMIfZeROejtfb4f4IdX9IAdmsIj/1gKuNiNak+ica4dgFIkXkV7imXUqh2R
vv/DSi/l6PybLKGh0gfF/hDT1UXa8RDaM5sJgNgeL8qPaNWptZ4gjTfgN5iDewoBjSTlnVONCTHu
QFGeVrnd5ajbESfb0TeAG1xyUwfrsZpt64m+SHLlVyzCPruNELCmakjlaXXqD+OM++/SS2HBZf6M
0po0AlyFOi3u8bGVLfzAVoB7+IT9Pp9a3y+c9bm2IEyecuozd9PQv6KWgZL7p5OMX6M7wB+oc7Z+
XlLgsxSOiI8vPmzmYtY+VP1FTAu4d9P/NeWA1TohQ4uFOFjMUbfxej7lkucck/AsD2OdjpbZeqtB
ILSck5r3CVCyP/PmWiYPSWfqbZFFYkp/c9am7JQKEu/o//w7qtnc1pXdx2O90VmRlsxzaTkWyf/s
78jl79T+IE64YcK+HsGWtaV5wU+4sRUc9l1swXexBdlBGbxHjBTJQCRSg5FiF5+Q7iV6HflhPX+O
EXl09k0Uu8BDfmMQ19iJk1Ftv9Q/WfuxPiZybzo7sVHX+tZe/uLnsThQ7UW5KyaPUTd0PINWmj7T
QYRrRLl7oztSO8fAujTB4QA7JWanAyuWlM9K5JeE92dBwNAKb3sXjPcI9QOBKxVQIQXtbdzEELrB
dlL90/hN+xf68P7olMcK3tpwxFBJFQoWFNhIl2PQcBHXjn4RD9J3v8Bh7twkT47mq75uvEE8H/zC
3gqscYtF+uOSFH3EBskynlXjcB+scGB+6dUWnAGMAZTd1I7nUe1fKLBeq4O1lEeccB5NFMIX+qDA
F45UZbXskTsbudyJ4uvBLUPiHuuSklUU1JsqwB1mXBauoo1XESVR9zCkUYmiLeDTWi4S5vvLsAQV
MB44vM9ZeQn/WRjKkWFJIQ==
`protect end_protected

