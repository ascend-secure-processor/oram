
`timescale 1ps/100fs

//==============================================================================
//	Section:	Includes
//==============================================================================
`include "Const.vh"
//==============================================================================

module TinyAESTopTestbench;

	localparam RESET_PERIOD = 200000; //in pSec  
	parameter CLKIN_PERIOD          = 5000;

	//**************************************************************************//
	// Wire Declarations
	//**************************************************************************//

	reg                                sys_rst_n;
	wire                               sys_rst;


	reg								sys_clk_i;
	wire                               sys_clk_p;
	wire                               sys_clk_n;

	//**************************************************************************//
	// Reset Generation
	//**************************************************************************//
	initial begin
	sys_rst_n = 1'b0;
	#RESET_PERIOD
	  sys_rst_n = 1'b1;
	end

	assign sys_rst = ~sys_rst_n;

	//**************************************************************************//
	// Clock Generation
	//**************************************************************************//

	initial
	sys_clk_i = 1'b0;
	always
	sys_clk_i = #(CLKIN_PERIOD/2.0) ~sys_clk_i;

	assign sys_clk_p = sys_clk_i;
	assign sys_clk_n = ~sys_clk_i;

	wire uart_txd;
	reg uart_rxd = 0;
	
	always @(posedge sys_clk_p) uart_rxd <= ~uart_rxd;
	
	//--------------------------------------------------------------------------
	//	CUT
	//--------------------------------------------------------------------------

	tiny_aes_vc707 CUT(		.sys_clk_p(				sys_clk_p),
							.sys_clk_n(				sys_clk_n),

							.sys_rst(				sys_rst),

							.uart_txd(				uart_txd),
							.uart_rxd(				uart_rxd));

	//--------------------------------------------------------------------------
endmodule
//--------------------------------------------------------------------------
