			
	parameter			StashDWidth =			128,
						StashCapacity =			100 // isn't restricted to be > path length
