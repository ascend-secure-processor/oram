

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p26Qkcl02DOR7cnF7rHCRVPjFdC7HaB9rwK4z8ZDgdqD+EBmIHjmszweIYBYopgfBX+o8PxCld8I
iUuHA1TMBw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BeG+ru1mEHFr0NIKY6hnAx/dh0OLktcuMhmziMJ2KDS16OWv2Mh1zZwldqN1Wap+jJfQw33GfHbS
XABG43+9CrdkmSel5iYvX1tV2xN8ztxgX0niM9PgyeTiqxsN00SI/EAhrw9QU8/AGmUF7msmDiye
Z/9oNRI1FwbSe+WY54Q=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lC/xzfBqJ3u97mkCbZyYuArFlvFE1v1BqN5C9UIuFtyZsz6zuwLD7ZtEfK0m5IHlr8/gejnC+njS
8YSns7L9/CskvdaGgdu8yh5L1MDrXNjj3QZ7+QXm+m4kDl+or7SJgEOGIHHqyC8VGfkbbMwZUSVz
z2aafjmuhGH0AKwOvJGWpKTyul84bu5i1p5I390R64Jp6uJhGehMSZ6V7Ien8rIO5dep26ftUUmD
g5D6arfdAVJY+US87+5RLqbIu7sowowj2h7HZOsKKfP4lygu1yKcBA8kQWlT69ni/iVuZk3Mk2mD
3wBhkKLpKwXh6+YzcJtMz9vHwaJ6amZrgF9t4g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cUNB6NBOqkU4rdOY3oHIejxB9RVu4/erq13pNOxw9+DPYrz2fy6+ixE1SZhI+WeNEczhylkPKDs5
//EcKLWs+FRUZvHBprDwbY4XSfpHW8ohb8FVoAbRg1Cwm1v2tgp9vscGefiQkw7w0b8jK3VJaUjh
RUFPilS76wZxLGiRNSI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hoHf3Rf98TPxZvwGeZxCG57b8bRSGi4JUlqCWjUNJ42Qq/feV8p4tRxZzi8YblNTkv+XUxo6rsd5
SYEXp6Nq+9RixCiWOBkuWdLdKO+qTHtHooQ7XR3g3JWRHvMKqFk++pysEeuGNXFZrNNN3+xs+aMD
yWN56FLkPufakUP3HI8gLdFThgmN5113hv9/yjDq3QWTtQqv/udKlWVdHnLD6kKw77BoYhhxttoY
k5tcDWMbM/ZdInENwVRYM0P4CbV1vv/jngLRQl5QXbwwgDzh1cCcUdSU6roEb8TM35vDx7UUsf3z
3r9Kk8e6V+TVk7mjfjZBgwwh3/vz3GMA51UUdA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
LzjGss4AvQ4aFfHkWnAsYBE9fkWo2UB3TsGDLIzRIAPOhgkso1843I5riQQqPe9oMv13oeaVFmPb
UC+XjAqlUq4vblfYltW9239uO6wzVhw129d0MvPNcZiWrBB8XqFsNWmeL5xCVfW5h+oy77LwARF+
27Mpg3cLQYl+mwC2TVL8R6sSoA+AHSx1k7U/jV7P0OlYdEeERqmBzRbW9wNEJQSpVC4INF6MSlW/
L6RDutFBxO65p7afu+5nxHJM6Iq/gyyHU300v4CnAlLQM6CQ0W12ktrIDazJEmOK2eEVL/Vofu4T
u+eWgolTSHAjdYmoYGysOI6V+mQnJ+sCfLcd1MLjccE7iXiKkf4D8KJhEjBQkEZlXdAxK+XY4UMi
HlVTLRSf+Czw+RpqtGj50H0VhZtks94pRI3Y0xgzBUJyzEI6tv415MPxE+hxON2/TvDhsXfa//WQ
x+tWMFezDjSAKRtPNzbhU/Q/Ei/OI26+GlQYQJSMkFguFbMIgM0l9QyDhJUtFzDlqTb5rvPINbrw
ligDGE3RF/Slt2Iy4KEio13GQ4hfiEZHVxJ95CGpQilrcSRBSJE8QdBzv0i4/FEoHi22XFzo3ODO
bu0227zYjyTNw5iQWuvSROB4E73gMhOVVfEzFE8qG0cEJfbUm0um/ev+27E5Xdjcv69GHHH8lvNS
NlrCm2DiwcE3S5/eT75CvQccZgGN1qtRoW/nOFYw0ipHM+bTrFUlAK4OgbDfc4F9Wagre9zaz+zX
nBqXqMxX4JG3sAtOPp55FMw0rUaSfHZoYANlYdEyafGV4g9FfJafpKMjjY33Fzlk+DUCgqr1Dyad
toGGtvmMQCGsAEOKsyjI4naLJDgK/z4zfHZL9ZhkFBtB3uLSWuho1w3tUnLJOrctATX94FyL4Jfk
UTXE2neRzcbrSrQR5ueuOS5q0k/w8P8BnyuXBZC1MNa+QkKYDv2oYCASiIrGGUeqYoif5KIZPA1l
nkXu2Eo7/BHN24houXT1OYhxFyvbbjxVxGK0BtprD6l1eX8PPm2O+vf0KnM2QJ1ohvu0XXR7jc3z
qrW1PuzET2HJCpvXYQHxasLTQKXdy3vSry5odDlXGRTqIa8fmJ/SSxk/VhoccrP5d6S1EM1c2Sch
fsM+kokPuImw8Ox/rSXpZtknzmSvJ3jp21PH1eZK0oLH3WgOwSh25jdKlfhBr7M9uN/nj2ws1YuC
1SmW3d6qWiv9+XeyJd6mEOzgD/lF7pQjKMu6wdsk1La9XctLrx5qlAr7i0prDTvRVPQXixFARse1
xSbn0unQNZ38IszVcqk+HUyAQKUWxoPH3TH9KN/K1zZ/FCK7JW2X6Cgi5qeYyVMlJBqJ7Q+dfAiH
HnLiAEa82B2aOSuBd3PLEHk1AX9PUTu+ffHOkMXWaIXsRKCFR4jcCwNJwG1wysvEsLDaKWsZI/vd
nimpBxHr3v8gicesXZDMRqVKd9UsM2Xfbn+Ti0w3K5suRHhqrpES4fH9vxg2faSBg0uwBb83PtQv
cV1A90FeLnrRYxyY1/bnTBlF2F3Hq7MOu/ZSIqoxsya372nEJOJDA76a4hvh4jA01Li7CmzOw6Hk
ozl6JDz2DQ4MCFDRdswM616LHWxPZzeFh36W8NPW89xldcCWQKjsBn9UGtfdXdaNH5mJaiGUSoyq
z+EYCWMxZjYuRE7YyFPrVo2brn3HXApqbZUhPV8qC3TWcjeQTZYZFzZs3H3u3oLH5aBCuPYWK8OM
Vv28xuWx4yiXNdk2RuUTHySXZpVoXtZ1SeDyqelt+exw6JD+EsKSQD5s2OSDjtjgt2SGay571SjL
3saoVUo3yLGZPPPPIYW4pZuqngruNQLbLhvgXT/QwnmPNEeXAxjKiwCW1+XAezcxoawobMd4ckB+
RepswLfx1bujEQJ1UT7npfuYJ2YalIFwQo5HIzPVhlAsX4LbWHgYSXpPL9DauUGg42AyEWxDK3iL
IstfEvkqN33kN/7/7FaIZMMD6W+cUbpQ61Q23EFMFSIT8P6uqvkbaIwnAt7XGGdMBY4sf6f87WNE
htg6o7wvXV7p1BxpdhUbeLFcK6gm/jvPH8pZ4B8MLiUnxLcuvbsRrdbcJlsxSTjOdSnnDZUXMHVc
Ez0fhuYQjJuHKn50o7Sk1ELASiyPxjXhbzTf2uqYZRq3xBOIKppMJCvfP9lK8cxb7XixfBgGaXc2
YtlDv0QOc33CBUClQyU9XLMMPzpqpUrG3nMJk3lYhSbfOVpIAI4Ihj1zN8xmdz74bxdKw0d4ZbGX
s2PH1NACqNK7jQWgl1+lwOONFJzScxkl2CtFGeunkRaLXS657EEB+e/1jQij5VOGsiuZ2BlacDek
CQLgFWgRevAAHo1QUskuRwe6uxgWGk1Fv+Z8VMZM89py1AEapt+QH+F2pzYkOdxSQIZpwvjl539f
/sq48x7RLA6q57O9/gr9t8wq9QLW9q90iCMVJhAn7XVeiHB5KMHQSPmYWJohcug5U7cI+W4SGS1L
Fv/s3KAA58MZ/G8iKCbNf7Z3mxGQyy/S0ZvZzvIsJC8RwShbSV7LiJ1rSovrmXLdonWLembcK7wH
mBrjFHpse19pLf2CbrHbMOw3pFOf1hQb/jErUAGuyasm1wK/wkkmBT+QdKZCLR2tvf9Hi61c7MTI
Z1MSybEO+5vmV3y2Jj+O7nwKBnQArIkwG+0scoB/4u+LVarvdmFKX1VTRIR9U3CsBqCmbMKt9Wl7
qNDgGBcJvzHdyZij+BzxwqGHOQZ9RKT4DcuoV6ta9Kod8lEGKzMaHHIPinQ8zwJxdUsdCJmkHBUf
5mVOQ2SOi38GQcDSjsX4Q2wY0Adueb/gee1d+BXC0xw5aOkyb6xnfgL+PFHUMCowgPox6TbdvZxI
VKkDUYYeChZfCsBQEd/VRw4IBxmMdu1mtndrMA6yZVw0HpfbYBgg+hN4yKMKQZnmzAIG/7eKfM9I
MzEX1lDA3ZBi4qUAUPXMrTLOzm/+x4EDbvevx3GF+X9qtcd9azSaiLp0DL5W+muvQum+hTztPF1m
RMitgpJ3MwncxkLURhJCy2G1IdxW3U29yfBZ++lRxP0faCpokbNpUXJRQ9YjtpaxwflElgaxL75a
QBi2g4lNf9lAGqHU1lCGgviuJIbvlhbthukg4lM+Zv2J7Q3rzXMonVd5FPORkSMxo+7u3LQQuBB3
vOr9XPLTsoaNC0OH1XnQoxtMhCR2AHLXGsY6TgD8B1ayjRmeyfgB0Y1FOH5Ysc0Wvgn9AivNOfp0
mT5uMprN5lpsA8SsNinG5rGDIANSywFFY2sc1LBtoQ+5AJAWhXbLvJ0nsj+tt0HAQVGLb/RULpEA
eloEVyzkYxSeVD1iL4YoTTcBpiSLryxI8FdeR22ghyzp57+E3BNREWg6PtxgrbmaS/4iXTtGdDto
ZYYDJT+IDVGBV8EXDyJNBMUvJVaZE4MoG2fEXOoaqEipiOXc7K9rFOO/VtrFBaBmdfjDNkYlGQuR
Ji9SpEdtBeyE+PcOllTs1e33Y0sFip54FNCUxdbiN2qz/S0WUkaYzwdVOwzUagoxtO3qYxjL01Sv
CB733zEyOFz8Fj/W5ZKvZ2K/44P1Qzvo8Ti5W5REE/Keyc9p69qhNRkd4sN/61tOCx3trvVGBP88
oBMO2Jl8qghWG5oobp9Uctt8X/Pz3Z2jmPKs7o8LBIzugbyRFtIlVm5LhRwgly37/ccdEAEofgt6
WJGAIIW3492kHrvTUJGC7R0yeouBi1/lgZcULTJzJCiocxdm0VEnlCNJ1AYSGJbQN5x1zUCoqTU3
vaC+BPvIf6ZbevsZHyC+mj6Yxcz4OHttDsk4C//aeOudE9vhjFLQIScTMHgMTmMp3D8Uj9Wb6Dc1
nTsD5GN9kuV6JSiibspF305ivuwyduuFgoVfdvyfGnbnp1CAXyLPZfrqYT7FNpO2VAXBQHB1DjyM
AXRDvP/Ko3oQuDROea4Eahvp2Mg0DViLZS01/NGtHCvmYhlHGG7nuImW2NQNwsL9G5xsvx+nAk+w
YKhkcg6XhmAQizg3Pbs5p5EFkcwvQarGzn8uRTWLrc1y4ZOM4fBtX1m7apq/9kfOdc2zeMlyFTGh
+wk18Y7EId3omdJGRqrVvdwdzF35EcgeGEwp0wlgsgllMWDGbKqVryGQB0Inj2pH5B+KFhiNN514
t8lZBzfHqXcxSPifh9littAjyyQAMUKoWyvI4Jt9SgCn6BSHw1i+FI3qq7OA/zNAX4eXcJUA2GZQ
GZEt9eQGzwufAFl9wcf1rdelF11D2jqHNZXtNPwu6QclM77Ho0el8Ep8ATzBaj/oJMhtbcEzWFsu
CaDxrzqhXLLpi/JxvIG+ZcySeQtnOsf/Ye2SK0HHvTMC8oEkGWqsJ4LNZjRhT4hmUyYXDP/b9fPN
ZI21WplR10Tt5RBtysETxWJ79hFscRV6vsSrYevHQTceg+9tS0oq/ulPex2MqJDcNuN70q0LuuRT
+hjVHpvprk1g9U9Q/uyhdAOUJg0RbGKlDEitPBemHnyB7f6IynCZ1ZZfZbbUW8HAbLHUkCCta5RK
tzdeYIipyTXHF/ByvJKxBzas77Aj0qEsyUx1furJ1e9f8txs0zIi3f/JDFzZiscDsxiBqeBlS1sN
wfzfA3HqMw/cUcqWDCDlPGTbdB4mqJRplMWS+BCuAYqmOyiG3bLE6BbqSG4/FniMk66anI1eiUUS
nGQBHqPaTjjc6wA1y04w+kKnTi2cyR2nOTyQeTu4z+NwMW1ijWmi2HN48nL7rEp07JK89c/hlfzh
CpXYVxitnb2U2OznllHuV4boMJlo7Xul0Qa/G/WQ96bFNOtTLPByc567+TJyMtkTIEuq90MJyiKO
kw2MEQX77VWF18Y+52V0kyOOa2BbEQXJfEl5Fu0XovWbi41tD7bITZ2nKdyEZOesc/+BWRaupZz6
uAnaRlINt5sq54U5W1rEOpRVY37M63vj2majwXxU0hdbQPnPUfgEsVRqOn/5axrmN10vB9lTIDw8
Lle7H8f4nZMEGSsubRpCnhzFnLYFiheT1L0nSAePSqI4ePqbe1vb/0IVs/uoUQDZsGuxS+FrqYUA
Q7SLZ/bUt9kANep5cmps/1pFu3pkB/OWkm/N2pBw0FzkIxoyhV/ge5Rid86gIbcoLt/Yq0RotPVb
rEhKoYm2TmaTWOHwpe1n1T9x8YXI7n4LEO3DqkBti7Ou5SapOuPVA751bzrrCpVlaZbSMyr/MS72
KglCpb3dgVBvH5O3xThfaagDYMPJTFG5NhxUEOPWF7Dfc1+9DRh5iTg3pbhGkjp2z5k7LlIwp5gj
MBuIlFZzZUbFtBaqVyWzH9TxRduERvh08apuTkvFC7zybg1cqyERyMWYn54ouyfdzXKoUfK6Ko7J
iUrUP/YCENOCIxoi/uC0YwaBfLIgo28PMGRdCp3JvmkqFtn8xbKsreVBdsK7Ipd03xXK+64MPjdu
PxpVFeytStpc7IUXGhKj4AjCRckxWOOeR3fhGs2Cm04hkVqAshQj6iqiEyHQXeRArrojj5C8+QZ4
AWYsv/j9S5+Ie1+b/a1wg4/z24YHqWk+e5axNXX5aQ4OCcCNX1eq1K+0E/csH5BCnaNRKi+YXNuJ
g9aCfbcJwueulDWBL8rW1fJhibQF+44kJgPt/+vM5kit8V9HoV8=
`protect end_protected

