
	parameter					IVEntropyWidth =	64