    parameter   PLBCapacity = 1024;     // in bits
                
