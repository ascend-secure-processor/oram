
//==============================================================================
//	Section:	Includes
//==============================================================================
`include "Const.vh"
//==============================================================================

`timescale 1ps/1ps

//==============================================================================
//	Module:		ascend_vc707
//	Desc: 		Top level module for the Ascend chip.
//==============================================================================
module tiny_aes_vc707(
			input			sys_clk_p,
			input			sys_clk_n,
			input			sys_rst, // SW8

			output			uart_txd,
			input			uart_rxd
	);
	
	//------------------------------------------------------------------------------
	//	Constants
	//------------------------------------------------------------------------------

	//------------------------------------------------------------------------------
	//	Wires & Regs
	//------------------------------------------------------------------------------

	wire	[127:0] 	CoreDataIn;
	wire	[127:0]		CoreKey;
	wire	[127:0] 	CoreDataOut;
		
	//------------------------------------------------------------------------------
	//	Clock
	//------------------------------------------------------------------------------

	wire Clock_Bufg, Clock, FastClock;
	wire Locked, FastReset;
	
    IBUFGDS 	ibufgds(	.I(						sys_clk_p),
							.IB(					sys_clk_n),
							.O(						Clock_Bufg));
    BUFG 		bufg(		.I(						Clock_Bufg),
							.O(						Clock));	
	
	aes_clock	ultra( 		.clk_in1(				Clock),
							.clk_out1(				FastClock),
							.reset(					sys_rst),
							.locked(				Locked));
	assign	FastReset =								~Locked;
	
	//------------------------------------------------------------------------------
	//	UART
	//------------------------------------------------------------------------------	
	
	UART#(					.ClockFreq(				300000000),
							.Baud(					9600),
							.Width(					256),
							.Parity(				0),
							.StopBits(				1))
				uart(		.Clock(					FastClock),
							.Reset(					FastReset),
							.DataIn(				{128'b1, CoreDataOut}),
							.DataInValid(			1'b1),
							.DataInReady(			),
							.DataOut(				{CoreKey, CoreDataIn}),
							.DataOutValid(			),
							.DataOutReady(			1'b1),
							.SIn(					uart_rxd),
							.SOut(					uart_txd));	
	
	//------------------------------------------------------------------------------
	//	AES
	//------------------------------------------------------------------------------
	
	aes_128 tiny_aes(		.clk(					FastClock),
							.state(					CoreDataIn), 
							.key(					CoreKey), 
							.out(					CoreDataOut));
								
	//------------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------