

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
caQ4kDNpC+yRhd9rT8TQRjEh5dHwq37lgHnP3RI5sQRwfA7zsWXwbZRhGD9ikfspHeHU7ayi3OmU
WfEoUTW8pw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VFnFlmJ3J1D3IRh9aa3aLQlPXF5So/7159XiX4axP65bRTF088ez5OE0uWO8ayvK4YW3ZqYiTOOw
6p9P2epqNjkH/N8i8ZN5SsgJ0WT/dq56xwITEDoGQp6E8y1M9iB5e3Zs60VN8QiK3xTd239Kb2Is
hT+s2ECmzEqJuVm3TI8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
24B4SGNCPgvOzh0vhtLN5279M65nzAa+XDLRI8Cw2pv0wf4YoOAqzpljAP3KvdJbt7+u5dUe+Abk
0bo9eO3SfhQi0EmJmr35x3y9MUFrD6V0qKHNSlcfavPNdn59fAyIql3Drt/x+RVhVZWrvhXBdq95
/5O1Yh2EeLrqlMpZtUAX3NuKrFlVe0pq950XXav0uroscTnf4/E8Loc8mG6O1sYv3UsREH32oL5E
V2Yt408Bk3rr0M8fm1mtKwXy/yHscGX0bfEtFlw2yBf/V2lqnPdBkOIdRFkZ+hc4vmgrL3zC+u3c
FSfumsObF4ymosR166ClBdZcC4XDGZtq5xGaNw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ovx259cNDtBFa/oJJBICxm0yvz+h/4r7qzgrTH4KP8268kcBQi/sVCMnbjohNqICo+/7l8gEaAFO
fqml5lkEdgGR/HZ3l3n9Ome0tTbBZiNnyAZ8QsE5/wugnKRozagtWPFRBwBNPboFN5JFDfQCNnW9
DNOUg+hIXZ6UYpUjvT8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K/IQQ0giJwfKqgjeL4+9+HSBTNKM2ovuq6Z+1C9A+q3EeDaIdaKKu/T+ZpCeDPYUyuKubgaG1HFN
MVGYVReTc8/zcsCueJF4SCCSjvLrqJpGqI+R1WxFRfqpheXCnilqSVpW+QXRhAznH/pS4qYWp6Br
JkX58ivBK7d0+qWjdNaVIgFAPQwa+zBDnB1rFqFki0yW8C9cHai+7CQXpP437jSGbX4UaE7vxDc8
7LtIslDy9Xexh+dRqaSdV+vbdqT0/gzea5XE+qxW4urG1TbURNc1dsqq819daBkpNlzlbTWrQi4E
NCnk/sVRC2oftsggT1HR7Wow02cXwEWoKGzwtA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12224)
`protect data_block
5e7eGg+opXV1tbo/prF0ybjYNrhN/w0T11LBZ0ObGC6kGVIjJa3Yh7DB1pbMI+5jaCY/edBPodB7
L9cETWN7PyBnoDtaValjS9dsoS37sm1U+18TSS6uVScnyjvFPO70lE5BXX6sq0b7BJ9qihkGysWP
irw15SLmyWIAqUxgxqJq0vHVN3B7xQuUNmFgMIE2+40uGWXN2AdSBE/AatFuBYS1kXoW1caQB01s
1s6okVpGvf55LbPqDmC0niyC7kEacYRLAtZ5zqGs3smxZh+f0/Dsqg5Z9PrqQ3MnnEia4ZrMzXMM
e6G3rXQ6/Ur7SI3j8mYPQLXlkpdYNheiK6HouppGwC63tlgPPSBEFdTlmnmTES5brizpwLle8wyE
cEbDRYlMGsoxxPQWClAOQsh7cj740cth7uvdVXxEWQyt2PmmHkcwDfgSRrBkANKUS8i0F2KRnpoU
xLHyl7gK2QlT6trVDzmHqCTi0y/QBmPNNDNSpp6OpREvnsZl3NEN/xpUjcGmWt2mF2ZcckyFIx/Y
TP9p0PO6vj93ZDCNEI9OPOS098EBModKBeyjeB17eXRP3goQ+2IBRI1vLy35suZE18LUslPkRXyQ
xTLOWlHoomwInAyqvP2L+fJfdeA0pOI9hrzjU4sAV+3Kg7a2Q3W8hxtD9jtPhn8dDQzcc/202M7O
5gPZDrxwdu5bxQi7hZ1l2cafF4pQuG4OQWg3MJL1vNcCR34aElLsXfUYH0UtGsf5hhNjGAaQ9xMM
8r7MSwtjQepl5tHPqP0JQ3nEeSy4sB0pwzE972k8QZyPyoQCpgI7v7vAPs3rROxVt472q3yX/Gy8
mwdk8W77wdvnytnOUktseGQwjVhqAJ0W8uUOdv2XqQAlEPCjUqYJZMkc7CeZpx5yjca9VPIm92gB
4+TlwXvI4Q423fdVSUJFLutoaUXyyiqhLX2pYC1X92x3KMFDk9F+0n8jLuoI/6552SECaVUhvv2U
A8LlQWwq15e+xe6wYi+Et51pNkxCfJYkdeUqFZpUQ1gUBoYuXWq6ED9b2qXAelCmZlBNuaXnyFvc
0jE77SQR0g4JoAx51CzV0aUj/qx05CpeJh0jDedmdLV5JeLWyAE5lbvxnoIaTvF4sJK4+iASBfze
n8iqCRQ6ay5Nb2LPty4NBsRGzMPFrfA3u9PJEeZ2pZ7/VTbAtZ2VXGy35FlJiY9OmtvTqIJiMkjY
AnP3C50HFOsivvj6fRKQ0T/fZIxCfpw3AVv3Zawy4EMaRhmqTG+EgHzDFnzZQ5WqM8srR0eYnNwB
lOql0sFTjGGeEn1H9BaQncm4oBB7oaAi6sqO7r0wDTy9WuxUse86bo77H/bLUXVVkEoKv1Qc1i3d
/yBrpLmOAVgC8H51e5W3pe11zDOhKO3y09U5eG6OWq7dQmaCsTLKn3OefLejcVAAWq/G4EO8M0CM
8gv2kpi2bX2llyjI+yecq2+qlThcLcfK7vZTXNuHJPVlhA1CR0ECri1CGAG8kPkktU04BADICov9
H8+8keFDW4tI6ZY+PXyhVcKRmLxLEysZFtGNm/6/4On5eQauEWAzNlNGqKMWXsyzUd9NDvlAZfke
5qk/vyQ+CdPAgbRLDOnrvTpaVIdaQ7WkOpfaAihP/6BsaLxu62nuxEP9/mCujaT52J2juAqmiuM2
vDtWdUn+cu1fjFoECfn8nm0slQMKung0J5yY56OfFiz0TZ9lw9OLFfMufSrIKrBLtLSrrh3PyJ77
maTCEznfFNzjeVmP+Z3Rsq7zu9iB8wKQDe0ersut4qlUj8O0AoVPGU9BZRTyS0hvyiUG3PNqxTLV
6KBnCJVhzaQYDbxXjC/i0BCEcrFkuUmxovqscBISrGYal6rQoVJ0xvo40TprujYrIEHpZJ+BlTXB
ASx5oHG5Pfi4fYyKg89x/yqPPwS7JOYawUTg2gU5PXL9C1+1hM4iXYHvTOE0QnKpm4HUJidmCBtZ
aJPKXNN/LSPK5qeLCfU6E11718ZZRM3wjWtHwtT+wCGOc71/P/6B8TMLCrt96HdyKfc1fEVWuhMR
DsJuuDLk1UAVnJiXa5frBRgYTBKcXH4/fEsibuAm9XQ0xKWr7XzWTYPwf49gD6zOoyfp3yrGYr4/
CUzFYt5R5JfPJFdBp0rzwxjwHZH7ml0Bi00n7y5XaWq4P20DnWZdgDa0mP4uWxYUO9A0Ca0usPJH
P9+PIPan8aS8fu3EZZoqoG6/fJqWcWBCmRGPTwRtYxpF+P4ZI9CgvHd9j801LG3Y1mv2fFaMuWPl
U4dYWs3uLUXx1JTA4NUYcoaN/+V1X1m4pMUGGdkLQ4Fjkv/moAqfx1GQONpp4IsOvlSHFE+M42q9
s0djTew3hrvyD76Oe/fhI6ZrYbX8xrRWkn2IDoEflTJfcxSX/uTEJ88DQGqo+Fm25sAZEgr8BR/C
Y9BY7LA+WSKxhnMTst/ji2BgXOaZkg8wc9/Rfm8LNXfGQzGIwrUHWFHFtrN5Vf187PJoeTUpB/KQ
KTEU3DeqgLIZ+rC2Ze2rSd2wWQPQ0VFASvLbnYPB7y/jEogAyzfRxEBeTQr+sTvHpPZSY8Dsy+EO
4a7JPHALOopR/DrDBW9ao1pRQQWmmdE6QFD/Rqkk2KPhFydvFYQ7MySesbYvE3fteF6GAzVe1CHD
MFfe5Um78D3U6J5CRBbjwAsFVBRIPc7NuWvL0NzbYAZAfX34Qxxkm+ps+3EP8Mnft7dhxb5E5o9d
jRK1cAo7WSorFwNtXSmKEOH2Ul8ir2zDG8WHRtvWSBNqb46xEUz2vUJLQ/cRJHCOdvFEQDTsECGy
huEGm95Sv2w5qN8H2KBXrQmYpSXQ7YythZCvM663UjELKswMZhdLuF48sdiCV9451femGfwEXlhe
PSwfwjGaEN61OOrayt1ay0diG9ZdDSoaYmng5xjmfN8mUtA1YGbK6oUvzX9YKADVxxTuk0hmK0fs
ckUNU8nvVW4wW9p7w1+5fNQnlSjLYmq2eYBN3Asr4sP2QRXCgp6YSt0z8QIwh4xar8pFIIqUc0+p
tJB2X5pDmTisgL0jaQ9SvP3ORQgh2nY2jHnbsxFT8t3XLJf6B58ROg5WXVo+mIWC+CCQSyhCSZgN
3Z5ARlQ5hW46UceddaQEJyYt0KOkMP5dh6ML7YRQWyzE03On5i8O3w9v4sYdgdLrvfrbx/Gs6gb7
EJ6/FLV47oJQDs9L9KXW6bDwF0ubSDmuBzNqCwgp9df517hA6vHMwwUdWHNPL45GojcBRx8992AI
FXr3G9FJzgzNRVUY75uP/V96fO91NXTsDUMnTQ3zqIRilhwWR6Q0bDN8LjwiKUhHZ3wD4G77F1wg
HDs9605baPEVrK6zUCIV023Ui6RoxHOAqkVSjbLiJbDKWyBtPkti+GOStX/Ga+tYeo75pf6IVsOR
5oMwxSsTWTRvOBmzGsOqpPbHbBpP5X+SX6jIodTwTJRMfhpetFfgbsw6U5u9af0td7NyZ79P1/zr
h9SJpYq8IQXmFQsZrlLoFxPC8g5dmwkBjYZFPGudoyzl1YnOYVySvZqfJIXuVnbB6D6pQznTpAtH
H/iQW6kSe5V7rDpiff0ATXFW8QdPnQRG+IOkAuorwh2V5j2OWidji+RQsFyfyc4Vh49Ax+R2/8M+
lVRr1GXO1jgtFFMqsOB3QzAK3M2/U2dF9oeklKqA1Rv4YcYvOMlSKHVR+qgZqSRqCKFZQfiS1xh3
Bb/WtnO/aMYbsCKui7ChhSUZh8gG3LzCGpAdKEjc2fLW+Ennyq7sY1/vf8CT6o5MUI0yx0S+QcdJ
ucRz8i9GSnlugpWKOXGqs5Izy4ID1qEFHuY/ZSNUYGszhJLvUnGFjT3aFaiMfukDIUCM8JbUoAkF
S8VpEvhdc91ItqyXG3rZEuWESFV5cu0OhWD9f2JFzS+tmxYazn/bp9gv/5Nj3+gBh1e6lyvxyAmF
9lFlfbcu+adXjf7jqWWG9VvwzKZ95hkcPNY0ZtG8rq9BVaV6SKqqZPxgtf9KOkV5UoGQp4+nCJ7k
vvrXUTQkaOhyvR5ZmnfyEAIGpH/mZUYwEQ3YAifnNEt7DIaXmyZQbRTDJt/IHY/IdZ3H7N4rmRAi
HszY5O4MzK0pX+Be4VrfwzufJuK2SSgoL3RGAJGnycNp5QNUcEmu4Br1XxeoUfp0MZ9Ifl2uC8GU
9Eb0nLA8RuenKy2D7w4iB1apOSrvyDQyj8AB/dKvTjNe4FPBRsGtmIEzcm3cCSckGOCdejU/QpkT
REDTfQJ8y7s4qs79PfYj0gMGJAus356/4UV542e33GM+bJUrl0Ol7oWtFAzuAYZyMMZPPNUL7ggr
UJbcOSAMtUQUeQkDHZBuJp2VN4ncqhNFouy2TwSxlDR4H60veTcud4SFEcex611Z7u+NjT8JEhV4
sKWrEDTI/06DT96+KUhMCTMFK9flZDFe2Q/yzvLDbXDHMH9pFH/t9VjzochMVZ1qWKBxdMdhflFU
E4JTCQol5Q8xaWwLLOV3UwXTaR4FSLx5+4Y1MUbNGe8vDI2YCvSd4pdXaG6m9QPtuD8F9GQbQn1X
YLgpqVOay+gUkiY6z4C9Wfq2gYR5SX31/s91lp0uP2evquuI640QdMkiDYjzwSJTQcViI5SUEhig
ny0Jil3IxBc8dRVn1eoOce55YGgdC8YmzsRnxFjWLklWzyMehyNEUu/0XM9+EZlckq7O+ZN37/i3
DYyqsqA+nsWdevHtSQOofFobh4OqzsGW2P2IaYD72MK0suhmPksLgBFVOFi+vzihzLpSCoacaGL4
I9gdvnYMjORIbmKAUUQ4v+NZTnn3b8oZO7/O7cZHssaJYEpvf3uTvyO+AADck9xQqoxs2TMmdFiq
NvAGCbnxZYwkwMEOgERZYUipmmPguWhyu0kQc1rqPLzyPOPNseRBVlBK28TZD49fXD7rxMg/rNTL
x5P94CkqdZnL4lIdmqVZCCjMVnxnGKArbMJZtL8U1bLX3Ux8i8ZUEQYYU4UYzDhVL+gfxQXJA2jK
zvf0E3DhwnjjMhReqIEHkgz8VBCrIBxPITuAwtvR4n3Zv+nWdenkSItTvtTgtNR4uYemkscb5lCF
Z/0Bk00p61S2wB0I3oiJhT3+QEBNtQCYCsVTuZmwUxEQ0Ki9FKi78w/LkS1CW1qM9dCDnVwGlEvS
F+qgT6XNJuvpJOqJfPr+kt5gKYTU56JeYAtMNsQrPXDukHiJFpbpfgD8V1DwTJk9PUBCBU0XH7ZL
Oa3iutPUVfgpO+MEqP4Z/ykpzio/v41fPAX/xl/k0ThjHOzs4N/AywlyH+VnKvpRO2vs/wYnp8RX
rgSVgHyae3vDs8uih1sKb2MllIKTR3Dh5bnjPYDlLrxkgI7wdCVFUPjKRV0HzXlT9ieXYvTMT6C5
e+pdccurbzR/PVEoVbBhAWtz5Vz7P69AIp+np7lqjigg15ObeB8fEtSv/Dh4mhqq2yrC3JV1f0MD
u+2lLi8sKlmSLfBapNQa9lyP54rvhUt7bxXxx31gPKdwYwcRrSphJpQ4/lewOrreDZMQMqqdww3r
DnZb2uXTWXvL+bwm+GUI0WKWYfvOnhyrSAwz6xWlVwwy8sxkLU5AWzn0WeBv871QVKXoskqjdSdp
3iypfxsTBTG1PSFkiWAZl+GnKVzQTrJwNrj9g1pEqzZZCty5huxto5m+dV4wq73F2qKGpTPG7aPV
Fpx93NqPg9NgK9Zf9OQ1FtdWBQBptF7OYFKu2B3OXR7shimdiF/McCfdlJpdp0RWqYOqb0zWIMsT
0HnoKDb8XE3ArBMcpDAwKxPRKCu11BR4SZBtzUuVJqXNS7/BRtsP4bip8ylvNskZeQLozKLMmieQ
i+9IJYa54eM8ZSS0SlmiFakJEF7LUhzOXLnCbQXyNdnUxJcG41QhPly1JqWTSwP1cpEGDA7zUWZd
y55jTk84HWT64FHtfaGt/+XsCcilSFquAMD+WPWotzXUPkIRaVYj7R1mSPfl+JIlDEzGYUsykUox
j610kRZVckvesF9pWpw74OxE8VkxwD11wdNlBoKyQJIbWDWi54y/9jRrwMHWJmY3gbSFPsk/obLz
2AjDpCwB18BZSVHUbYKqubFFHiyf9qdu2VFWcjRGGUGcSGve0DjLc0TOc4GWsSxdvVKimxNw+2hY
eFuaKyout2+pWa4xpr0SE6tHCqXS/X4qFdEN8mMagiULh70wV7N6wZiHhpSDjwxvnRRGv+QmkxLh
HoHBblhSQ4U0mbpbwAf6r+gykUc3tOQXWLTtW87cdOBlqmZV4nQGNTnJY9a3njtV6IQy62pX6gLF
aQ6FdsujlalX4xvv05VuWZac1+SGnzFxAE4VuHovjeoIWY8RBQQhNu1kT7Fvl98MNDSVSvDytPIc
zkpYRl042iz1FF5ZmbDuXL2nzIt5X0DYg5829OfFCXCM97nyxWrY7wYIbzmOFjPyVS4K/alDRFIl
C8WOc2HmaD+ytJA8rSoSQM7aGShKNrB+3PJbPWntX/2rk0pPx6pg/RqpkeHJ+MhDtZ63zspFjbdT
t2gNN17GPt8D7m3XGcBbJOCJRylMFP4+Tp5FTGXVNVwyS8XroPIabGf/PL3H0meh9Nk9ueK5MiSL
IwMVPebxOZYtMH7qKrELTDI15dloer8v3HHnN6oB5g1FeL5/g/nJh3JzMuiHLNwCTB+/GyQ75oQw
RuEr7Xouxa/scQnzWfGhUmIJeDPa9EPf0zEgApXJDl1uG5vrGEMO6I/Z5w4t7unQG4AfK1HDV2mw
niUEY2Zc/q4pfVZPKWtkbF0TJM2EuyB/4qDy3s6mn8HwaqjjPy/ytbLow0Au3MqscqF8G3pDtcCP
cIa4MNW4vNleRnvnARygUj8Ur0qPb07NqyMK7Zbpn/ZabL0ULR1dQNyDu1NIMAmKSBP4cA+a24vV
+cWuPbyP+zMiNCtMS3kRUJfLPyq3v3ZIpyVXu4rM4NWA8SUgwtcNjJww0BXWh+tHJFWmvR36C+O0
Z+Un/MnmDyvZ++aGAN6wm9IG7uSP3mj83w8up4yJLzgmR3XVU0Pj7npipwMnn/8h17FyNp7pyEwR
PQJpCrWAfHAFUY7jKGMNLY5MVs2Jt6jI8/iWyjNYLqp8BCbuCDG2Q/NEmEXqSPFzpwlaD8xHNU+l
G0+TgL6Py7X73nyF8Y1MjSulfqdDabHUCt7cmhD37mRntR/RkAQIron0OnnUVtINs3me0Neqpuub
XfNW/XX8eawe1pQmKIejWn2Dqrylj2XSi9ceiDUhiaqdRpC+KRXEi9ktydg8JkoDaSPTXmTlGrBL
qSohgQIrReEcEIHzG0CZn9OVnGJptDNYoxnOX/1SexW9q2l5wXiR4Xr1V+r8PBPWp834O3nLcvHR
LmuzWTqLprSR1/E40PTS3A6rtHgpLF4QO5uFcxJlDAylp2JTJGE80BqbNs/UDYhwRF9egOdfpiJ7
q4OcKI8gWwwphnh++FOZxmzSPQhU3nLy9JtHZ0nLMfLMT8YYu9p6Z7vIJq3hMzGvDEZkKUpbYfRL
ujIdV+Z1IC92AIMV8kz9m/DldPTU5tYCHvrFp+DB2Eh379JH03YwIbjnAJUs6D0q8Cg+VkZMj69e
sjSom1/iLc5RHrd+ZKPk7C4pYAO/XmsLEs2h2s36NoR7ICcbcST3ZmfjpKDj9qm88NpmSIig5laA
o98ck6paKmv7cfvz9Z/wPyP+RzNZydMPT0TJJE9Siapv3Oar/ZhL5PuW0t49wXeo/9dqiCNH72W5
kzEqYhb/6Gh6U4JDj8UKh9qXRb1eOC7deBL9AEy851dFecX3tI/mJRcp8/xIoQ7/JY9bK0vDyGH+
cYp1LK1tXyXWZpq/9km9uqKz0Wlchz+Gt4l+yAm29Qd2GcdwDs1VVmF9HVPSctNlHvWGBrTbaJsm
hYgZSbCktGBewFbMGs1dtYFAtGnRheALgKM5DLcNcQqas2yzyaW0fY2zsZgb/MhCx10F/75zwG3g
G4+nHsmliGtBvY3kRVDwU1V7Ulz4w3mJEmVMUZ0mEht9X3SLVUe8PoBuJMSX07GRi/M4C5y+8/3S
gd9joJ6QwqtG24VhDCX3iHYSKIGpdWOMhm6ac7Hj4QU2sL+NBK+35VIZnljoPWb5fGIushu5rLAJ
vFBn5CqwuODe0FFli+miIlPY7SHeQ3fqb+X8Pwlp6XEFOCiPhX8u+oLJho6rK1MkaZTsHTl5Jlly
MrkPXdDAtYbZ6adIpY0/O23XaTaddsVwGt9SRHpgZcoMNlXBtENJMQp/3QjP9ZEyIfiUsjTsWJ9Z
pzzARo0fbEFp01SWtfQj6hMMNXUbdbCUMYGlb61ynZPf66bFOoFlAT1D/AjLRYAxqV2R2Y658E/g
BMq288YEjXkeZVwA+Lqk5xS79oV5QTWBJ5uD+kZ+UpCCwe6gfRwF4o3Il9ddXPbVMn9nptYGaSfI
xhyo3qqQocz0fSkYcHIJi4ovC+P6LUS5hAUU1nr/iys03AmoNRqOgLggnW4IGc+bpyaDbEIq02xW
NfqFhGfnVD3QDHaHAzWNaGABwPSTd/jr6OPEj7EavqZYKlfGJJ/jPqqEAVax+y6HdqBsJAA6CTsZ
/nOGDDd6gLKGE3bFup6cmcggXRNbgehQckkRs5lVgcs6HLse586N1KZa50h9Q8mlch8fn0RFh6N+
obhabKkhSTJuZOlWWZLrgn3LO15OjNjMiAbXlnjTuc8ltK4lslbnko/zGeBizHDDjXiaU9ohm0/j
lAN1cb8+AOy10RhdNm8HesQoNCQNxdG54SHScDrMg/Iw62+1gaMGHAIUSQt/27KX3YqBDfo/GfcE
MaFuuqAFmREexQqz1RZooaaqy56A72jhp03ty8Tvl0b7/NtNvQazHHIjikWw70+Dfc/oNqOj/Zc3
LC2k8EynSkVlzWroLROjbvBFUziLxGi14oiPSGUQqHKO/UnkfQohK58N8ot6SBQOMyL2NFlf2UZC
KnWqUhDO8fNPZh6Dn705qV0rDyszvKXA/N6OzpeHsea3ib4CuWzG7SBKOnFKnIYT/4Kyyo62JQ93
nqLN8+HuxKC9FyxLAHiApt8HB/Zs2b6LxnTKjAouLFmpfjJ9mrB94oDfglf532BftIll8tDBSLil
MEuDJex30LyOh3TvvctazJ5luRI7RfTE/V4SbtAK7UBTg3ZWeEP2Ev1AmaUPbnzSsMGAvNPZqih5
C+Axe3WXveMtZfuTb2RY8na8DcUkU3tbeEq7TOZnBFDkwBBEKnyL25y7NC954WQ+ohvZWMQ61jtk
EnQFohksoigS1d8DnHQlT2nG3X+AZaF9GjxUyhNMy4KD4nnHh3vnJNlL9rBWijKep/EpM7VmBCiP
fvYIihNd/DJR9kglYLuSVSZTchRMBKOGG6pQnyPT1fCYtj0XzY9axZV25GSXZ50EcZFCKBUqzKwq
+BIr9Mymf7lhohaETTotRHeeZttEq62G7UXuBNS6MqdIUavD3vcAa25hT7ebSCgP4VKLAUN+DHDT
cUwWMo1caMd0DC1zMi3rhyEoqms78oLJjpiUQOYLosUOEfjlv3+iUppGm/4enDuaBTXg8txdBQOs
A6fUQtM/4ag/HtyieXqXDi+6eOR7mO4gWiv6zmZNaSwOqGYd4eLm+sDfZ6PiK0EqogkMsg715JoL
Xr8flZmr/oSxJ0vhol2FOrahuJJZWHba8LWSnfDOnqVEWuE/LEuIl15ZwRiSF8QFcClRPiTGj+Cn
ZDN49sYENetrnpyf458Kmrp6g93/Us2ScUyBzWRBEUSq6ZzCtRQSLvzo7zXI/3DxiVP5yshFXhUH
M3BxzilNBvKyHkCToKzy8igD9aCg+wxskdV/50XNzkpr6Mb1if3Q+ahEJDGOp3cS9379jwopuVR0
Oub83WUli4cozz9Bns5jCnfzIisn9eVwyP01jchejhS/tl87oxberNaWF6PZ2Jt+00W5ma3i0xjQ
yGUEuzLCBbPFGeYzRsgrs10YDeAEQRakrlFKctQfKrCwC/6cPM5DDiPePT4U4gy3GAC3FuCO+JgC
krDoH2OsaeVXC08lY1uv1ZlI+qeiByi6p3dmYIXfFZCeB29ayx1k0cWAohW4jEJF0ga5crnLCcAO
jt6Ar+TpNSxI+6n1okf3UoyC/VDJcwdFgtU4erlcKpqgCjR9Tm4kkwrjcVlfgsfyCPvKjfiZfHfY
+nQLYId/gAKdbRrx+XBr8a1DETxiBOsL0ls+Zsm+zlAHxzUmGvYVbjBgStjOQpbuE6ifUuae6fVH
i2xame1GZ/s9KfxrN7uljll1LR1LVqQeuBnR5Aci/U6EuzN0liFgmdf9MfqVoBKksxn86C4NOTGE
dG4z0mqZeHb4583de26j//pmzeH6CgwzEzVz+onx+VkzyvLshOHTdM9CsO7zTG8f7T2+pTvRttLR
R/c5x142zg9R0Utz6T6ueCejjNXQoZgIm48uOVCWzG++2UkJQ1NUAyfuSZ9okKmkoGJ168vLaSu0
HziKTGf+1mU7GXJaSK+b0zkZU79R5DmJGtFz+Yzmdyvd6xRfpV0cGgxeqybRF2XuoC5lgR3gEhUE
73TjHFIXBhVY+uwvUBCv6dANG9a5Y+YUWhFQOxRxo+YCGKi1V+Rd5uM9KYvBoSKSHxn0A82ZGRNx
g7zjR7WJ7V+kAHHOsMG2D9TJ2YCAe+vP+scUFo5/U2e8hgMq96Uy4zne5oAjpKMD7o9V4jv65sWO
UelvaWrHpPAfQxC//fe3A/K398suZCSOf22PA2k0MTBzr1JCp/FqsODg8o5RKl1cMzlSWBw6If9i
ykH3BTntpB3KLCcoBJKVNi5M3NqxdYcoGAOfHeuwwaA++dB9G6iiVE4GIjPLDuF/ZOJOLwTWDUSh
Eh4QZtyq/oGSRDxs3fgSh405dg1fTfU3MHTQPqYMSfk5V/hycqDPcMDjESNnWCkNL0CCqhjEJRy7
lV6u05zbi4Iykor7eTED+HljUWh6j4VijppArM3BMsrvEnGzcxXfkyAlonsFUMXtKWiS0KCkV/y9
gOXINY4XP4S20xB/DbJoz6kek5IjFiuRhDPCnZHHbVAG/21r4yRkxYhdM7oF+VEHSlkNmFybsLHr
miwevY9TjWjZgiqteTxmu+KC2Q2sV6bGiCPTyQdKnWB410FzYJFnQb7t2Vuqxx+o33/x6dlp+aBH
f6e32Wo1q2T+Z6pZSHHbmEdpgST1d3iVulbF4iP3+oZypy7j7bb2e8EB+VkbYbD6X4lWILhBHwxU
PUYaepp64FJhAFljU55d+Atyl2YAn48kPmEIDN7fDKzlGlALUtD8A7eavO4TPQIcsbfoA+SE8XIT
wxSeK3xNtMr4YIz7wXW3vOsv6tmZzh7KBULiYRURTQOkJvAGdFlNIqZLz+5yIOdX9y2/VferLhu9
cGnauGRCF1g0GBFe8+GTQjf/zV53cGbDm4gPXiTPJDBXYhYmsWc/J//IbC/VnXL++4vRRRNbDjFk
uAxJYL+74TA33uExxjjCJ0URh2KivzNRkyeKAbrMm8Gq6A98PzbC2J5LI7ISaIvTFLIUKq7dtvHV
y/3uFw7tEgLaecuZQKGdigVo+yZRRIxzDk9A4Cmgak/1cXt6M03x6nGmvGfle3h7N1aHcccjqolp
zu7VkhKsF7MEhBaiamASK0cwisBexK+Bmp7EFMcEff72/5qdMLz50DjqvlcbOkfwvqxdTt3XDzBy
WhS7HBBaLsGO0+s4cam3lrusQdThajm5q4Xpget4D5Fmt4+KMyrAW7MJMXwtvXnI4AVf93DozUkW
94K1BOHMp/2ghpoj8qp0lguYqZxDhahCEKysMaynKj12VncQeIl7TKpFYtVFHh66bxPOwVQ86OpO
7eUqOhGvC6Jf+7sCvBB5/4p1P/Q8Hk3dmLm0wK1Md6sxtSCXpNpe+NfT+ysPWL9Y2/17PFnNGgXr
+IfeatcnxPp6uUhsDRal4m8MP7nTO8FcG+OPntRg+F17vNR8nLX4VmrtCJnLLyrMJ2dsJhzYJRDs
pxALl1KcWR7TyAerna5M9433Y4pUivRdTBe++wuF4hLmBoNFjvZmAWPckHuNghDpcZQwKgYRssEZ
okkfTgZEcfeL54EHqRI2MncetkQGOHSVTmx1EpsmJX1O8MlevAHTuuImNNaLY4dWBm0kA9JVKdXm
Ck+iyRbBCGKsQVBIIdGQMHwZXEmrI3Cd5NWuyq0jiDD27nKHY6KdjGi1LvUHcIHxaZGGe7PsChQ8
8dHqLO0Ydu7VXKktK2Hgc/vhY5Fv4RzO368MsBh11t3n1t3MI+vk/udDAYlwJ3e+EbleCECVJeK0
aMKWVtB7X7yWGFXeCk2TDnBJCUlJF18WNBRNr535zxZKT+8T1VyT25SjFbJyBRoEwAEVfvONEDd9
Jf+DMGIf4QA4bTx3h5MCpHN+9GmFWaY3mmVOeAQlhyiA2sn2yY/A3l8f6P5agL2HbukFzzk5JE2x
yGO9Y3ZJ6eJ8FRYqKPg7CbhihQQ6zcns4hdENU9PKMPdf/BRzxygSVVk+pht7khH+nnSTI72+9/8
JuLbLMgZ9hEBDsQMBSRIls9FU7QrlAnI1fzZb8BwIF5mE7Awaccdkyzakcn1826QCRLbMjDJMGjC
KK98MJjnLAfHAC8AN/pnz5d3zR6Fqbcx/vQB76e/O+E7fGxuzkWda3gKQ3Na+dKFyjaAQowe+IjW
AEyH1Qa2QFEwDLwMAb2DgttQ9g3u4z3Qa6ziEcPHBtWgcNPK3OUVtunp09ELBSkaEjrxYGevbQ6j
ds8U+5ogyxet3d2NS4MS2W+WC3MIj2rZQr0ILYbudJcTtZhuJ0H6hDnX6czFYPcvkMTILqlOEuwj
co8kXl5iFXd4fAQG2xXdIwAskz5wIR1Hfi6BeQclF3heqI03vUQS0srmMkKTTNUhNk+tr6eLWJDR
zZIT4VEKVcgnV6fNxPR22V+KNmVMxiMI79uycwZa5/GCfxcFlawiLp5M5FKhnUnQ4vCPUrJrCGEm
jtYRF+2J9rqfLc70aH9M9AG6J14AcXK5go4dkuJnIlsBfJcfSr+ouAxAqJNp00Roq+1Hp/5Mw9zV
pOxKRCJvJsL67A2ByKFIFGWrquL8/1YcaJfK9XPMj7VNQERMpI3pqZaiOhSnJxFd7PF738AQXMol
ZM7DT/j55/S1ZEHlqnuClw4yiri1cXDTc0Q3iEG8ZR4pHe/EETLlYPDf9BKgQSLWDPxByoZISury
JCpF5K+9cNT0HwC/Q4Hdc+LDx77alumA9CnqXK7H1LARBhdw+TS5Bjwh5QQ+Of1gC5kqqVe+okIV
axU0KqRebV6ISLnQTv+mix9+O5E8FY4IXZJbIiIm6Cq3iCK3ocyUW/VuLzs4Vfkvci9k2Nvz88dj
BtnZMFVY6Ep1Fb7GT2YA7xtlcMspHQNIbUydV3EW1SD4j8QJxuNxh0xkqWdq5eQAusQ84dwKXA8O
gVyNQnLEQFY1RCPBDg4NPDwItY8qLQ/82s3kUfHdQQRr23czYu6dcIH207OP15nmOCi8vrCCVPd0
5WohH7JXl6uyzs8K3Zq7JX3x+cN+X0gWfl412eCfsK/5vzsqTTee62zoho53O1KDHqMibQHeDrNT
hamn6+30BXMzEXereIdaQ/S4AXg4o60GwrmYLD4flaWwWDZD1qEp1i56yOj1cL7qPw4dO4BwS5qX
YSi3M1t2gY04vPG1p3vhXvOWcqB+H1q/sXltTSAppSN/j8exR9iaM2CrovS8aj15Eg2rjfQkvP8H
uwlgE6dC67rjJqlqUYT3F9rrCDGtwv4xNMyH2Vy25Z+wsU8AsLXhAX2o3K273T+S85q52bivu3KR
NiyX/XUe00ozH0sUybnAT0uZ6uVcB0LVOhobKQyYlH1XEjSQSNJMhdxEK1f9t1Q9s/OXeEjRp6dy
DJZgN0AswI3d0jibYDV90BzZv7aVQgbCd/GjxTgoS0JtFHERv9dC4a2rn2bQFIEjtacUcl52PSFb
zu1vaz/C0z8dA+hjghoqMhQeK7MDH6/b3Pas5OfcD32+GbXh7NYcmKA06gapFEwQG/6j0KiKXiwY
RZcQRlJmgXjUsN0j4k6yhUEgDz4ys1awttNoPkfdzoiVCt6c9n3zWVMjp4NqUn/f09t/OIGzsO8x
LzCNs7RtaLlJgqN60moIwYvMMyyJIC3gyUP0EudLeg3vOBbJqDW7jIqAm0sMefJclQxEazSA4xo6
cgcf+wzxjIGwgTg8w6mGcjTuoVA0cycan994Bq2iJ2buucu+SFDBGQBH1cmLu4ZM6wo5pPuY74rt
juafdT16nnJSgq+y8VGInr4OjRJaaQ0EEz5kxfk4zoL7nHky6TUT9uzIIMJC+wpHK/Or7U2nnwvQ
EOl3vGii5ZwSK9svK6Vf/9tfo0ujOhF7kjtyR3xRFaRpoGp/2agSSjxmAQWTh4bkEUdGNbdKPHf3
cCM0ooFMr2re9nO6+Gk49q0+IZBkKK2sKDbSEJwq4ADdGjvWJhG/wtUJfbM3EF4f1ypiFF4XUdti
Pwd+fiQDNGgkP91SAZUrFefQfEJ/dQPm4hJcI5eqec86gKCTG1D4hr2HHCpIH3dzCBnJBwlDAzVJ
y3ArRXqRSdAy0Z5yvof/uODHFUtPpBhiT0lhOb5FB1Qx1pw26HWIgBmtmbhO3mC/K+zXgBjaFyQR
vNu//U5vVxzVpKtzqpWBr66U+wzCqc08xScXGLFufQfimXf6ynjm8sPF9hQTT10kCyeqibf0egXB
8r1kNE0N+zQ33376jkEsj63YuX3mr5CpYq+Y1hTh/jFUhw51rUkCws4B/Y/wlHH//a+TjmFF0OMX
PpoXd9ML/4mjiJNkNbIXONwXShACQvFPuxyH6mjacShvwBwED0tLDuhnvnEoXr5JXbdMApy8LaNj
O9ZTL1isY7TGTMTBkziniRtj4Vj6hr1DTSKBiFZHrCrvBuOVxkyF739Z8PkSpcDFuCCriGMSQxvz
hG2eEE9gDS6JxAohECRMJQRmJkqtxtZTANGEbgFDV1UU53SGAvf8g53GRGpDtERtCl4lvJFijmBr
sDb8sdzAChVFimkCujOdjd3z5dZY4LwhEEgWMI+sOCanRrjFbqwSZp8xPeFeRRR6IZsFZfgDwufa
rtYXiVcG422BDV5vyzosc7e0qX1zupbySDKxkqUOcuCF6355cb0P/lHfMWtEGqO+hhKNjTuOD3GH
Lho1Lbs/xQgyJWcJAbKiCOcvUKoEC1BmchrwUgWJYq9E/78kSKX7rABn0XtuJTFcv6yHI+HuoK53
G8/gI5jAopQC7wXgZ4pL7vCyPGR9iK4U77adIZakuStrohCTY3dY4WhyE056MyIUwJXZzPYawkqN
0Xr0lWeFYZgW1OBCOCcAZHqCZkgEVH48RHPZ9v3K1ew/zOv/pfH1h+25194fi9O13FIpnpCnoQXV
EHHuTOD0rwEqk7+WA6082Ah6zAgc6XvL1YCNldkoeFbQ2UiYf9JuQkXNgbrtdXWvA/8ZFe+L3D5w
poQ4nbKDlLt0V3z8FSBtyks80gzMSQR9T0eSWKSGHdLj8fFAfKzuYQrIJaWWf0gx0RlhxRoCKUzo
CXwXzOBTkMKdwfL1F2KltEmtcBAOn0Q+R2IzsrT/r+EYMxYqHFCrH8XVMz7Ge+zQ1Il2vw5Dzjzz
TNyLF9OAhZNBVTMgh2gPimVMvbBekm9V38lVNeT93KvGinAgsI5tPmRhLrvZd7+GCSrsguPmNQ+H
1b7tj+z+hos4IyMwCizeTZ+8u4dM+vSdW7RlvItSPLc9fs7T4qNBhKfK/CfkLavPfOhJW0X6TuhK
hRKoQ3xcPeztQILrN7C2pqafXUB+RVpoCNLsI+7c6RIiOU3MxRyQALsglvNvndjA94ATmuMXtbgH
ZIpyEuO1n4hdjLxvRKPZYlgw4DOIGsTZ2QlCL4pONFw7BQYoPd5lJpPpUNWNPEcGpfN/vz6OH0WY
W2DG9Fgqe+xGtuyUmLsTP4Lz7owKE8QGmuzLJnDLxMr/Lu09YPiBJ+RlUFwwQN4x+KnUK1w0596J
VlqHGCyTrh/pYgC5iA7lIts//fKINMFmlZgFOfDNO0/rO7Lrusl/e976PXoSewgEhlZ8qiqQ9CCa
lfZzZO9+71KW1ZN87nmBkgNB7tIaH31rdGBn434oVuBbnmrVIl1M+IT4ebYr/al9cr0C4xXljK8W
xOiNWFrzNK7L6HrWH7dcqp1ceddJoBq5XHLbrY3w+iCynLJtVIb6thbKtNrXkV4F8rKpxWar2/bj
PD0CHlAPH45f6AzbMv20Lo+fFcRGWIC1Z+w=
`protect end_protected

