

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Aeow6Dar+wPwyCuZ3CpouVllPxC4llA1Ukm5brPkUf6jbA6jqKC6lQwebzsMw19h5bccH9idRwDY
jemL0fBrsQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fhH+aqlEoKE+JZq9qghNfSjPHdRv5hlwG+33iOnHAwoQz3JLEXCjbjK+/OkJ0VZ47mEYRGFh4AMB
Kd5bYAsHBVfJU7e93cOCmqMi6q1NZ1B4TYSa9cbXieENl3lcMAWDjVXehJfBz/WX6Dwe2sYVqHas
VIMFb+sNilgPS6HDJY8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XK10objy6h7oUNp7hJFakI8VyHyBjdmYLutHMeS7A+cEBZkpecVT07LulHHgQ6KKziOF+tKEi8wJ
SseDgde3hi0l4iPQkOV10LTfLrRvJhBfeIZ8giQp1t0SrhVy6N2SSqAn2eht9NkZHhhTN2ptQWFp
0WxnKaCc1sV3GIghFpbS5rrPhG5y92GuyT5FWa/h5Ldzc5bI7CyoJ9vYfzMq58minDKJ0Jm4Y+wp
yHLZA+Ov0xHxm9GrfwhCkATL3ruMGZYQt2s5zV4QI9wQ2UIEz+JYy8mzm4GwHollMtB5NRf5scWn
l79oM70wWXF4vtffYUC8HG3KNp96Na4QKpBYPQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ykye4tSzDCZpeQ8JRXb0ob3ATquwfCaSG/ly4GVsy4bD2TWi/SlkZna7zRiLnZAzCamGizuqrWRL
lhFyzoZ23CkJDaAHrP4R0DVjNPCXgacmijI2x8zSxwjKptfeusObi+G4cJ4ea9XYuXHdvqkbssiN
HQHbZSHeJPlG8zIt/vw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j5byzLdNMnEoE5qwywfZ7XMWUUDa/vRU12ws0qpEN4GtoTZgc2FboDnnBkgSUXUolpwgKX2KPVWw
P1VJmwcR15FUwZQrqh9sbS63mL7WHPSLNYElbx4uy534LVuKyABLlnHKjoHmVUtp/4E0ZuLGoImt
/zsHn4GgLIE+tuBcZ3jTd5dxjmeQWJivwwjH/wFwCAVczK+9bLnUfJbXp5EAOTA495Anp3M7uHef
CqLawyLHuTbCQrqf9W/UvFrFP4vYRwsEsllUJ8mnvN8qELVwvhBehS0LrP1gDGa4Rus4OZzQgGv3
gxc6OKVuHGv/NA5wtcEC907wTYphLFlAs3rhjw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
1nCdOUl5Ydufa4PWbHbKN5gEkDRDujZTCw9Wc9j52Qz4ntlR7Eq9V7C2+aKKsETXybbk9lwWZGfW
5tP8Ef7776PQ467zDcOfXfrOhR8KUL+xP1AnYGyQRTOqv7ZDE7LLuCV6XxkZ1lb1WqDk11a8451P
+EpLOtCM8q7uz0iYLTSB17NKlEwDv7sOKX6gpwiTTI9VRjMu8pAGI7bi8pX2NZe433pmyHF1FEyu
1GNqToSEwz7UgoMdq23TrPn+7fyFmSMl7N2TlgzrhZinh8Cezw7y0aGjO+dxSODixhJUpFOOVUPB
SvXRvE8ttUWS89DolLE8aX57M0UHjtxbRq/Ol2OVouf/EpOwDzAoMjJLOZKcJSKpAaY33UcdcvaA
YFV+8M5ZNbtFHPIGhGAq+PBOu4x93tRH8CI/fGqvMvjHaeNbDh3/tsvL/aDYjU59DxrbYbm5ZA9A
lKrxBNaaxe2XB5RzXxiI1m/n7Yx6G2CO2EbkKRaLgqZXjYNUGRfug/rtUlNXm+FOTxA5hNwwVY4J
Ph3uAmGYly8Zf4cqwoFc7Xb3R+8FlzFuCtdsTj0rngASUXogVgP8rakSqsvg/+SSvp3t4wI2kKm2
mgHK3Z1tEB0tv8QYnWyjY9g6pGHBNx0ECjtNGgW21zIaKiXk5E1w7wXriFIZPkvY1Nx2ZRufrN0J
HrpZTSW0rWfHiP39yz0sIcMLqFqiTsyP+epeCwjOC4O6oC0BpZitgg0l98BjX5bQxTA78dr/OTTC
pGrUN6Mevp8fEf+yzk0o9wTrmynuQdcT7aFwm9cSYimuiSUTs/1sv16zXANrdUAGRN9UrZiTUMWG
WLb5PnpkltsfdBAs85eU6+HWWJehi1uVu6WljOkqKAno1b+7Prx3trYsdhwi7lSMfYd7szPBQ6w3
dmEpTWD+XsJ5GTdxoH8I9kAB4RiUCAhdSTFDYxhfEUQqbM/TujJfZlHMhsvRxrUUJpAVAB+gLype
BAfX8AEuSZuCia3UJbDr6qA5jhz9fmV1UBf27ZirfKHCO5jz5140rm5PAEev97MtDe/LamaJZaQv
Nqrovqb1J6bYuoFm4I9ItNAqmBbZRyYgvQsnbiQOSbqj+ahgttSR25/Ndi5OfM0Wvr3UrS4AE83m
tshxNoMsv+rUCLxlru1va13P9yycww4PRpxdc892W+AHJic9SgRkLaLSY31FJSAjcYUp/oTXy2uR
/cioHfbM/F2l7wEejwGxVl2u+95WujIrkN/wz6hnxsR2mcDXdjvQriGGhHtM9HUMbqmodK+qEFiK
54ueqMnrvtZmJxt6GDDFeP7BMgEp6S5u7awRdUUqSqfDhYB0OwfMA+2/g/IoAb1BDs1/pwv1nFDB
q/DTfZ6dMLRjEn2ii9cgOLPdImpTvWmJXqwgc5d/wvTh8/F03ZZkGBxv2EZZgTGANPEl2YGoOs3l
9ZADKaKgsrhXx5UDTYHhHqNucPCsUGZDl45qwFAnK+2oPtN9/KWw0hrKdnZ+tOxuX37BbaEm9lpl
STo5Wsx6HZerVo+fQj2Vr9elv3zNkIaEZL6l9RIqCRi++U9ES/FGJh2vLTL+OVyco4zDgyl6Dq/T
yfiQHhDHy4mE/y0bcb0UI3LPXd9Rs7UroNqCTOcr/ppR9NMqZEKp4tGSi22iOSlionoaHBxFMLsB
Pw82TJivEAIgTdsXac4aua570NSSNjDBpa6hlV3PdjV4hsXBSYpWvPfWY7W/r1gaWNy/zrgYaKUY
I7RxS/qWj79pl7fg51ePBki8zAzP1Z6Z60fT/0zwDkHJMXprg0jSv8y1XQeqLQ2/cgV7rfGdu4BR
LYrDYBhWHyN7wOiN6TGjlhdvHKvb8EE9RODV5tCM/NM6nfcfYgXpYxHL8xdy7+iu2Oi+qo1swIIG
/6Xcg2XyD3FHF3o46EwozDFfF6S95O2X4JQSy+1LbTmua/fSg1SopbvXhUBWaN3WA1Vnzq0Z7NpM
hYP/eeI+NxyelkVdukpRx86DJYBXbJuDWd1GIcoqHIDriXV4UYe5QKVobhyBoop53xoz8Dn3n2wM
BsgA5EwUzVbt6Tf/egEQgBdY0yYFOkS3uueVirSxvGbSyWrY2zVmw1QHJTqJ+v8ra7bJ79va82hK
JasywprW8ccdE9p2OjPzbKOT35UAhYNOhsFkzq4THQTyl4bC65Vyhr07/PVZkGJB6kzoRD/dfQUW
MqxpWjB0o3X451ovNcDxxHyMWVfejXJ71w3kNswcYI3ofbXclZvuVx9+mOMK5qMl+bMIzO6eYjCw
Cq22fzMNIZnpvswThyfIJUrmEaqqGcR4+heqP4oZyQljmAEnk1pz2MOOS0wlFNib0E1AezFt69R1
nzMRvIiR7+K1xYrKaq4epCv9AHq8dGE2BZDVFqSMgA385qJFwQ3mJ4aPSWphbQovby9xnb9coNNH
KDEl4lg4bh8PZEBdDfN8IGx1SKgZUg66eiVMhejLGeBKfmLyygyPhQ5dV+oeupTshzPPuidho+YN
LyLcAdVv+fMqflN1S7hpIqoAQUb1y+rOE9RY59AopMyfNqphwXv5QfmQHaxfoLsxwALFoIZzKPx4
dVYQ0EJ+eD7NUImVdy41vpo4849C9IZ+jPUnlKKsbVK7n++pDd2uGRWzgYm6xPsh8ZAvA/5tSbsM
VWhtN3+q6y29d4iE06/pbZaYL+AZNsR9rBqsGKoF//o5IWMLiYUpu/7Ayi0DPpsncGFyEuHtxMJu
deCvOzFNRtIiy11Wes3gswF9xlYDiFfX245ui6k4voGrhkz9QkToj6MHDb0PobYI9qi666KdZho8
r4p6fRAxH27YfE5dx4bxL5tBlv4SluuZFhxKI1ajLp7jS0kA4Pog/suUT4T5nC+5VoEpDwRABX6O
rV04mfnwM+p3RpsUcfOsU+MQEnmwJOTTcduBC2aphFAaomE18+837cI2QIZw+Hgc/JGR+846g2BW
uUnkRTyDZIIQl9g3ti2lnnH1MP0/RqsFVSOP06+1b2SPbVm1ifbyFIQuwtd9CdkwCSjJWkWi9xdV
VF0u6QZXjw5a9hUG7yOA/UvevLy5UuhCso1h+/JtxSFKTV2Ezk+S8gv7qXxx38IqdDOsLDTOnCrh
AX/OneX79b/VPcXVJqTIT/lBqHkqUTwdyRidyi8BEARKHSWb8NSEn5V1651wrrQw8TzIgh9vZPxb
vfKotMXVSdQ2Ivwp33eExgI6++NDrniZHAuIq0AkrY1zcp4nvf1q9qXhr55pJ7dlS5cXy/YuJ4Ze
hjE4JBQKCGpjAOhsuAZq4MF6M66GWaGJPLfAPgRqyFiSGDtHrSx+E5RU6mf0kbO+/bUjSHJrUISW
sNjlf+GSfiKTiHg3VN6GRVZh4ovj+u5yZz4348DPG+g/BURNRar6Y+kWgZ//aYS9upJDvH+oPQQB
yAxw0+4NoAwHyiCHGa2jBqZ2NWNgWUMtzAnFFGdauYuTlPgS8h4u3aTG4qTk3K8KFWqX2pv84hK5
W385VG5xiKwAt5YSSppd1T4OxScMau+UuDhWmpKMfmIMA4S7B3S+e57FrTZjhGdLXcKV3eW7G9Le
cxF9WdmYpIChj8i9yHdJuR5Hqm8LIO+ljjIh6UN3dimxPsuqvRhVRUqv8AmgeIMN3JneLJXhJbAQ
Ii/X2PbvRrxwFYuRlYzbuUAzc53wi2WO2GyuDCweE938FFc4cxewy9aPs20AfvAdff2JXNx8Hhhk
Lk6c+XNEYGUx8TpSStGtUULRURiZs/7b1+P3rAyJsvq3jHd1F0n3pbsQoVhhgJEAs/KMJHoJecUV
eTlfb62C6aQYJYgd2idZ0Kn/0K8IIBuXUIv5KAVA7j+uExfw/ZCbGzb8IRbbqvUMs34aVpS8vqMS
KYl6weWvpYxbHF/BF0T7nZS3omz7d6ceIj+PlFH4MwnWjOUCdV3afIyi0r0e9gVdp8jQULapCxr+
zIqFeHQdxolXOzkbhSejSHyHu/7Y1IWVqD8uEZNRdHIsmTo3w2sNhbagdGkcoTlwa1+Ze+3xqaHl
tb67muK0IchvHcdi0+zK0Xy8E8L/cJfzXabHfQBztm8pivUzsDuu8Zvz75QyNn+v/6lz306Hk9S+
bR99DtDBTdYe5CF4q9d5e/IvnRE1JIpNpNbKj73ZL5wwEfx3oC3KuAIK3ayZKEHPnFlfgf2Akbg0
hJiirLrhPzP2n+QO4csn/jTWO97aGpf0kVu4OuUyFEVWzTFitmcOyNpHIgYX4Ku+YFZ20VM/4Fv8
6/Yqr4fx53EzEfTRYLUDnsD8192FeXJRFCEWGKh/e2z2WiCOaoCbUJDnD6W6MGKDGY/LzRbNdtAD
LEqG01Y/FdTpJx/qKb29bDG9qzkDIfQWc0GId85EgT632caanx6rHrd5Zj2JcpaQKVtigvPDViW4
4BWLQbr9UbymfAkWgLqa5nSNF675D5/0nH8KpwT4ziqF0ku+VRr2GBlECpo8M+wKUzw37vPe4Tww
FVDqSuZpx5aeVcGbjUo614hnr/QIaolWC2kBI4PPuKLtiELNszvI+uXLPsr9f02LC9ygqafXjPpF
e0ZljuMQf/qUIAop7Fh04RWd5efofrYU7ZEtb67FrP9Bu1vgsy1sZU3VTc66Fx6/DqZqYod/rdQm
EnvsQqykpm8H2StQKIvTN8uFGYHbCRC2axE/N/T7LSZyjdmaYg5DoEoGa7WxCIQ6tI5FH03C/EAU
cYkZj+TkYHXy1HPsywvAts61ks3/mkxNVd5XEccK+CjMHLVAk90MSzyZ11oNR/HWDJJ5Elxx2BrJ
t+aDE+AflgNJJ7VYtXa3G7wTCcCw0l5Lj1auvLm9imeZjPK29ljYsAx1H6S3bQBKMMhparM8i+ni
SzwaM98m9zWP0cXX7DnKU/Ci/nC/huyUaeT25CPtXyMKj5r9pcwrfekAoc/ZD0zqYE6Cv0c4+ER+
R9Cc3h/7wThdvajCHkS5f0loHoRDq4XBRPeoM3TgiwuL0Qq6Fh3Puh1tcTm5PbvWGg26y4JI7Wq/
2ASujX1ThM4sWVbf8Qa9lnWz0L7RkP4JCnAuoOXAJijPGebUO7S3FqJ9pTT56RCECRuoY9dy1Hy5
HsZ0kUuzd1wlvzI1WqtgnKiXwp3sypR4xJLtF3KssqM/3Sw2qhz80EJr2EXbvmGmiNFmDyMAnujQ
VPnRrUYuUncCSxHc8UhwkFLg19DDlATCiiMPKbbHPROtrQb8sO/LMOIx1cxrxihAnTlWVnbo0PFM
tZhm5R4AjhnvDV10kHkofpXgLCLk6EmTuKJ8VrRHptP6z6if6m3v57ZxIXkuTI4rp35tt/6/Qn3H
mgzh8eefflsRti1MAOkNpNux0aQjb9sWjfwLgGvygCs6KUOwoLwRgFOvpLOkQhnDB4JVYxsKic9O
c5TDZ2Ahrqqlrt3u09SO3J2zkfMjD4oTZ6htUOzeOUVR07TNMrla4gQXtqngSS9lEQH7P1y6wtHE
+c3lyPaPH6MZdmUSWO8KF9Y9KxmoItXCKVLBtFKXBK4B29UKyOTOPmwrKwE2SrGUdkUOBmKupIRd
Z46x3KHZo/pmsAPh08sAkygAyYwHmN5T2ETmBSp4smmG0hArs2vC0vk8qxvtdNsRXE1djPJNpTZ2
3UxNSiIwZR8shKYFP8d/ilhzOrNVQElbo7+KT34lpjwKSTl5FQB6hBWnz1PkjxX7c37+TVfdhz1L
T/lqNoEO3cgjEdR49+UwKVe4DEMQdVsdSYWdDxXAKzlQxi1WOcNOVMPn46E7aGvLwSDgDA2AREHY
vhUnJeO3tLd8djoIsYmYS2OJizwo7XF6VB8ORl+ew3RZr3nMwQAbZp7bTJDqHAJ5N+p0MAbclA3q
ocmOi0mkTbXLMf9raCI87RYMx7pUOBAIsO2I0VE2ViVqRZ35UDWVH6yAYyzO30UyGGZFWtdCKuCE
40G9CmrzZvYKavopxzQGvKsTWpafNyutLVEZCLaG5RaJTXqC9opkp/3fNgXNWLvNwNCpN8xlE399
YaMRvSW0wI7Z9YpMakrf0JUGqy80D9pJQuaZBihlx10lhEkmt+zivDPbVAtEeK7g2hVk0Tk03Z9V
Y21feReRSWA81/z/9iN3joZ7LTxl77NzOed75XpcVnIWYLqvOeI6MQ2K+5jdNmRXCw5AJzeNeObn
XXihQAzfJL0ccBBAUleSExIcxQoSS9v3duSLJpvmxWfSFMUeTUTVRNHnxvWEw0Epd8bpzrdqJVz6
kvp59zejb8QMTMGwIAzedzYPfZ5Z1SCVaYK5gvyWgS8EJThO5SAf1y/UEpPvppBJS1ZVAD9wh08r
iUO3sdpVnVThJyoTzgaRYHKVxFC7iXR41DtTrATxudfiK+AyeKHJ+iqiPmN4aoEGQqRsxLQZvwIL
OBGbwZ81FOPjs548brANZmGyuIlOi0mSLL/XhIWf7UotMKiNGxeE9ScpJ/YybV8Hl5qR1HZ1Kvbz
HXgzEWGqRISXT+5KmZ27B83wKrI32SqxaY7rtywsxy86X2IpqdZSPb6+Ufr6Qtiwc67Nrhb9ANhB
t6oeAHVjPlt/hN3x1YF/BgaxC0ERcwCBT/kmq5+6PBpte7YZE9GDogWgep8g2FJelcPZhrxBDo/d
X5HQF0cSu/Nu8u1i7YjOfxY6yK39W4M9dyyP/4+oJ2/shJQ9tfvSXtPSwsYruiJuuT0gHtnr7wq0
ZcvVrcojmoPtG2ND4fRDZcma47xUJ2vFsT3c/4yb7MtUJYaowRXsGkqtZb1WvB0TtY0Pwg2SrsYy
awUPcDukeENIOwJHXO7cmq1KQzQ2Daa7bZnKOclQSr/ndOs8yS2KOQN7u25w+H9hSTutVYXNAiBF
cnZhGD8lpXSXWYHL14qm0jL6BQVidj6YLIYvJ7rKB5oQYt6JeklLgyHnyMKKDYKpMNJVmiJHAs/3
VkELS4oWT2d6lEEwkTTlM/UirCeKzG8vNY6GCxGv52mssWgscK3x9ZoN1MeQfmXQk9OSFUlIp0Oi
crmx0JoI8JsXPQIQdiKBRdzJanbetwzjZUvowATO5MS+/4IQM07z1lIPiMzDIdoLy68VyBkwDmqq
LZe5T9kpj2GO8rc1IfR0OJi8C4S4hQKv1o0YG/RP6lRtmAmixJQFUyMWP6aaE3sgjTioezEL5uDv
cZIS2rWFtoId51NdweArNVh2koke26e2eZB8eYRBqQOvLigQslSeK8hZdTe/hjAoFYddjowG6gGR
WVzsiBAkDdqyWdMQlqRFW4gPFC9cYdnGYiEcQ9ljyG6PdH75RAIClw9JevamLTNYkVc/MFz6aY/Z
AIPolud60LQYV6yJGuhAojVwIFLXc4uzkYlPLoF9xdXvQBh3QXUwqk9qrkwP2bGNP7U3f2N7m/IY
3rV+huOuTPCRB0GOFIngIpTSqTuBYNsdRhOADcyBL2uXDlSMHcygoHTLKUens2cSCrutG8ZqoXil
0t1Skl+pPzizAiT6TlrWcYae+PHVsllV4852REAeRWiaANNINaKrH9edR4XxmQm9OrkK1bj8cYC5
K+s+69IXqZrdE1rcqvOJuS/Y21mbcrHGx0yZGmdKsD6vvnbbkkPP+siyfvogQV9RsQXnPsoWK2g1
ipcjJLqToTl/fm6YYnwVaEz/TKC/v/SIYNHLqhfudZSLbQwqgI6MzTQJxYIQqDBvW/qN7v64fxE9
c3nbWPFwCv7d2u4Uyll1NSjr1P74D66IwPCrXurK1sTulkQBuV+aMDhIZw8zWzbD5+poI4NtE04f
DC6A1O/6IOEdgibXZLyxSzuUN6PVoaLs+vwV4QWf0bJkMw2/y9ERpvi23fZxGowp2cyN9Z3kp0cx
G3VzPEKsp3P67BXvWzjD0J0u7i5zXiE6noO2KIj0S8zSUohK3T775IGJw7hBEvwm1/vq99HlV+lY
Nwl3IE2OSFoNoY5Io9yi7iYZ+khSnBu2rZlvQb73mXmCz48J2Cn5brOXm2ambXqAqfWsH5RT0yeT
ZozkqwXadWM0MMcygp1AOkjuIaHZGgOvD9d2FvOufI/ragkZxp2/R+jcCKyVuQG6Vfavygok2oLL
pDsTgRNUpWXD0FEmic4JRYaB9muloIXqMAOF9yANlbiwgDiRSHbh+DFaoqK+F1rC7N4atNLL64dL
cufq+foyau/sGpTIglfTiJycnkmjXeZZqWtmNSCuImkrfveAX+VZ/gNoGf+ArpqNG8uGvt3WfYmS
uehLJU+eZiEXl5A47ahk7a4iS3EDCgIVIog+r5vvXXHecDp64vvEiO3xsf4+DzR+UgkM98/kW+TB
JJV1edkwKT37iqK3B8KEwfh8zh8nUPDfGupZo8sR2VhJVg4E6l9lruJBk9ZGbVpoybv2+Dxc2tCp
K/rmU6zGyPAH5Hz8Yq5K8YFjtzpZn+KeecR50jhsbQs9vKatkX2ddSp1w/BM0/qT/Gf6HwfM6YPh
xfzDpKNOXc1tkMaHKgxF3oiRBMU+YqaPF7SL6/UuSkuwTKwuHFCResZQ+LXC72tlE8REqEuSAz/C
WyzwS8GgzezH1QhzONfftyXn7+wMgmgkE4hq9Sjt/WozzmGTG78qlYf1BoQ2daQqQQJ6T9WWra+z
wBzM+oVkSIEo5adOV470+EGX5m88HFYXiQKeBEiMbvTybGC7/JEFx9TH4VXZf3nE7fpUw4zsktQW
zwDSsVTl/9Q+k1ARcSdcemAsC5EmFzVGk3K/fb8jo/axV/QdjjCyHvmz5qOuCAuEgSJzxdMGIoHw
Fa+PcN4JL3/a+Rsh/WvzI6uKZCL6/OsHnRf3OX9gSVUff5Wy+BTkKumCfewGpW4U4aGZzQSxPy0G
g8svyd5nYpqw8qU0V179vdgyUgsgwWzlTqHM9zdbU+YDhm0S54KOMCTV/+RGycFIjgzVENDUpKzq
xITNCDEwr3kpzbdM04UyK5D0EgjiLQtzDVrIW6VLTyEYfnP4oz0+8Hxtt+bwGzBqplqR4HMIHTaz
mbpxwiNMl9dGRxlcSufEef61OPZenlOf5NTcRyHGTl23V30utjqqT2qoZEa5c656oFHN1o8peZjw
MvTkX5grXdeHxJomAjh0NkPw9+WKvja1FHnIvrsyvtabyJGSzu5yi5I2HZ948FP8/uy7xLYzIfM/
5ynkGTVHTMve8N69W4gzSPqGhg3EYiLhTD2nw5EMv3y4FkzTU84lQKmalcIA9ctrMFdAb5w8zMV3
oNOZckwnpLr8+NIY+BXd5y3sdRKaaD6gJt3U19Wqyt4SacnuZ1risBVsRghPX3LLRb++w5bZF4sZ
YsPDRMbit9gN1lmC2yWEe0fDZepjQQdTGWjI28vaaieYpkBzLETnHrvCGFhXYrVCqvAhLq2dNaPD
59np/gwJ9XcMbDgbrhyAV2++dLCdxfR4Z6j/EutL4ecV4LHGKQR0Y4ISL8U49ramXxDKKUGL/kfq
MQij5q2cL1vu5ov6SyMj3Ah4VBUgCXFszxGlfeJOt2k+1q+d9NhBZ4VPakbCVvu6RNpe1gdUB64b
VDNcGykKplGyWqCHr2JwsCO3wQGR9kyeCkJmEgpOtVrT9wJTk2MsVvP28qWTn3qnAcEGTAO1ozeB
GZBITv4uSXCBp2fcPvqDwP3WfruQTrQ/Bloz1KVpBOVrKFMXU+o1ufHJop4BZUCR8FZ/k6iZBYIm
52GxdmsFJuAP+hQ6YYmSxnSqTi/jokQv6pAXwPm06fWfER4uujnG6PO+EO45Q3gJE3kq+kUVlIj2
1b/r/gEVzDTO903cDN+vKv9wyl15VQ5+ISvHAd23tL/NLhaPPpQFIthod4PyXRBOUWXfgxXUh4Wv
/GZpLenHFUwd+4oYzmszyANJuW0KTRnjDkvDGw7Ew5GgnZQpGIRVqclIfvGT+EEvjCR5dHhks9zJ
pm/GTpORe5SISdYLw8F4bmpB3N/EnHGAw+a5rXkpVkAwubH877v0+VFCoRcgq0Q73DRYNXJg8rEp
g/Plmx4vmsjATdzfp7BTg68lt3q40a5lNbf3c6iwqk3zsyqk583yqcVkJ4I3s+XBKrCLoRja9BrF
M5zPsrLz0glQxUUHWjWXBdfG+vw4mrXVZXucGIIpGeBiTuMGTBi1WsglkP/VG+ow1a7UHShhXEB1
gxt2ZcmRLbmFro7EY4BxyGALATTrrKOQe819TqRr+uksOvXXhlLVW1hBnQAGlTyglUv3S3WgfbIJ
i2z34V5fTJGnM6weo1BRAmm7YLl2Kytc3T7tEEhGxMTstIqrB9VJWnSxzeqSBFvQkpv7QkP9X/me
9CvI8HRBLAcCkS+ajH+Ac+NastjpxNHsJv/8t0TqcHGrw+TMWiOqjRN3fkP0hlBYuHW/vN7iwa2+
s52bHHwdatDE/WS0U9Ym1/oS+7MwI92ZpeOIKQ+bBznViQXAlVPHGSQ/O0Wp19Y1/2zWRBsTI+lM
PhDLMPZdtYa2liPaukdF7KxRBLpvkRwB3XP9WrhWxTMIsJqU1uox6nUvgMuPOIoGzxfoaFLOySH9
DXieFJWoYvMFqaSddNfrwk9rsohFEmjSo9rxpEv5RcSmTfkKeRzlM26MJht0hRtClmQtlSlfrCZU
J8Btt6E7aYu5QY1trXQCXAeWoG3D3rHJ1fzJYJS/kT6De7genwvLmoikn4o11FDhvWLaAvmj2skz
iKqgXY0xlnocUtEzsxVw3NY0VJfXpWSbLUp0ZorOrY7/BK/eCb5YIrwLalkxuuJatipr/srVkWCW
gyx9sN/BZ3ckqFDY0P52bQnOPM/PWfasbeYVNbGSGvvy8I/vFDzbdv4JNSwBPAnGZlD2bc+jZJJM
fDbbYCeU+Wm86d+axG+YMdyuZQPP2sSFq91YOsPioVtwSkF4r4GUVcfmZDeladWAhWev3XiWntp5
R7qvRadTPaEqLpUthwvsSjqOGEjfdoIQaR9V/uPKxF8vsVfGK3h3xdL7Dib75s+tcUqSqgZlIRBh
WDyHtgjA3MrAAnlSE7+Q03Udy0ITD7ZCKlEfNR5C6TNgUigjGvlWh2hyZal331RxHe9mS5nxeT/B
sKulI+iDD0x11oWwqEB39jpMtB/l/LDIyfN5i/eP22NtvSIj/yP27OltsaXzlWT8U+6T9wR8pXBs
7lmEguEk9C3PS4wO/0Y7DLSgN13gNtSYHWIfWk01o1Bwly6HUc7FUXleWdHLZTqekTPLFZt9MZ2N
DoR0aDYjOdViHp7IpPPXUiTLw4e5QGmRagF2c+ZTQpX1KcONGS4hjPKlVdgIAqRYulMJceK09yek
7h1gpbHhZ3zyPABlkjDbwuL/vt16fw6CGjGA7Mw/NdQkT4GHX7gH14Nvx+v1fava8WJ17Vk42/rY
rWFXgbm63QLdBbS0qUwfnKP+wF0/lX8G+RQ/qeLaxHRMGfH8Zk2diw1C+aqwfKisyjuUAXn+Dgru
cFy5T5TpIaIHIyyxAteK5x+0Rl4SaczEs/5f3XCvJdQ6V/CXZUioNf9Nay/Bf+iML/n2Y8Yo+GHI
cn1o0xZ5i65XPfkmCT3v+DNKXt+OkNV6uVAQvtTqiDXZ7NrOABnUBnxhnnOH5d9QHnHVB+VTasWY
zsdiqntsSn7LwIXgdQ7uGuYvjLK21TsjO2ry2VJdcemym4WjOWd0SXwQuUbKKieDVeV+CnggbWQa
wD9cMwDmvJodA5CGg7YVYpHTMpKU393qGpPvZ4+oKWO0r/NmOXtWcSVcHxS/1IK+OtvRSipOHULi
Jc9KhwkDofcpuf0GpHmmddy8sTomg4HDNI6fIhD84TMGlgzaSQJCFAusf/ms7P6Ez22j97uUJ3ja
joVvs37B6lvKBqUBGtyExWk6+jYSPZ3yxxa6y0szKcpeAZzJgDQRx+y2W4O2hpIERfbBoPALMlG4
GXB+CfMzN5+A0PwnesVytGUZWaiHrHNvnTVNjnGlqotfl3uVYBHnjcSs3602gvQk6NmwW0qyX3dl
ifgRLZodBH6P9nh0nhpPPsG9BiyIr/T6POUx/VNDoUu9Y/q2/E+FsDq1Y3w0se4roEEtscBsf8sG
PYJ9Akz2ccLXORRHXZl4jolu+fDO0d5GI+8dQ5I904+ES+NmPd0h0rS0G33NlETBlk20Le3J+F8g
RcvMCFuORVM9vXIWkAbcydMaiPHtUIsIC5mWFD9p4DGm3JnOCYB9yVsa5z1Kx87zJKQr+dOWHrS3
QjGYCcWcjTh+ORg6aubIg/0fMG0hzk9M5s4cZTu23mmErcwG/6cfbSeL70J9ZK9Kdmy/DLoIfhY3
XV8i9fjRp6ZcOrQqMuUPJUbRWwRSs/NDmWrpfVV+GKqjrSDmOyIgpHdx4fp7rqgEAoSoPlZ0z5h4
eKP+ICv/xkz4+ymcFM5aaPgnjsczAL8hcpz+dqP5MPOhhyQtO1lrpVGlBJtPdnD/EUzNtNAAk//8
276pZoGImdQPkpAZeIgRKc85NZxJXYO6jaL+KLbpbWzqOAqWELhGPMsa9xpihFIk7/3HG0X5WHSl
mgsyECCKhbx3+sNLmX5e86NuTHdDeuuCsZXRIl8lwuDXdLT4cTIQlpIRAsX2Q6z7vgzgWffuHnAH
FYRwLhy4C9IkRb2izWLWFwbv9o6itG+lmpUU0dR7nJroZL3pghvL3BY4IBN4f+0Wg11y9SnwC4v0
RKooWU/YILxhYPSk6ICoNFK2yTVirnmpJBT1N5k2t3chQz8rSeBDmCdeRFFnuAFKq9ycDeSXr/5W
x+pHuG6tft+Rs8a/H9hLj2MSpBA88QW9xq/Cu9XqpABmnQml+wTlRQMG8j3X8y5g3MkRCTU/BM1T
PuqjvChN/n5VsDs6O0Fx59zr/sSquMaXRQ8s7Mwif0QvhRNNHO5dKXoaDX3iZuEsd+ZqwulOTJ5X
ZqeR6Y+URxPab6eVHRvhZBE0YQxoRWEFXHFeh6M9FkkMkeqp4FUdaEKVnFB8jOTQBHRasvMowHeY
VJmvUt0QD6MzOPWGyPHG50QX6ZAaD/Ol3zpODQ2KxyftGUqB4VoOyg/xMOypXJUyw9IRTP5FRrxY
833opAsQzxayccNwMJ1JaaRrTRt7CDIaLLOCGLfeqM8xA4Hok7q6uGeYQTTFpAxIC/DoPATSwX04
3iKXNXZh8xOhLF6K6t+cmcLWAjbO4GNiwQ8qD+E/2p476d7kZuOf6il9JbKk6S2RS6+4Gjj1ejv3
wSVZaLP+f6Ae3sqrbFdKhD78pyB68JgoPSrjglR4UOebZYLS+RFVcHsqdDvd1Mtk3uYo2Ce4VI7y
wKoF9tYHDRtKHwYI82TQ+MGNn+8pYw+UNSyTWBtLCh5L97k8PM8EEca0ylD1iTFNpdwbJa5GpztK
VpplCem5Pqt/gNR26UxcAsugU5OuO/NCdAMYuJw/cTTKOE5QPZp7lC1NOtMnukJG6F8SRnil7H1R
hlfB9N6DVYxVS0L3VqyDVRJpU8BUqQQ2pYsrvjhgTPNG419U2ILWlLs+W1UUIwmazl7qrdP9Odgv
wGjiWVIwXaChdm9dtpabyZsrIhXo/CoM6GNONu/5+Zl5gkVfvqPTZT0li5YltiZ5aQFkk53v0uIy
io2Knsp2yPeeJz2Hy78jAMvR9wPKsHb1JNAv66um7EMW+F4irYZ6mlO0yi5vTaZoaSP3phsotLMj
zkEZsEOv2hYXGC2Z5viguLFtsds/IRFr20Wz6pbMeqmaFy/AffetpVvYZRMLjqBdFdZUzffOw9Zt
kinTNWlQXj0sxYlflkyXMHq6/zyLxspw2MiGSzih4zoY+Px945sVMjAvx/eWg+WIHHfvZyxjkBrA
ZVj82GHPNqY+VyVeRaSyER/udz/44oc4zBPXAps1oxLN/JdYyTVdiA7KA9adICHeuzH6HGZm1SVg
Ct558eseyyU6HPJdawA3SQnwyYxoCoZVwITriH32WDJtp87NnpM1G6kt1h/JTZs6bW1VA0GsFjOU
1VkQ4lCotCnEVNlBq9u0QOYhwKZLIreuk1mtxv7ApYudivcPzl/MTk0uFvLZr3W34DTYozaMZJA/
yWTWkEgof5JL5br5EVoi9Bh3yuY1v+1bt0avz1RqBd4B6izFlEKq+e2gr8UIiLrYHX3PSTGirm74
Kj/9kNwzWFaaXfjIXmnSgA1HcPaY1zg++VKh+WW9MfCyfjcvIo0LyhCU/dXEbCokNJF6oR3s6Q4Q
alWdLslrsWQR24z09Ca3rUX6o8RLFYZsufOlqjsEkRL4hCv6KYA=
`protect end_protected

