    parameter   LeafWidth = 32,         // in bits       
                PLBCapacity = 32768     // in bits