

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BLQaKZsH4asejKznGC3MqRlTiz7BcudfJJscBLiMA0xMqmZb2NnzsT/xLigT/CZ3d0+qNYyx/rny
eLoJ247NGA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OsLcopJPXayiJfcVLCnf1kmX3JIo+z3eHtfdMz43bjypBxd3CwO/tVcXGMc6dJmHdZ/Noymq2iTo
9GUwsW963Xk1NFWAofj748NTimVafVoo0sJKPFHpHucNbZIlYygAQkqAYe2yeBJlnSqZhs6gdR8W
25Zj0I9h9nbg3tDj6xU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l66+uTOPhXeiKCvyaah3L4u1ckedhS/MpJHzIp4T3afloSG40AKvW4LnkPr5xeQ6UxCDlUEr+5zR
vEA5uStVMU2GDpMAJqnSleinU0EQHBIsM0d8cyq3D8/gGjqB2O/kX7nkLMcxDdXrDcvPV4AKLSsw
6EVA7ivNjg3fNIqbu2+zHKSkhP18GnuvtvE7C8sxIfhRFzgWschVJD03Jz/3S8b3NL3L2A6DiXRT
jvBE7P01tf4ikbHHH8nlhvdJFVMrYH1VWPgU6wAEEjyfa4CcFcqM+5ONmD5OPnHblwvgdPcWKzsL
wfOByf8V5k9bmNYvNJWuYFlO362iV8DdFOKUAg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JIfbjaO/Nua5r44GtyHauPsGGypbV4w0opy1x4qFLvqSrDfVjJmq1LuT0i2ufdY+i9fb2XxqQckE
4p12fYTQVYCk7DTHk3n09qxhrStTQ2hk8Me9Wxi8fgn4s4QsTXA0CspFzXnowgY2ZNmG6Mm5iOJh
fMtxhLDOBzJt2RuuxMg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DifpRpqTfEncZknfvKTMRJDfeJ8lK+rNN8XMz8NuSfhC/7MGMIyt1EZBQtB3/5z+4f+CPY25JEAP
kwaigZF0fTqe/vxUg0IwlCNsRUTvv/JiZ9c8q7gZSdWhkKEecrdKfmsY2tk52RPbTPaxLmK6fMoF
cW0SteGFpV9tXeEybrJKpX1RkRzdccS6EP2N0g0P1tMzZJil/fUxZxEsqH0F2jxYPmAMkf6BFxPf
iyy7U//d0VRAD8ceTvR7RQfjSyxiaj7FnbUWhB51lBtz/h9rWbAxscy4UA/ujxTMgl7Vrzz1vKwP
9KcAc3hX6JnriLlgDd+qVKOGU8Ojd3JfghCeWQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3584)
`protect data_block
p+joIfoh8iby+TwtBSHLKmQ4Sl6EOQzS+yimz99qHv9ZEnRVh7n0gXnkkyIa50tb/F4cZVT/fU0T
MLBwrhS4sq/SWkL+0cfuCwAthaoywbZExvoQeZ8UKDtQqlJzjnFAxvtWzKg//MkzMl0dWa3248gA
Vjwpe+8v9Ss31qZJaTW6n6e38fYerSf76QRB3GlU21tfApeHYz/0ES1cIFz9s9oCRDmlQNTLqRI7
hCy6JX+4XMDT8w6KpVH2xKDfAUcfuH9GYoS3TII8rKaf69BWDV/2lBb37F7/RsFDooAOED6Tel2p
r6xUDK6CA2gmpLnGkzD+qEhnA/NAtQxKgTUwhPYxP6WflLd2JshveBgYtSKjH+J12p9kgRYERZkS
HpAPHA0yqnf056U/KRxk/+i3ek8A5bFh/+3UsIXRV5Zf3S2VM79Pe+aHfScZL93ypeeimimJ6lLZ
lKXnSqhjGesWFOJYFAqRCtKtaair6meI3LB8VgO+8wwq5B9eojEUyZ1g7QJMaleDTW0vUxl4pxsI
cANQ/5W2eCrF4mlACyIk187Agbww7AxFE9uCiCgnHC25yfcj0f1DcFthH1f/dKqfoSQlyLin4ACY
bYBqxURDakKofg4HEah1eTjUb09jP64b8oKGN2FFOqUse1vGwACSX06ZTuAzw8sHteTljRlCm2fy
Vdis8n/9LZFGYUQsTUVW5mibW79N2rt0EoP3hXhzac13Ldu/zCrtn5Oc6CtNC+LEXY1iuREe0FCJ
qP0ifFvwfGjLGEif1ddNKUa0DTjzue9C/9fHzfLZ7rUn3qN1v1D5oKQWVlSLBEpNUCSh+HXmpJ6U
J6JmT1IeSVJwHlgFkdC8RQh3erTnqTp/noRTJZoIjIk9hooh9d8TNvC6+zZGaPDbrcygqAwvTN4F
6dP0z75KJnHLiNyk6wvcbGnB0vHtc51Ba2Y3hjLCxedPGaF1jwDd7vsaFLJps9dDy2TJxl2Y9A3S
WteVVCbG4SURl6cUt+YOpcSh1Ioh6az6xmKOHH0CeMJaYmnOuGWIeQ3ft6w9jrtG80TTPG/BqOA8
Kz/eZIIanEt5xRDnZpxatx3cfZkWmELCVy0QUylKOeHJueJO+IzDZNxKKMKRgnsc4cSsj74Vq2rA
3e8rNpObFgrUIBGR7JOgFiGno66sde9Hoy15rBrj6EN/lLcaNQsUTBN/71jnTpwfk1U11m00lF9D
EkWUaEV5X7uUkW4/1ZdAnOF8zASOgfnWUiROpwlE1h0ZQEkSl5PknXrZvdrArp9UhxQQwk3nLQOx
8sYdCkLQaaHTlVyuaDEoUmo7dq8dI/WSOPwvxCDvCjaL59X9kAXS+CKOzQAn9DeNKM5LkvqEssFy
zn/WgOoB7qW6IE+N6jRxZJQoUd/M9kU4jd4PTMxaiDqmL6PphacN7cbsqFUDPMplKw5zp2CvhycP
vrAe0H0RACe0iRJdBzHiiKA2HmjL0FLdoIWy6u9ggrUtkVeH66QjDs0MbJjRfYBu3Nu48zCXdnXm
d9lSsWCTVF456hxGTa7BxyoFRwmI15Ar1NZ8dvTnLywpbaIzg6MUB7lP0i1ip4m4XCo61bPGDSux
yLxKXf2Yemm+raqVNPduAybdqni/ZOReR11YKwfNlqMopDyKP8d+niT9VfQ1Ewj+8MGx6fsHlZe/
/0WnAOU1ql2cyFwvD9DddRw2Em423Bf4+K2GFAbWbwUSPHWFwoj4b1Fz3xfHdxxTlnDuFXaFAzst
CW8ik+VVQWzsu7mMFTkdVx3aGMqhroiYLnSRaxytooODcNZE2i3vKqlXZmOB/P1G1ZDyWG6MmfVa
vBJLlgXKiYRmR6YL2qZyTlRszR7elCbdMokmaKbi8YVqaQ0+5NwQ5XdylOwsu/h2XGlBrrf1Ryrv
50aJnACAK8EddK0+hleYJlq4W0bLOcSueFV96f+KxUUzC+H2PkqBrT1nztDsHzFzHlcNCPplzQ1K
xehlXdRG6kKT3gTpx9C4lo8X9VcnyDHtugvfIVJlaAXaRkoZOJlOqUZIH+qIXeeSiFAzS9gyB/kb
YT/oyRxNf6uQdf/9sMBNdlUvWnAetdQNUR5ydf6sazUwAnoyJuomDhl181dFLYj4GjJtVJoLLY6D
x9QSh38A65qtHIMF3SjRmaNhHXwxKIY42kiXrQeH/sK3orJP58GqB6d47fCXe+ums4gPRiwpJ4Jp
eedV2bdSrnrlZOmUixZuPqCzHMLp7cRlE4Rs30RqnnmPLHF3TaVLU+TQTahyoXI4Lxfn6OHXkEnQ
RvGRUEKpUW/bZiwr2+O8tEPAf42QVbuQSiovjhwfo2huPVU/itgtg+2cE2ZgX1dgN5TLCqiindsa
rQ/WKucN74IKChTpGihr3Kspb1Sq5XkoJcDps/lk816mel9o+p/UzFWttppBezGnozahzHPn6Cve
v8Ha6NKb04aE2SvV+l6HV5/j6u72d4IDFf3/E9YgNwoa2Tebqv8zxtxgR7W6Toi/39S/s2L8ci9+
5hwjhH385S/HTEQi8M1Ki6yawWgMh1RHHFPfiXn25CK/SBEZmW720ZSBqeLyZbMBHfW+kMnTsHJy
10meBoO7FmLTGxecjDDScZP3cJWumCwU7+LMYX423Ur25RvTlBA5dPy6tLP/rJR/5lxOJt7UuTCb
mux2//rxew8MKB7fMzxgziBjUAF5L3lWb5+eI1YHrkRCmmmCZVyIPxXIxJo4eDxdnt9+Rr8LqEA4
XxXhJfOEyhbrq8wbf85ACbC/Hdffucr+CWulXco88uBKjxUmVUuXPelgpIh9uXOPdVTRxrMM2BIe
ELDZPkTuVuVed358dXsgUkaajkAXdsvgLGuqIYy+3EyrmLjMomSBBCa+3YZ77gtU1kUbBN0NeR3g
8ywGmDWfY3z236g6uXPas19r0UhOWLMsxdEqD0TE3EU9TB7BRs1ZJWN4lYG20hRTQak3hEOvJHrS
uqQkKTI7jym0bBp3V0t2I7v088h6s8HjQ1BvrNIH3VC9MBRMHm7POJCwjazmNwSZW12l4RGaoQ5l
/vTAVBevLym29w1KtZ5LiqoOrtW4qKZ/Ocv/E6OhRx3gQbgD5xxo3x4wofLMNxeSfobPe95l7z8N
fxfkVRWdZ4bkbJD3PN1J7oi3zoipjS/jVrYSgaHn3ihVh6mz96u/9NZtNiekuulqpZToRJ6jaOdD
kSjbpJLv7HxhYmfakiwdsM0sPLJtjfsGxISMGOwa/rEF4tKxqqIcCQJdVPXV9Fr+JUtM0TS39pRY
b9Um3jtpZXN3WZERLg+qJO66fiUn6gSnzIetAHbo4QfEw8iKFb/tdHiDusdlMMpkkEmoXpbA8P8q
XdmJaz1WVMVT4bmas/tqEtU4caP8q4ZN7DogPKKPbgfN9pXuG6BpLgOf1XfxZ1JWL2WnWrjlbzkV
MQAKziOylgSM0XUr7V81sN+SANCNHSBRz2sM42A/ez8IFcYJSpRVnglNnMiDUFbZI+XVLvQl2edQ
0llCpY2JySapjlHTE0aAvV27JoPpFpkgCIvi6d9xxpe1qnOQ5n/Y4lfDwvBC69C1sAZ++b3ixtt/
WY2m5edKY6UnJz6Z+0icmX73OrkYZYcTJ711DoE8+PbJTMrrnfZ1mFoLolHaWM+ppISKrkW9emNo
8Phk/8J/47ezJeSoh1YshGwsr1RMXet0n3OvK4dN7cWyXVjzyTgxbF2hWC2zjOI7AoTpve3d0lbL
OFEkfV8CRM8Q4WnkOraCJJ1Gik4PEtqiYESJDFzTikfnlk+T9VOLoQ8PblkmCcidL7TfF4WxUWB0
hDd5Xu1Vx3J29+drYEk81pK4//VkEQGjLPqsTcp1Z2UkW9cjBZK5KSF1p9CxgAAITRIYRwfKzzEe
x+1f/6o+m/R06nhLOzH4C2t8L8oGqjcjpFA/q6IfWQbr6cXqKHXzJCYnMIUH0P3MrwuYoVqBNcG4
uxVQvlMQ6Ei5zZoYVOYtra3YA1hwMAusoMUjucDEjx8d1cqPJ1O4Disll+RvmnirDhWE1LPcASHK
WN9lmQ3h7WqMXHtIsurRMiKKAn8TlcC0mAcI4AolAfOkytwzi/IccUIfsqD7jUQZNZy/qM1OdCWf
O4ysLwQFuZfzap+yzmVadTbibmTT2B7CBJJeqxfKXDq2ULLBr62af79llJ7MAdH8rl/DhVQJSsWE
giuMjkECCnW3gVr3rJ9/zgFdACy+fcYjngA/annjI/uiI+RopMdotbeaAqkRe3na7oSWhUATUOBq
+iEm6ukEqoZP7sr8rniN8NnN4ohQ8UXoqbRflYb+bETuYGUiGOwM1X1n7UbV80kMURQNHTzXpajk
0vyK1KkQw3ch2lsq8WfMmWpn3Qe9UCBblw0IN3U+4RMTTp6WXRS9Vfz0DqOHODzObTOmh94lKa64
/EO39tv4zw4TjDU68Q87rm9k8KWuP9dZ3+j9P0dNm7UhuEAp4803XPXLk0HM0sWheveSYMCLvsmh
cVgCvUDYsMhzJjBvftRLJZrnFHAQehMORDPDdzqLiIBvdh32pNTa3BSNcw3WBALHT4DM/YXcAgyQ
SqHkP1EckZGNtp5pCHdXNWdll/s/WBng6nuNygK6gyYbs4ITCDjYZt/nSttevv1VhbzNhDA+tjwA
ifZVB8pG0DwNkBSz+qC8DEdWrcmt8m4bAfTGHZiC32Zq9V9Tp794b1nJU8FhLyYZZdoTgiJQaArB
aUtk6jlpfjuXtRYZrsq889F6tNCdrvaJpIAoJn9F0V0gPvXdVSbWr2A63s7n67N70Ug=
`protect end_protected

