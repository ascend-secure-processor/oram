
	parameter			ORAMB =					512,
						ORAMU =					32,
						ORAML =					32,
						ORAMZ =					2