
	// Sent by BackendInner and understood  by StashTop
	localparam					STCMDWidth =		2,
								STCMD_StartRead =	2'd0,
								STCMD_StartWrite =	2'd1,
								STCMD_Append =		2'd2;