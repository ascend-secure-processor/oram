

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NzFmjUD8XE+w/HVEVMfaU9nkNsJWEUWVUNbVxiK3QiEwiP/WmsdUvJ8Z6jnVm7jsbvSC/rMUaRet
3uaC4ntk6Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jYEf5kI4ImQZvrctQraRnaUgJPv0gSBqo/n5n+T6iwJIy22NQ3qViYqi8EHK5HEDhY3KFAL+XLqD
4x1trPAk7hTjgEVwSQ5IJCWv4AGN4BlbBba+2oHqWWt0F00+XCNnov+ahL6IDhEBrfN4mGSJuOr2
ccZdQVIQHm3JdUfFcqQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T30nECWqgr+bIRTvxuxwYCspGLIzFQA944zxoh2arkYtu2A3XXGhIxuAmc1sTJdbKigKmrCEVyth
OBAIAlMN7xNEhO+U8LYVspu4Jw/2WIiWS6Vnh90/2xyW3Y3Y+MyypHT8zcQLbu6os3MBxL8Jgwvf
xSJSrKRQfzQ+QrS6unidP/j51GQCFDhQw10sTvxDlnlqXT8aH6fCR78reGs2sMWiMKrywz5TIF3p
O3gihOjuNhZjeNYXoNkiYo3sr9Nx22k4cxy3/ENAmOTkyMgCJ1teRC5rqBeAwYTnFmmRBXbE4Pat
O8qDENLDrsKg4VNQ580tb1e6LM4Ant1nFHQwuA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ePJ0fef9vfpot5dvQD3hvTQw49srRBBiZ5iBY44CNqTSvNkUXzoICtyoorLMeCZsKzWZEku+nI7L
XyQ8mIi51EhBzEiukPYQBO3S7JV1l7oCucCb/YahoZF5BYd62j6mPGK588ql1xNEp/Tx3GRyZqcR
CD8Zac+/nGI1k5beFKw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nlAJ40uREisM97Yshfus7G8shucFbDE1pvTolpclmxI6y/Z8AhMhjK53m2fFJrmRoJBUou59alwE
OJLzGao1PVHRPPLspuGsJvn1QCRfvEGGRpVHjXqepUmjanUYTl9kIHYuJ9NyU9CMfxuMfji//j1T
5c2bOk251uAdoPVjNHauQUQyaAFw9lEHS+HcYrGDYlcTsSEThRkvZ9HvlzpiqgWYHJPd38bZC4Tt
GxVMtASEwS8FKiv6d17Ndy2M9jC0aLBoN/PYVnso1LD8flghCPRD9RuW8hV11NlqUbx42BCItefQ
wSbhXo1Z1iwVDqsDVvM5NceXT+bMUmMBEuvWMQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103856)
`protect data_block
qkQvY7T6VZEJCb8EPeHGDPDZ21UJyMVbgIwbRJEaEyJ/jFgImRruEL3FERYB/5cfz3frA/ixYP80
leyRXtjVB5Dt5tlIM6xUC5XPlZmgVnQRkNeQZePHbUTtJHe5uAnSCEjMSllo1xNbs2e8515w4UY7
lJNqIetxhPn3Vvm8qXufgVSqO3ifPi7bCu9atH5Wz4WXh8+Kl0uIH32Qr1YJEyXcGtEJObufG8wf
XLAaXWy3RNxmA9WtqaVoP0C1jLy9apFSpN87Ed+gdXrUzTCmQU+sbFY2uaqW5wZvg4kSobYRRPvE
wXfuoXbPeDLwanvyAbNyEm1N4O07U5OhhZqB6c9vXPACm7f4AaKRlNL9SX2pY5K3IxxebLGyA/Ze
ZsXy2kkGN1F6zEvc2gNPz2MmGUxZEOvytTmwKAptm3WTaLDDDbpG+FGSYeL8uA/GctRuX/+YAsex
saqlaJy+eY8gf1Aci4XuDjCBKLiLAws8v8bBWsWQbdp7JDu/GuCcgN+iHd8pDuNaVcZDYNBOsSyK
OfRZV/bppKSJywfeJx8rEMKGdQ+zbHT6VXiNKqx1WbS23nKTSa/6r4az6J2GxdvLNm+GEXI7aByk
3klVNvMjBulN62QSVgQwY5Z9TEyL9Tk8WbSfz1flaTQGVXEDKOinFXSa+x180Jw78ZbTVRsDRljL
RLIxogApOTdsqSr9EvMACsWzyaBTTDoTbtIx6F8t2gra7awFN10Bp8dWdxaf0oHOzw+ptCGsmiVA
piQrJL6SD+faMjJOozzzi8guUvzQ7YKubMKFgCMZQoKOtKVecoZDjoYghphvo6WbJneUYxjB2p1r
yUJRMFs3meI+1ZtmKua5BDrt+iWybjEPCuypgG1EtP+07M/aWvwrxegPMms3/hIkkhCI8MPZkD9C
aaaVxP8rkhdteeU9lk78deLUmdiLsONecbrkXE8zI9GIyevo1T8QTElf0CtyRjWY8mwEK67BRwzX
gu/h6Liq/ckb1OLeVt+q3P4uGJ5iQ/bxqtHhlsUCpZAG6PrpIvoLjJLAM2xDUpDEQwkt8/E4g2QS
+E9HP9bGVwfL7pbH8MyFrA5o2Ac9Qwn8e3QBV7pL1ayhVTkB6xcAQhLeR6UFlVDKI4aJZt/GU5Ge
IQHfNf3XZKmfQIJZYz9tuGKWW3I7u1dBukB9n9RBX8VH/fYclIvG+JKb2P9Z/Fh02p9LfFajKfci
R7tnBehpAF7To+2gVqm/f3Jb8QKjV3Xg8GkDyGSYJ8onnP3FJpAmYo2lVZ79oMbIxQWl1+xDHMpQ
bj5YAM7KWEdCodExaDhlZ3blZrBccJq89oIIRxPFIYPLNvrTWSCbcaxHh7ZEP0eB8o0jz8uxb4xP
llg4shpPrfjL5vlfJEEdY3UgBG0wzYYt+iY8ZtrgUBGnp7HLZ2oJuGZf0EiArQsZkeItYjj23NF6
BCORoZs2dVwZqrne345ODGX78ZBH6I0avFIpBgLYEt4+gEqcPvPZ0Zk94boTsc9T0lp8V6uXriFD
l+TcXTJqJzla7YiHNmKUy4DydVoROmre1kCiElsTqGgQO7O3iBFb8/Vjk13QfaEgBw7DeflXbVMI
OYA1+pvha8jxZs8Vdcf5dCIK0aD+FFu/UFjOyimf35QVZk9cJXwuKGVu7f5x2eUztcTB3gRTT2Xr
uE1Ik+fJRa2Y2JgJIEGFhq6sLKkc/1sGQDWS3jDpiB54dYo3kN0FKk4a8JuH9J1f254sPEjMY+b9
m/lHElnePiqbqhtTcpucES1i0GvHqIGYMloNpRgtc5e/EPgi9OU70BUgQ7rlAtYfu4k99HB4XmY7
veIMpPfa+KirGlc5FGLzD/LtoRUhn0Kszzn9xbd4OmemgjkgDfNZ4ZxJNWef1I86rIkabRliZnGs
szU4szXAok+i2UMPNNS2w474CcYrHrqqeXDotMeY/9UiycyAeRWOI5Lmiuocv6P1It6ntbVmRBdk
OjFeFHZUERkKZVSxFB/+ojiLrcPhSKSQvxE1EMvyQ1j+i/ahX8RuE/OZH2US0zW68Vc0BxzxmOOZ
p1hervKRf0t8Z8oIDZSNPFkTM0FMouxivH0lx5uSN18Q+SoGQgcYHm3LYNjDmbRWwLtid6RJaqhO
yCPsNxpXNLqyt2LJbYxYKCf5KND4GhasBnhhuGmAC3MDQQuMN+vchRm59LBQr5gwhFJk/NXfemq+
WvmTWw76yQfvgQWkvdsFBSr0CmpNsx+ouSZlvBuPuiL1cyL+TbkCa4wfd653bGKium/SqUMvWiU9
/Lp6iko00KexO4rmXc4rKHhS6Z+VgnLOwBDeWUNFci+HrLBG7JaUK7avDkiIyxHbM5xKqlYRQvq1
Hs73P7w0zPC6BmKDOhLiq8tU9IP55cFoJg2voiWSIIb/SB+zymAOaNnEEcKNJXc69XgFP7NmAiju
Zh5zAiF0N5GlbL6vVhEkKDMAlBQjIUHP6GczOxfTDpM1kLttX/hiPJg403fvhow5sS1PGq0e35U6
+r9EOXdY+5rBXeN8lWsIhizpBAzoEafJKDrK9AgFrycKY6aWjHbEQV6kEBpXo7JK50VE115/MTzA
eSyCQBjQgjHlM+qiOSR5XC1ITBhGKFU6j+/mP24GCwsXTZDZ3vNVbMOrDxhSzmhgvq+UZQ7gvdiD
Gjb6T2jfRpdh7/yTuJNTy1TWobD5jCpbVRHhREiZGjbUcWSy5K3gZulRKMtZzIMPFDmF/YOlcfcD
+HVr9OtCSraJyoeltIWZVgq0tc/wDH65T9IrooXRXXhINqhpH4i/3dVOmbi7a5g/DtBgeaY9NHzO
EKFqaE0EcpEQnEj/KZeSlrXV+NR1acTwPvJv85vIBi8FyA4gU6Pru5BwQnTHqSpGnErj2DVlbe69
O20bDSbC2GTrc82/aKve1VEOn56SJ0pZK9M+QI4UdhWT88Wd7VGQyNBxJmzGo/b5PANOy5W7ipyx
HIZDkjctx6fjZAB7APwH2wtnFcPx50ei88y0/BsKTTBBenJZsdV0nqk0kaPI0RSHKKctOLLZYBPw
uXH6DmgUjGlA4gSwC1ktVPyqAOTgc77Sn8jtUTUvATFJh1N8YE+dhKgGKPI4hgUepMa2YVrYdVtx
gXWtYD3HBGVQNOY12IZNsu52mYkzTFPyslvKe8imLXCkU+9cfjo1kgwUUl1zY/aaabyMZYSLpaFH
YSLra7kyx9AyBQvFQHgdEhAo9Ku730Y6D2yiVQZsBB/5Pqsiq12y/ygNTDEU92xqrvJS2Q/L9ZEd
NenbB1I+v+8m/Y6k1Ze7HJdr3srzZECA+mRMjZObw706znwq7DYib05I29nv1Athz86CXyxjBhVT
BNxBwnewgXiYD5Gl4tpSuxg7xuD0lxs2cIAqjnOtteHiItGtfbipRoer9m06WqqT2EZPwo8pGk5G
5QNxNFhZJd7BoohyQDvKW36dnOCWftKhaa3foldEWlHbKhvmfZHcWmRpeTxWkvlWffBHKCLL7PH4
C8CenlNGuGop6Ymah0yWn3RjYwnxlpBOGPDWvG3KhtUgf1CepcvrEX+HIXU5ozTezAxuQYAQzDsf
L+kPQPzTB/cK8VV/LVcPuNe36dyDoMnbIb+N3IdndVqRrMVr+fmfQOriRw2TERybY+utXdYMAYqS
qiPw2ZKL4WUjt4iZ2KyqGTGMvDapXGH4hP99p/tMH4MUxcDDC1zTUFreBjAdxNELcRlpqpR+m2Ub
ZqivLG9HJ/TsWJ0CMKTQ8gK5szCg2ZkF2x84ihbuIKiPh6x6nAr5PKZ2PoNrO4bYwY+1lUOntsPY
V9jpUTMabvxilk1jUIkPW5lnh7zoPjZMQxfGCp5pqlmPVB+P3+KR5RtKQ78k+q1g2sxG85j8qYY4
0uYZ3FW1sHZ2P0k/GoMqsvA1olPC8sfNWBkEplEQnFpMCE2E/dCsMw5qoSX5wi81d7u2UwASKG6S
LRSqhPG+Xrz5+xl5n4s/Z0aJQRnu4oLNRFgMyA7wTb3EZPCljm+JTJbdMwj/a7JW7F/kB6wXV4cN
QfKF/d994ihtVH2i/XQpIiwv2tWH4rGKqjwQfWV3mS6YyQOIZs38hXYVxahn3uymLot9zpFAhrKF
HOODiVxrxFes0YcSXHCiwGYnMCVsKf5Xs2k4prqoAG8AvQmoQtQI2TcA8UOzUTkocGVYpRvQWaU3
nJX33evKCsGJ5G4KzLgyjdy1weu49KnV8k7XZCVKyea2TK1FKPeEx1Fg5t4As1i1sUOisBFTmGfw
Mnwq/fjxrUw16ns1dWpsD36xMF92zRG5K4kYwjRlqYi2OVgGjLjiNya99wV+8okwxrsAd7bxB6Zw
iWnbA2xcBgBuuDfnHJUSJiFBp2WsK4dqiSVlQJeAMxCP8MPv+XnBGWI1eQSLC0KJjjgaNqHIRIOd
BELO723xJviSgHroHHZU0NRkV7EsAMRFzakpq+iuX97bVSub3kdJTl/ciXCYIM6YcnalzvnF5cyL
yhmS/2aXK1N+AjonmndrP1AadM38aEh76ZfNM84f80Xi+87HuebieALCN16AlbMhxInUwWmUk9wZ
jlqSZ8dYwV6uAakJe3hFB/mkCGn++3REuJMHKzX0W7SlfJFDbDoACpoeiMJPe/+ItAtCHgi7e3os
nU13ZU/X5UjpMRKmEZC1gTy64nc4IsToL+4fDiRjdDX3CmsbRPoipMdcZndfQyazi5y8ius3Qm1J
S8n7oAoYQySRgIUudcGuMp0MndgYpYrWWOV+bhz+HCxBrVqcMhG9tsfWl0uqPTuUaSGTc+MeJga8
g8bUrk1EZCUIWxB3d0nsOrRV7xFrE4ISQqp0wvhDgGozntF1lZ/KaoIIsnmytQSoR9+508I/VZh/
/UTqoiQ6udc/nDr8bIhj4gIlY2be2gYSTupfxBrEgG65sfj9xM6XQpA+ChO6c9BRstSVlkEeOjYt
7RgbIw1+G2v0xy2NMfcCk68NjSyMvtka/chIjF0c7cPf9r991x7H3Txavh5c99W1uE5pkIxzIKjK
yjgRcM+hVq7Ahlmm2xUqPydHfjdYesDAa38EUvfeOCwyMedrhefnI6KLqKqlTtFjJZSVTBkdCELN
Y3cCROvaQlkRdNEzDM939LRDxL5TSK9NDvpng3B1+JPNgnIy9XO/XsgAryizsOPzaIu30VHs3P3U
CieKa+D6rGe5EXM4HhHhgnjK/91zHKiGMN3Cql1iT+ppZlUjVcpWF2ww9UzAgzsxgQnI9lUjBLsf
xh4v6nmCv5sGelFtgjjuxVEQEFyW5m0wDdu0PxP7CuYrdqHOhF+RZH8ddwblmpGNBWOAlNGi5uiF
KFcrWDzqBpD5WO0feKvTpDOM9w4vBmFLaB7zl2Bj+6kPvOkf7Vl9wiQbuH4cDrlLIloi3GJ+Ac7f
VTaTEAI48rJGtXbrvAmv2xC/KK5l9b6lYjF3oX3p/M8a4zDFHGDsKr1OHX8CPznaumXFvY17THOT
NDycMD5Ay2w8t1ujYd2sIMVi+QRLg2yTljfC0JoMqJS+Vqt+FhjC5A4wNB8VkxC9Ucj/T60Ekwbg
oT4Uqin+B1MH/ZUqPH9DO3ISl/CZhxB1sZritgqQCelVrPcZ/ZZ7t8byqru0yYyc1CyJqqAo1cB2
0GebXwlAYcffHxEYv3BPkg9MyFFPeUIwYSRStH1L5NKniwr9aK54YuoKbBzcOb/x7XeaDsNZL6TO
uukCjoUT4bZOLb3BixINjxkQ8fZKcIAQdf7Ly4ffC5LaGNFA3/To2O8YMEZvB1H4lXvatdMz//aJ
3s/pSUDCr1tGvK9wCG1lXK0wzTNTLXfgMqA7utm19OAGwkSig6Q2w7yjXddPE6tw4ajK63fTQFbX
fSIX6ECHVJoPGxpq2F/rDP7WqNVermS7ueYCu3otb5LBPEQi9BLmN1hHPhDqoJ4QkPFPEH/V4SB2
hq17vk27D2gevf6XBqHmDaqr5RlKlbo8Z1DbIVgH4YFkzL1X3sGPIjI4PrpdJ+1Bv6/QXd9hUTkD
Bv7nstERBmxLJuwzsyQDM6EZBeio8UTQUQQJYGSWvMx/yENkoeENwNXyA5W+9a1NQQi64TiUmZZ6
dpQnIRWwDJXUDX1Ariy8u5WA0IEeGHOWI7ofaR3uCmrXjCetnIUFbCfFAOzEmsno+Df29MqK9q2+
NF5QTiTWKFDRTaGjSAcR5KhI5l0ghmkBrO0/WUv22tVWEzZMGeWAeVJ6dxq3ZiAZ8ullg6pEGZgl
8aJaUP2/vg39L7oGZW1lO9jjHAUljYby/MmBmgQVS8dM3bkSAWpteCtF92OQ4rCGu96cTI5QC7m+
iPJ1PgTxOGwnVpv8ek/UXsJdW+JJiuy+LBgPITrQQB8w7YFdhsOZRon2pMnrOOM5zeaQWu05O2Nq
H0YVbmLZeZH2Gg4gzczc0tOYAKCz6q2iouEHPA9HrqV8DDYCCeR22EQhYPWHrDGwpvhGd22+Me9R
2E8psqIfvx+el7zCuYVfPJDGWxMS9UggcUuwmlQiHjEjIgrHhjnolftY1ibLtpdABlXK+7YQOziU
U3/pjLmEIUFS7w+ZiC3fp2ofdnYB/uUku/5BRNZte8fjozM+YIEF725dwlG7P1Hxdcv9c1VAhV6f
rU7U0u4x8mhRN0+lRuzLR0dHHfh0SSRHaR7QhaSltzB4X5CI26PDMKf5ubs0ImB7S6JsZ7qGezU1
0NJQYflGfpvWFhZ8JyfJGZO1CIYwGoLzkpmXjFcwmeZpKViPuN7eKXGlTVZZwePKms8w//nx/3Uy
58aEu6N0egmFmZg0XsmpObWkyMUki/HO8WkKYNhbsHbZQuYyArTqVehXlMpteyCvSgQRTlLcMe5P
smUXZaMKC8PVIUGAiOBJvfNjcX/dPLgrEZ4AEOq+t3ODalejlnJevAnirdQVfVw/ZqYX8NmcjlJu
Vdkhlj2H7+wQNP1Sua+n2UwLYRBdyENYWgB7NImCAOJ3vMB5N9Nev3108dBOGxBb1j39PRkWfvag
1z2CvzpRFz1wibmpPHzCgVgV2AZ+N7/QCRI2+JyqBAFvbYqTVY9x+RJpPAehjdMlvvlPQzP75ZWe
PWDUNhk8YrQ+SlCou/yo2jM0A04fERxd5VwwOqM7Pghs9n+w0klz4X933oXFBfRQ8vPtXB2/YHNk
muhQ03ZVpEfft36f3dqhfNBeYMgnpWrPQ9UBpka6x2HWr6P7lXUHtn8WL0myWzB15XbPfHC/jJB4
yXipfXX1982xooZ0KfVCXpN7V5oBRGcC/4V/Qi02F8IqxnVWLTTsmIUrZgB8QrgU3RJ4fXPZaBCS
lGK88LE+2euLg5iTldIkCTtnf2xNL9ATWOo4/qS57F1CQINW1FbboIQBjuhQWy8CF3sOlZDJNU5F
3yLW2ygAG1ZJAJcS5ZsTjCjwcvE7AEfStVtGbzyoyQyW98rCQlpf/46xU8LvKbfo2s4D40kn318d
UaULzNTR741/dHBx1Kc9yynQnTQzEHvUrYop/MrZLJ7lz2cGb44zdGMNs1RMr9eEe7KgHORTtc5t
Y4DZ8fSQDsUTlPbR7eQs6L/u3UuUgFIMs/1vgA2E+/jhtwvHBwTl8Rji9Lqn15oVDpwFpZsx6I0n
/3h45k2NjizYysbUZ9GDIKg1WAkVCy7PPJovsnb70QUnzORvdbkERdAPTi0aB6BckSmfN0NWM9BW
OBvfkxL+5mhEdX5MemLHTVnNu0/Pfr8U1Jz37i6ySknmRrWuC7m4oSiP1J1NAJUbXa4A04mfW2Ap
TwFT26yTUxH+2hPrDRaITVoqRelGrzl5ltb+V0o9YQOuK3bwEIGmYZ/zGJMa/9Y1zhJtzrPmdDpN
p3RSjQS5jgeL4H266j2j0dNZgD2YGUa0ZNytX6XPW7hkXKpkIfr1ZosRqIo5wELZ600QY5Q0dZkQ
2+xs5l9NHBXX71jRP7Aq/mxv2L7HQkPLc7lXaWZVFLwCpMDX8Vs2TFZuIhrIP0hp/YCEvEfdfjhs
zvAGqb3V+5XkebSoDOYz4p7Ghr59xfSlaJBW2O3uFOnxeNlrn4O2oB72K0WhMoo9G4YiRWugOFnp
BbkT0YE69DrMaPhE2Cf3bMxyD9ouM8eZWwpLG1d+ZRISSqlc59pLBllpjWR2xx/m19mpJsoF4N+5
iWdBhbkz6D8Xzn/5Ip1rlit2cHAP/iIp5WvbFNOWEnb3O5IQrl1nE9dWXyHL6MMr0ukE0JBw5sGv
3rZFgEbPrk8ovSp93qiueSWBBrpUHA2NnKudbDFDGHH9Mu7BwZkANv6uEbFZ1LyFsyqrs4IHVMwj
2pSvBU9WIdrj5FpN4OOurh/7xJ/EurcRAbu9UEZPL/UCovBnYJQCKRUy755IzjZCNTezmO3+P+4a
DQQZRS9376vtPFhR973nW311G1QJL7B6n9sQI07OyoomucHFh2eXKXn0QUt+KtT3ArAcjsYptWMr
pFnPZ9Tk6F290aYft5lO0x89aYjZphdMG7J64V/rVPsrMTJqHc3qRNs9Fg4XaucYnHv9rlKZjn5y
uIjPZjGOKinixgPhRNfjpT4/6L/yiDG5KZbnA7v8uqn5DXOA+V7kOOFOU+lLXwFcnEe7tDI4k3A4
8aVdJZbVzm7kGPqb1ExKOg6ABGFfAMSPfxZlUqq9LAes2Qf8t0NgfnVIoy1RUomeAXldio12a+38
f+JyCsCy46hoyACRtxL/bGNAhELN6sTvnbfBy8ZFQxvjjhyXps0lUenTr2JrxqInxgr64bsdcShw
qc/aeAlWUdD2D+4/HUOy4qAy8l/iNmgaAx3AIm/514EXJ6wkNUmpCu+Xt7lQf499l4en/rVp3p0N
/U+7zmlgWl7tRw8w8lQkA0EWf38+tCp4o24AU0foPHecF6dHpSxG97+PZbplagfzblV1iwVqCPah
8gLkIV+DSpCGYQytSwwuMOUyCGzoM+2vQ6RfneibRtj0cVMLBQE6umZ6xR5CasPhtv9HKQBI3yBh
uOoyQXQIS7AJtpmZ5WpnR6GUvzUc3qf2JjkThybO/qNC04SsegXRNqtwKF6ZIvAdJdjcGQr0Hugi
jiH6ohObEzleHMLslUIzKxX/hYFhgo1110T9RmlSGOHPqPEz1e4ZXRft24nVI9hcKbBsplttyFzj
YyQfyum7m/UET9cjvAnhyfb14HqW0SSEEBM2IIqxNmUgXspuuhS603vdIW5FcyO7GPT2hMNRbfQk
pT5pAEpGUh5B0bCan1yFfVaZVVv22n7UAjqxKY/gOlzMNxkaD9P0HnQ9nZ/4+XHaHOLlGnERav9G
W20oYxqOdSvANEM9RM4xelRXpqazb3BRuYS14qMOOteYcuphPIeUkVvCMU+16LjzeNzhV4bDu/FK
UQ8HmJVyHX2o/bycFWsIduLLbyK8a6ugy7F0m+6ktp+IICIwsuPKAT9+Y09DBx0+pyzR5VvmM68W
201o70MZt7lYWWDuP2Onqkox5By1a8IPJ59gey81GJifukMyRLT0BMvbIiDenMO2i3HgZBrl/Obb
+tirqvaRzbEi+F9VwJ3L0SAJlsuyUSWAgZHEAFGiLFFXonq2UVyb0vm6r3FxO/heCNwXBwIvajmZ
94M9GSK4ygpFUgnhAUZGLl5mnHl2KGAZhJkHngnc7vOl/gWVGo/v8oLdGALx4WNAt4j5CpyL1qWx
6DsH6TF+HqKfvGnekMZ/ZnFs0GpAqeQo/fo5XeNMsuGVROYdFyPUTjx1BN6qcR/TxLfqyNvMBkc+
vqif77X/UffeQSYGVBjSSbcr4E/257LFl85RwHYLoLwahsjHcj2xX8qxv43ysRYi6E7iC/eN3g0T
mTFgm1Le/iYGVcDqm1D9ygXqnKOh6uprNaRFHA94FFKBHFNppo87tJXuN2Q6YakRXQ334tZPevM0
iNBkT91SAKuhoX91oO7qIsFzD50AU3mMyJekvfC0AJa55Pw+Nw6CL9h5Pldx/TnYoJ38mY0ksFxc
fPCf7xyW0AMAGp1/cLiV2RF5b2YGBgh4a1gvZOiVFYgipkfAB8iZU6HIe7IlgVZbKO2Ucj+kZKGk
dGCCkth+1/x0xEwT/mEA0x/qzKmBMZ1M4/Zcu93FidBcdcsGlxFr/r0ZKjE1UKlos9zt1lt/n0jq
MRtdzN3GPgtawOBirSK83fErJj9qcjTc7vctrDHuoweIMEIKAgeUHUnyOv2H0d4M/99EJs2ybtWX
gIb7jA7gJrD5ELe6D1bENiIPrLNWGnYWkz+O+Sc/IkONLthFPY5kptjFBJju3T9suGf1D4HSvTcG
4yVzcTmLfCOvEVp9+L2AjgkLIC1h7ffQpA7zEJ85ryrlUdQ76E0RuE8hwNG95M/UH+9Im+A9tami
NMyzKHTT15Jc5Mcc2Etz8aoDP8Spvi/LatYoHvrL6x0kMftntWfb5etkJ74b5anvsI3zXNAcFtDY
0o0Dk3MQDOqJkLXTatvnn8p8V20oxBqLXwuQd9p0c0YgepeQdZ5jKMXqqMum2epGFQRRMl9EHlVR
8Crzzt4bewO4AQj+5HYSFSZHygEXSUwxy0mT4yg0zNRvVlfom10WbSs2Py3VbVaBy/TC9aYjtpti
oJwKjB6GT+tOjFEYYaN5H4iAjK0gZZuwIeRaHQqlkZYiasrL/ys17oO9pmCS+bFDyj64f0/QD/4q
rDbG+6TOS52vvyppfh6P6p1SA6kbKZPCvV92u7pXPPCMh2B9Ul6TvehgFcZrPUAVoONmh/2bFhlq
3z4gjrNbMtauLTsysLeGAjzdmCIW2DSsuSrQO+wyiUXqbuOT/PSzPcWvwm85XSu6MLHU6PkDR6AO
IDeMVqyHx5mffhJWFKPMMaeXCvd5fFjoO4Ek7K4eZwH+VVujtYbSkYfjuWxAri2O1KyWdmetxQ93
WkjLB1wVpUbn/6PWuEhIV0IW5CRT4nri51XOUFm040zwTnNdqyMF/5zrrsc8eiT7Yvgj0WTqGbFv
KYrvNrp0GfFhmen4XCit3TPWetNegfI6blxaoMiXBv9vWjashViSGkZRwTXDg1d2FBn4E3JHA3tF
D6a1Jp4oXilLiDTQhwAZGiwOaYIOTQpITrsjc1lGlX+/7tH+3E4oD99Aximv8UP12TTiiyrI3rb6
6FK347uKA/kXvA5E/G5Jaq/bCRNkZVNE2Eeb9REZNog1rs5D3SyI/bKH24upI820+Vx5DpPu4eKo
tNj/gf9NmxbLUyFWz3K9lcniVm1mxZ5ccDU9c1dwH+XtipAkrVFrAGStYOF0YqHaxNyJnD8pV9I5
pdAm/6YJf4/SyM8TMAqlMdj+v+Ye6JJ36EM/TscLddNEzHej25NBacT/RHegOWgsrGzy8DQHNEp0
9gFBK2C/UCKPQ/AjNAqjZaHmVp0oSDg2TO+TBxXgXy9Mk5DqEXhC1bV3RtHbpRWWPB0e3w83b20x
prAnGJvkrw6BtXtNKXrURuak2qcsu/7CBbNDH7MBFBKpQLgowe+5dhumKkqNgzqStuJPtMwP/fll
5JGlxRKnKonGDXvry2EOZ5azLegnIdC7edm+QECQEbuva5wWZ/vdEqe+6vj9r21awDyYUDIR8Sp4
0vfswYW0uZk7/6ADPGHTLKDVoV6uNbnMrasK6rWiOja9O73RTdTMi9GKie/3av+Gg44VUla/sBrH
I97OSJe7BRGnzMTQFzX79oOC3rS8PmKV7z23Zjn2qIgEpjOlAlfzcNul/5Wn+FNtfFNs4h4R+CrT
hwsQxVe+g7tBbZpcnfyJrpm/0tcrAHS2ZUYA3GwXEmoqvpNOQzMiZ3CVUkZWJLcJksN6jZdxZ67i
k2MrR68we10uNaHplXCLdRDZAYVhpVsNNTObwPahJQR1C/WiR7QUlc1NaeZtgkpdw7IUc21rO3Ba
CSn30/4kUkybU1qvtbTbHTxUdsP5igqp2tPsOTKKG5sal0kv147eMmxHzzHmDmjdnITg9q8HusS8
ifWpRZbtUwrxXquiF4/LbGA0f1tsZnYing76HNFLRW9Wu2fbNtWOXevywwtLNlaA2hI08QNa67c5
4hhLtXDdMpt+7ukE6vAs7xFVCCmnh7WtKyzuy5caSWLN3CoPNBYtVHDLEx2ZXuegW+bhkaPOdPBL
+ozXAWSUNmK4yRl8aOqRvfKbYixvft9J1U1UZ3/SbuCen/qztHre9KIValvv6hpWOJnWEKAmVE+L
DujpwgSqanxnU0m8FyGutW6tC6ZBzrclcoFdez3IcK5LHis1GTchGpQeOl+1JURu/f+9V88zqvdu
+yYqNNB/Zfd7nIF0jlnR2f2meR0yVMRsbTwj85ZQeey6tcTjRTgUTVPNjFiunMgOO06rP6BuUvkr
U2yBOEIGDUg81hz02D/XpUWWZQc7ujDrcQvNLq9F8O0DIQX1Q+lvIx3HKtaRECnR5oLtsgDFXCSu
062FHOG0TfUKwHQ4FJikgOzhR1HL7rnvRl0MklKCySSYY7YEUu6SgsJ45ut9ief81q6tc54+JbXZ
kbt1tTl1spSUEKnzAWhCeezQnFHDmhVH1l9XJkXqL6QYTVhDTN8iWQxNahiHhYhs0uQwF7k+2SOF
wAcD6bbnvnyz9wlrlA1tP93E5tovM5ydo3Zgg5+yrOzcILxPpXAPSSsFrtaKM+BbPvRk8NH0+jOd
a8KCC1lqnqMce4LuaBlu0liOmB7Nrw8WackV3hJLmrruDdDUAhWxns/Qu0g7rt5zB1IExN1Itft3
wz6jOfnA47BuId/+htHrEo9LYkPk8zEF4+rPhwB5frqmleGkwUi/6+ouX0O34k/IMXufFFTl6KJp
kSAUva53eoVhZNc4W7kGs11rRRE6taQoNRVeMj1u521V9GShZS2Hlne70HBSUn5mXCGIdAsyzdpJ
OP0Azg2te2p88WD/fdHGqXuGV/fvcA5xlGkwWBRJi3CLObe4bCEmZkPwshuIjlkuQoE8es2Er/sI
K6oeFaS1/o7Zzvk6QnctgSnGcHClwSMyqZEO2UZF0H5wMnwn4dY870hxJ4kegd497oviOSjG5/6o
hkatxppIEMgrDkvIdPJX16ARKvs093qcUmGERGfbBRBBZWN4RM9CW3GRffG/zuJM9lX1hE82o2Sc
dFxavX/L7YdE0gqKu/rCahzlFMShWHxPxFSv40tgKJP0wV2wU7rvwMdKohv5cd2SYls49YdUnkiB
Zsybo/r7M8QSMNaSuN9ZEj1uxtYAgBz0+njbsxS8cwrcctYiC0hTsehi1lvWA02j3kO6p5wRu49P
TK0f+YBZPBdZNNluBPjA8Z2aH+3a+vCs477oLlho3QwsToYr93jaZtB0jShw2w8JAi0bl/kL/6lF
YGUtUEsVjZGv/5BcB6gy5qFzsjcJOjhxeZkF4XqBGXn2EPHAxdmG/A5gemjQ6wQYGNhGbfJXv+fu
qG9WvLTqd5rpEjbGTRHIOJ+hbILW2OSncmu9MKi57Ww6Q0oxzHbnlJdfndAtmjB0bHHyRQupPux2
kv0Jz+GWrRMH/GkSfOOCPbl8RLBXxdBgBOt7+x0zxPJUqXviuun/KtyBa1Yhafx/B9j5zuKAsC2p
eYpJuvgxyjeQTfFohvoIOsSk2N0uvbLRhS+j2JgYTLvpcjibMPivuF3ckE/vPfLU4kxbFLviJkFZ
th2fwbFvbpkt3s5nbJ/m5bM5iVN3Z6x1GSSGDbrylbFVndsX3JaCLiFR2AC5zPpOky6qwmwDN91Y
q1x1sVfLXfb6XDnMDXH5sBzYRiAS0kIOYhPHOND/k8IyVbDwCq465/4OEzQziGLkn8JjqorirT74
+lvIthoh3MYuF2S/e5EO5ZgRc0F/Uq5imKMK3f/0jKTfQmSyGKYorMqyrO0XPM231x7yS5yDerUk
b03hmEHRVdryiZaM89cXhIyvflSG1wpQj6AFWmCBO5Lg1TiaffmohxbY1b6jQ25aCmBHQKgsu2m8
SKJ70lIAYxn5IYnHot4MA6YER1MsfO4nO6D+hGCbZuoWJS6Acz6nhjllFInUVWMzlsaMMiYCSSB9
XnrQ8pEDTRMDGLZ3YxMMNcdz0tJjyncm/1C1bzxh8Wgwqdv5+s23ArBJobA/nUfGBs2Zv2pLReGP
5XnydhEjZgxkldsxLrhTWjzBEcfcr4x7+L8Kbud5SqNygF+d+cnhW6pP9pVWihRhX99o5B32MJqz
GNVf4xJf6OAO2ydSw6ilBDduJbL2Nr6vfhX5Ch7mWfuUzt0/SZ6kmC9/hfjyA+k4Qz5Z8PgE0FSr
swYugLp+FYnt+FLG66fDP0+ki7aFuh2uB1PeCjyYjpF/ed+lPehj9ip/LxZO6CGvqDQx5wrpvDPK
iaZ9Nom1C+7jCZCWpytpbhLnQt1gDEikOHG2vc/TlZOZSjz5oHaH3yX+Q6khWdVxPDaq5c5dEe5k
jEzf5J/jYa1nb5by8x48n9M66HLY3q3NUqZxSPHua7im2ntMqbf96IaEfsTswZb/xTTafjyRvlPC
VzQ2LN7ZeUkyH8naYIgjbc+IF78/wA3aOZMTMtR+QZ6gc/NbZttC+L1RjgLer2AUm1sjonUwfk3g
mitpoK92RedR4SoTOXx/d5IfGLI1UW87HamDN6EmyL1w6njHabqzocFORK8jM40Zh8EKOFVH1cSy
C9Nc5rP38D/fUlKS4PvPX/nd0HSwSXORWg5OycWovnK4176/ka4yXbB6Y+wTs9XmmlbjgYHlF6yb
2HpPHYrVqPWfZi3NbU/S407VNzZe7vYrO7ShLxprqwSu/Mwds0IDHhzb5Z4vk/omCIxzg5Y0Gbyn
lljJEsp5PF4PnZuf3Zr5acV3Q3/zoWlXe7+qU/BCBWopaF+NLwXbXQxxkqiCVew36Tot00TMPSDc
tLN51hHbp5uPSWDvs/TXfAKFTOLRAqdtnQVO9CAPqxYQWux5JspPpRVxEh2T9/4sBLzXevx5DaUC
3n6aFdB6JQSepMJPPtuDW9ppKbGU2tf7wOCbDl8K7lHr5HX4UdzvaG8En0xNE+C8Jt3Dr4xZuGJE
G0whC4Zl8N22U6jVGttnuqPa3UZcCLALGlcRNVhsB7BBmp+ndUpij9fGCtMU/cQ4dFvpuniFsPPP
k4jkGfHN74xq2n1DDBD4au/6RcWDwUlR2qaOuJBkTgKokxenzmIoyT3qV5TkW0C0ykm8/DtO8rpT
Eo9rYbfnipxH0bfmSNFxOpjcmxLzFqYqOnacjY4FghJArtGXfb/l1sb7wT+sMmNFPgbC+d5jVf3p
e1cZooYYymunhM/tVzvQypq7xKoVp9vRWplLhQTahh1cqpqXXEKX5s5WMLVcK45I41FlC/p2tkm5
AorZ7PLxQlnkrkr+Lx+HMwhAUggAY3VYjoJuLThhie6olk8n0U/kXsTiQYn+LZN4FNjdv0EpXFER
Ne9Ti9AkntPOq5ACKR726EobJhx5JxbWc5O08LOfslPE1A8mYOKlojPEoiYfsIracomSwQPayG4D
Qa2LvEyyt4/p1+mjZ1aWOjoItNkJ9DCq9GaxTfclZRMyYJCTk2qn4fTbBbwq+K0OqJDqHTJV/rWR
z2QeqmTl2F6dkZvCs7YVExgBFmCJncUTGPHqp8wJh/Wx4JJa41SCMdJPc72vT/sfHYB1tqezV7Vt
FLkFPZSK2JZsriCjFiJsymam+5nOfFE646ocWNSVr7mDW7MQP/IwCCtUv9SKqw6RHbHdQIcPvEx6
QoP74nl/p52TTzTrF7lyao//mZv0o67IFq57OSBALftYSCrEUOZIylD46CU2Xd6BK/jiqB+m6dCz
AEh7RkFLrWvBVyrLrsqPsa0LaSL5qjhbtBdR/6CfeGeI75WjaI6ZlCUuGzrDkh7eI+i1tZ1e/NLA
kKrbcX31gigUK9V1ebFiU7zLyUpqUB0NI0hQiF2JHadEMmgEcND7A3Zqp9+oiPlPkiyYKJJYvo/Z
JwzzScZaOCMiOwMg/g6MWIRsh/vPETHh/GwMX0iOVaP8EhIvkBQhV+M2ZIkIbc2ejfz1GvhKElcR
gtMHvc5gluQ96yQhdpQexMOMFwpsTYdQ0peKQLWsLkp2xedcCvF0DCPIs0U8/P4nejw2zpSPacbx
AIBPTzOxHk2WmTDxQuOU7whrqNJ0iUrunma/XPrl9+3oo85UEebyb1kRu+Qw+dFIIcjcT9n9B6Bk
Kp0Mh7/pmoEOxc4QM9M5eksie1VMYwGi8lN2GQPPylj4fjMIY2J6HxJTTgImmc2DKuo/TUVsEwLg
hmh59XEJ3SPI0FtBODp358v13C8G2txeoRtquxu/I8F/UuMVRwW3iGFGDk5fDR9XwC3A+Kegs+rn
MuY6kOaEfw43Yuk447JKauSKAe+FGdL6ZU3dJEjAveuBCMOoF/aJbMJ76jNuqmLnqOExJOwedtCW
lMqtqwCDzqT1aQVHtLrShjVCMW385NOdGrUmXtSHQ86L23J18h+rbb4eIGtlqZY1gMuh8wZBhO5R
fVLcb5C19oRkrphpYwdA+sgjSyLqORXUxNR5Cgm9XMy2U4qL1jklc6iHBBEo4K1ut8X3w7/kiFkC
xSai+LCMFut2a79ldzo7Ekgyf5nRca++fz7xiiL20Bp1YsdPgLTBxrFmuARk2t0TtuR4cxdE10eu
ibtVRdWy+NfFt15IdtZKfd+IH5TZWBsWYHSIB21FKJQEcfDcR5kjCKTQEs4VpQaDJ5uj6DLC8HZo
8elG9EohZ+cpd7WGV5HFFKk4pSY8caxc5cpTVq/PZEzKhTS7+OWGlUyDEsofHJEy+LX2U4qoGXxE
hq1rQKJucOf6utt+u7DIt3JpVy0Mcry6NwyGGV1W82qOwYJhl0p1aZDnK2mjBfgIDechkV85PHoh
ipt+Tvvg8DPvfxHvec2UhcVBYM6owg+3qzAoX91bbiKot/OtHAdpficF/7ux1yFIzQz5QmGmq2yK
F9SpNmeytp7krancUChhaJ0/WQUZPp52KOD3CEYooiB80LhdD/SHVoIhTgbyrj8+xRnQrHevZlVD
VUPODY/3Xy8CTb9CEhH8j1WbgV/bij3kcMqS6+0HE6G+dHf113wcCcciFNS0qn1CT87BiFV9FMXI
lm9lqWLF6C0MiQZRlNakE5U7yVSpMIFKO2V+vOJ3I1tkp7I9tgxbXXfgP/S8OKQk3oZwLGl9bPGJ
P6QE5PEAI1WaYgFrjtPaeiZMZQ4FaPSaP/olT6NPpi3dkapova0CGRHjcvYZIM0vLmZplMOfBFl8
oxSPPceXPT5fDT56HoNdvCCCQrgYZNum7dbaWohe9IMrtMKC6b2pXujMbGHB7ex0nPdS9G8BzRLk
yYPf2NuVKk6Yx8CodjmWgrcS3IJ32mPR1RIpfX10teglZh90VSZUo5uDWvY7cy2K3x1FhnKCzKYW
H0Ub/xp9yRd1M4ZUwkQYa0xZ2Tzqnvr25x1cPK/a7IHCjyDgsK1Z6eGTJm8zM67h9bYVNJLGdHF+
L+CzVjTnAGjcgxT6TPqx//uwcCAv4qxa6TvvuhGFcGA9ApXXxIyDCaP+ZV8bdKJC7vAxur/EfFlG
3nwWJLXwJn/YjHPy+mMQ0EgK0CkzwH0u1r1oBXWjkaSpOvOao2z18KsXGj3S6htchQed938nEhWY
TJSDP496Ol5l76+5mPiSd0EKMmCvdu30YcJ2ey7nmCtYT2jpfrWLPySlkmHTyRj03bYolIoG6Uds
KFmhDhp663qjhig3qgmi6tE5h9wYnWvAaA6xGOWlVpAmkiBFZ/p1xCXOhcrTypV6xOCKXZPMhrMG
a7BOQ1kU6KCN4j1RTDws165OEZUScJ8/Di2pE0TcbKsqB04mO9PWs1cJEMAVIwBlqTSElXDc0G3O
O35yMIDUZ0kO1jS7DX3h2WlcVarsrmaxDKrKV//eECHKd1ZHuYubfvWZ0wgQ6ldbqpEA7msUMW13
FsBSjS6wcfDCS/Y0gZGoOxbpWTRUv5cJyZ/7u8mGqVpEM7R5GbbAUXuxBbQR1ODZoztk9LI8oSmw
cDw16HDZ9ekUgb7Ay7SU+ILJnMvSsjfmZdK8jN9A2MN+qlUvCBFJcuf6zeGP0qSqUKrh6DX6b65C
4jcVARbk8De458mnx3OKUZ2IpMy8nVVynOfeVKgYY7q6ERG9C+xc/nhgnlIcp17NqKH5FlVeoMxY
mA2WxwF/3zwG0DR3FLSyxt9L4k/cesH/9u9tLtvMDAXKVrIIGE3dJlEFLKdUwvoRPkZIwYZmY6Mi
OZschIs5gKsL+mLgOdwZETylzahoCsvWGHSpcuyXObeOv5BIiKPZSuG5FAkTY/p5tQ5/luzLzPwz
54jetMQb5uP4Mu30L4ozZ5qCdgh4X3SWUZSU8mZoBCD1fxYT8slvlT+ecRL3Fge0Whpjx9bquxLB
T0tb8UNcI35P/dgXelLsnWHEqLqnmpVxhstA2TobF3k2nDE4krJVL1TqMCU1i4psK3bBvc3MPWkK
+ic9HIgK+2MWlGXQmfaxkr1jH7hQwYo7LTtoLEFtZ3eL4sco/OMWYkVIwSrWBJyuXukyRuEZyeAe
8NHpyv9ss9ptES3MgRYlEnQcMQfAhzwm5WSWhZbFrnD2OsZesg9bCXgv8Hz90kxCw5Z3YPWjwGt3
89GBGcrJq00gGAKcGCz4MULMG0SSRwBMokZaOWMFwpuBprtr/Db1xBY3OjKY1Ry1QULpBiLH7TCf
RHHD2ra6bkhKtMhTEEZSo4iXzhy5C6anVX4a55uZTelZG33LjVz3ePm7i3ck9CuJILRmrYeNzhkL
hw3UROxFxoVRTJ0KI1dnWNlUh1Y1yTCZtvdYUwUABoGI2UvJktbOIElgu4gP8r2QJpYyqYjIRA2a
+IjsvgBCEVDbaFgHRcJ9bY/oK8KDhgmXlwiRUEamVJs1V/1pbuL4au0QoEBiDx7W9JtrM/6cuj3E
npJtRS8QKwe05kMIbPtQ4WzqlkU92ntFnyTvm1WGHnAynq++pWzxHpN3EUJe/A2KuYpEp97BSm8R
WjVMEMYx0Ibn0SzoiJYVyDXTdGGuogvXskZ0Pi/CvfhZAkOm4JxdiJvDQzlJTyOG39rbgoqRqSK8
KdT5vPBOgFweRPrbGcTdwmMNYCDechAAL5CUT+Eh3BeZ0F8OPB5I8fcbZq79ToMbt5GWgpTeFrOK
HP/rn/NrV1EEKkTbmPlYa7aanT+H4dZx5gdwkxzrj+vxDq96PFQjASfcZPd40CEgGisq/oJ2zKHr
Rsbuw1yKLRZ6fB2nF71przPPg5Y61qpBuAu+C2WDopJsXVWSzt1B76S0Ioet4JFjfJN1lnUuDq+I
7qRUvBtlI8rLBdfupybcFn+XPxGbrb/tf4gk0F00tlXjo9QJ5iqERBZ1q0G8bsrSf0Sso2uyIUv6
Fvcn5umW1x49/uAtUtfPBBBWkQD+05V/2V3eba+srUSA2mwxQWQGOS3+pZIIltQ2wX9wDamAwheM
olXraxYCvjzKmo3jZWgJkyw+4dBT/AOhytiqOKTdGuip1gPQFNcp8eAKCPzXSKFedkz/BniCI05o
0+xbnBTMzcx4/cb+OdSI/TGH32yoJSNwstu5RFfvFovD7vXpzpD++q5goOACj5ZZDCbKmPadegmO
sPs8ZVTfTsDuXaojCpRiDu5fex2UUtNQhab3uUMHm38VXv16F3j7DBhfRNGEvXvymdvt2uM9zOa/
JvyNglotki298YbevzTytGybR5EpYYoqMROh9/LV3z0fWhjHvoi7l3mdUppNgq2ZzINutxUXyGP0
ye0io4RxLEwbWZIpSZ6PvrDBP+KNc28pwKXooQVXSdLpspWNN2wkwFZTCjIZeafAsvj0olWrhfwL
/OQx6i/iq4ewQrE9XXeS+RYgzO4HN8gDZ58pheNnL0JoRLv+NeJ/RgQT4ShzJ25/29enlV2SVYE/
Gc5jNUpgSyLRSAxxGOFkicLqpHogRmKzNOqrfSzd46O094CbUo5TwAApJf3MoimGgB79LoJBjIo4
b/ZvnGHTA4BaGUDU3CvvD/8ZKSCSbh2AeGXIbnI0Hn+gGrGqHNTxWJljSqVqS0t7hMNFs/qRXq7T
eeptFO5Qf5Zkgp3BC2aznSNbTAUojpMUxg1JV1vjNMGrbD1LbfD2lNEgl7bwjVsASSypmd4gcO12
BTaHmOXYKX0UHGmQ4ZI5F6pu5Miq5EjgFA5tRK6fmNetKko7vp6hEP8tk+vmiAQR+0VdvBAqogOd
XLidhn383lWl/K9VlxSFuXTS+rc1WCVcKteIFrQm96RrU/K09QuJcVuWfvc8/7JogHjrwtHz+ZZg
wW7oZkHBJYxHw9QODu+o2vv1244+K0OfT7Wbdcr8A/Entcr+HKvJjAtoOj0pMcNqNa9W5L/FOGnr
I0IaqTBAeg8GSq+C2UtC737fdh8M7Xl7KELYQP332ry6ra8yCU97snsGIGhlIHKOIuomrewNCRg/
u1l94OYnwmCwBa6QvQ83kRBIQ2h3oySM5CRGAaQnP9+8Y45OjiUkRhrEyUuSRhk/UziM6qUf42ZJ
kawLjgQqdWrgPImt3HNBwwzzVz2jDlPv8eJ8+IW9OtQW9JXQaEAuhkA8HthVDDcUqeJKT6wTco0V
iCz0BIk7dXUDlProjaobAU7tL3GCOM3Vx6bWvdEua6Ycev4yB0XktzGW76XD7724qEpCt+OBgf59
H8+ElPOsGWURHuZxfcE5Rr7RH60Xiej/xj6BOWudW+VZ3gl2+n1MEDOEuq6dusoKklQorZ0BYFnA
RtJWLpsV8ByxF7idwk7U3+GvZDnkDaWEin+EFXropkjrUoykLttm3jA0mTpeWQsYt+IemJw5SlKk
/UGek8qLiZfyu/p5tHZd9vuk029qg83NoAAQwOr3i8g+7NeOaA169tUrOdJqPHIlYwCrh8wkRuio
uHwY4NsqZIMwVoK07pTmSBxfElKIgdwn3wk2xmYR1rVLnSi4CwP8dJ1/w5DoWg1dY9UMtcsI51Cg
w0tTA9ci5IbIcrtPXqmmsvT4PMo7+/hV3GtEeIGi709mrnPe6v05eQ9TFYpEqZm3kz6CXc2WeKrO
QbPGjxSzP/hU6AwNl7dlxW/RNZ3QfayldEAwStvvM8v/f4qbFpZj8j5lq0Ox5Er4nO8yglWp2yPz
xPy/gxLyBBgiIsdkgSchAiNxZC8GG77FzQhM0dho/iBzyKy99tsBkmAie4dHnG/i94fELAK/C1Wm
uIyzs2fLPCKdtx1xy3BrNinjx8OVNXmkdLixz2/jg7EdgHm5g8/aAkAmQkNoT/C8c/wXZpd9cEoW
S/xWhLRSY3MfWFQcqcKBtgk4qZFNm6QnjyGJqESwaonZa48uW1m8UhdZ5olTKXPqOacLlpPbARCb
Y/K8/yhKsmEOvscKwL9VlIpx80fnxJ9bHOxC1xxdWJ8p5jg8fB5l/Kfcoo47S/ume+tJig4noDAG
Z/Z+cI4MdK1DmfC/MCyiJW9sbsUDaYL6zUhVAvbgJ7uP5LrbJiL9S23+/MVmBLPaqRBswQceuOsF
4FsVXcjognM1b3XnrOIiUDA5i9QATQSsZYU2piLYHZvnjbjV9YEeRyUzzBrPVN9/H73D9veYGI5B
LBfBixA+cMggOyrljr2e9xrjmEPX9aDHSF/DharhzkOlpFkcFniRpEza2jsJQC4lZcfw9biNeLF5
c1QMnB3OaPFimTjbAt3eXdm2WXsVxXYTL8AnizpBD2xg2bKXkBve3WfYdoU7xrW2tora0gwbCPgt
0DaG2lYNriVvHcn5+/AgKad060gYb64idIuEYvZTUcukFNl9sz29HX2UeuovqlmPZ4/KhNqMklMc
SkG440ilaeCCZahmGm73eiWXrqUGKo1v9k0JW4UM1wESge0WT9/cXFCtPhLwna10/pfh4K18tObT
rwBt77W7AS+r85l1Pj5VJKDaKY/eJkVO+NBroD32IT8EmSOuw/YUqiiR69ESInpMtqOwiVX3lIAl
5/vK0Sn0WzZbU/q7tXSMzKup52WM2PlXLuRKHLuguu05xMq+McubAjwlhI1ds+MTolkzzh4Zocdx
/m779ftKFEb8u3HaAlyLxht6bkxqv9UWuzbCAjnQ3d+/I80+nChl3qThOfeWfgjwHZumXGMm/g54
smyedALwsMdbMcV+3OcEvxR2zZkOW6In62FIeRTkwtHzqHvoNN/tLDrun64LoKTU7Gp8LwxIwpYJ
SpY05ihIvAzxCKZ6YCIrDhvEmIBRTy/16InVVWB6g/k6JPqqsK0AeVCgGIh2FX1FMHWERmAxO+HQ
eGx5/gSRSUxhlOG5Hxi6l4p1i28bAMYAg3nQ7vBaI8dizECGbsU/QbiDIluxIuYXAEPRx3DyxdTK
amXDm46MzAnp7YIZ27K4g2hBiVNpV0Vqc4TqUbUSbYZlntuz1T51MeUkf/u50gZhThmn+I5HJxb8
s9gCltZ+2wDU9WJnQ9s3B3PFxpVru19qjCBKhWW079o0YRIZpokGFkrm1JZUB2nOSAvoNby+L3Cy
VfxLHeLKqodV9eqCXu/UznwsNN3eQMceYoaCPodA+bqmkCWHeI67/yna3Rk9B/bXhKYf9vprgVW6
6+ZyxRSB81+BRMrq+PWIT4z3NyRvngH7ZaXiD0zCVN5u3f6gjRnWDe6bmvvEFaxafzbKtv/3b0Zb
ElYpykRBr0qNrMBzeb9DbT1tl8575Kbg0gEa57OBVTBt7lEZUGPk/zNcTtzDoYuwuHsmPuWt0NW2
P0iVb+ST1YeOmXkGoIkNfOeQU8pGng2vaoEbOmX0S1npiRDx9UPVumeqRd8bmfjvRNndlnz6oXH5
0G5b8cNd2L0ookhOiiPPVD+g4dpTJgLMn8VlEGM5/TvCL3LoAvNGwbtWoVLSuCHlT82+k5gvJxEx
u9+xpE5m5z8r5iMaIVT8rfs6ZiqbTuChqcJTkL0H2m9KvIICvXxRDc1pPhle+pGMnGKmFlNO79NH
fHLxYECQckAA/0wBaaDUt610Ex2F9qAf84kMvfxVp8Kz53YsBY1jea7ANDwfv2ReTrnFYGL9Odz2
MQu2Mej8DCM7eUq56jhene7kLAShyRk5iokaHKkc2/KkWkVBQe1ACXINUaaCVACZCp04fpXYOSHd
FVHMgb4bscRRPSri72Ao2qZ8LC4VU0Z6sTPfMrxUGlfhT0cMKkaP4OmCV7v5E5OvJlok3AI5eXmR
wBXY6pNYWgc/3NLetSfz5/G0ZTQ3172mcvAF8OAWaUgfYzmloTrrc26xRPumN7vk/T1tKwWXq52y
Tp0vfp66aEFU+PEOrPELzbfuDOYNARK0ZDBd7ix8PEBIVhsQR3SvPLFNQMsH9HiPSzL1GBzUAcMn
TKkTNYg61KIoLT2vFPdtJwm0HR9BfLdlax69Ht5yhfpeedKH8Mdj99AAjfo78dKhDprJEJpFJeGK
T/ruh5S7JjuiJKIwgAdsQzZi7A88YrXk/6QvCwlAC9g5WvYNyXpAYvi3XaJ4ZrddbHbQdFN5en2a
fugHa5UpfUrm4/jj+Qgs03CV6XPTh49850FzprXZjNZkxz9mEGMwWvhCrcQuYEMo7egVX5STkifF
fkjOpMsZ610SXvgREOq46uhjg0kl4coDc5l8uU39jGlw7E39x1sBhFT8/M4H/4zFLpsVe54AK15x
PT8PQmyZLg2dJ56xFb+6bd2HUW7jorajs8Gs3Vp7kta1tDay976O+cXPtU/4GrolPmbZdtcCJMXU
F4H+CPHCop2orPu0qKIsQDdIMtm7enN4Dx8Pho0vgLRxY1roWUHVm6f/Y0YiVq9KK9MVAcMfa8vq
fRlIYLvqpJXqVbUIAPCALpASmJKUD/imiGwmpL5t4mJW48zISfyLUcOkxgUmu7ok7dP3AvyKWfAi
3i+QHeuUHzorD4XO8w33gpZ4eCbb9bw4IIFFSa/hXNI+7/jKigwTR+33dj3h6lhiS1hAhakaZa8v
cd/EtqzlNF4n4BPzeqhPhx2jHVCF9HLNO9vSx8QcpZOS/SAiXeWoIQSAwTB1ZDd4EBfyO0qQjJRi
IdJEWcILNBDTYItPsfl6fpTtMv1qoaZIi0GpbRZlR2uQvUS31IiVKrup/Y61FxKBqZzgHnhu8Jj8
ircn/7kqPzE88DisGLX4zJlZ0zIe9KvFQMBVCQG240dfAe+7yt9HAHdZxLNXbbsztCoo5o4oWGTX
WL3Key5VbaDS23CopgdvgWMrcCW/RRZ0yAg6j5Z4TEEPvL7s8+9tD9AkgfhE4uAY6leCyL/Bh8V7
B+WInBKX8ss7lGNGn8yOeSwf/9VpDlzzVnEG7Wn+eJCVUG3RpsDhgnDwlSbeANQrm5F6/f2JPf1D
LnCXOlj2+cljp2xz3PiH1WKTJRoJWsn4DDRCkttEIfDIn+15yvg4sEYa+XXPnUqxcwGgVl1K0KbN
Is7MBfqqwKMhGnGOBNbBrnAfclYSZUXUSjOWNjg6/M91GgBxL/DnUQRoYtdCz+eHJhJQ9mLaZD53
rrPQNOwQVgwUx1+gvOL4/CtscrOxpbi4ALmcOEGqHdxi/qKtSl+CvXWeQuQF/OWE+ktgqQ/CC2v/
N34Q7HT3SLG7u2nr2QJRQGTG4NyxlsU3M8D7vJbvdyWoaXKI2wFXhGzCrW3T9zOE3jpHrikTRgwi
NGTftjBUT4vx0fkbrDotchtc2bpH2pMYtLg7dzbl3gY8VHW6n6xK+/dnYX4do2eJmEhJUi2CxQFe
eWOBR8/1GbLEOu+AHqvteOTo2xbLp22vVRdxdIPj+ueNcW5+rI55R162K6kLE8eKlhvMG8I2sS5y
QuUf9bRPg7S1c5N72Jk2sbLYW0EZ7JnxPfgr/Zpeoshhg7NvzkukTSqUlDG9wNckcuqJ171J0FCL
ATA69a1fd8YMeGNBcyi3RLrDTze3Z3SdmcrKfY2g4PK4fgiaPbQ5iq3dmq2GAl1mG43BpvdH1znK
xEmuisjMKXh78jqLxmtwgis0O12dlXiLDVBlafKPItzFQisJzPYtj6KkL7OPrEQJBGvjRzI4Bj4w
YLwc5zVLzSfgTvONdaus5IQViJ0ey4ANHawyY+EQih247jWS2DPJ+W2w/6moANxhz/2ipumPyEIa
avJ/J8ifGqxRrKxWfC9fYepBcUFqc0RBlI/yHNWRUj+LkbibEGs7wtCn4urPsuPIFTRaSa8ChGNc
/5JfM3HdjJzuO7CaJH+KTvNOtU1IoU2L0NlpNwPP4bmadOkEURHJyb7YRg4eIgBV3I0WEGWyIa8B
zAtdHCSmqhjIDE2NY7bfn34yUqMb79UEJGd5aIz+IyIi0kkbOlCpmvcGz4JD6pE2sGo8CWCbhJtN
7BSPsrIERLhCmSZElpTPSshzYpb8CJtrkDulc4vYqxtB3uTAhcsV5uZyCH5BHF4YTrrJxST373+i
EXF0MhiweYWcU3b35geA6vTmVgP9ILtUdE01lgqoey9M2X1+3k2t4GMFzQt3f8TqHOydj1hWL2MY
xXRQcdnGplKoGbUYebtJTBBhtQLQpwm+2OrN4brteev0utqzkOqLWuUZexTwfi42qcByA8PS1WMZ
RsOtC9VqNtKi3peWzZOA8P9H017CFkhdZ+eslOTG9DzURoau5d1xo+EY+8ec77MyAvm+IDRFdnw9
D4BE3BR2aO9Qt0GSEPJ1jxMTHS/5lx64cWVljhoSF0VTNWn0unM0UP93QolZnGmQ/x2J1XzEA5Xc
J7g3ppTyR5T88xim5T8PyDk+g17hM0kx40oek0S4B0EE2kOWk52qr0G9tWhBi7e4QNDre36ebPC7
WMx7P4vaHtV53lxroEPzXFAGLdgSthdXW7rUvY2qSatn8YfCPdp1dzWeFapLLIULwPLeIbtvlXu0
ngE1wPEvfqKnpdLlzlEDRvq9qSkUDIK07dgDOjDIYIxNOFseNMJgLLfexM2ebr2Knsbo1/hd16v0
XGn5ErihcNjTNE1cTPEYgvXtQAJGnhLXjG7Wdny2c5zgwoPSPut1uknQDK+bSj94AdAlwLtNyuzv
OWmp3eXhyBHRY/gstpsqfgKVraPk/6sobc8MsvcrqZYfzY7vv2IbC4zrGP1mINZRItD0wQ97l6jr
58ktBhORkKQdR8zhW3nMRPTUyvkA2nUQ1GsNizUa9LPpL+c2d8I2UftxUg+bm0Mdq2yauxkik8ld
hc3PUbok+D+9tkYCrAQ1yd5DprRfZjk104kHpLOflV9YP3KJD4myh+wCpqDXgjkESLBxp5m5Hxs/
oZBA48SQx0m7sk6OfZZO0FEeekR1Kiz/esVez3Z+Ora7yjHUTJACwfAb7RDWG0l/eO1dnTHXycYB
94twoQakz6Sv9RnfcZ4YONs1EciEGitdH/rq3yuaeiG6UAm7sWEGJpkvp9vwNwpe78q+YsjivGtx
cD9O9akSnhXfSJFXasEbHSgWS6dED2nsaFUGfVm8CgbApjoq2wCg5BZw28KIlIqqmgY+1vaqPL+x
3fqiUYeYiLkGQkgCYLISE8FA7sEMUxVBuAr9uSQUCQBI5pBbJjZlmEzITkKXSAzokesA+MqW/nYJ
6bxzQewi7es2x5ADsUiJTJhHjiEGEMXgRopzPv9haviksbl8HTcuxFN2GsaBzvJFHMSVaR+Ow28v
2gLJXR85FO9dIn6Tc1kKpZmV7nT7OsoqjYVSyyS3zr7mT1Eb4rcVeZxU1jIRPqwEETDWDZt1s/zW
S2hYhBGegIX2/KxzTCWoH1vVbEZ0V/lNnN9NjOhWaa2rYeyUNnYYi5dB6q1QkiYki/nM2C+TZB/o
9lCUL0WuQi0k2MnpwYY+cbGgg0zwAVadXZTlwkrNrR/oLtufUkhxqG0eL2OP3AKn7aZTvHmSY4SA
NgwVRRmiU29atVFmY4urdvZUgBniymcH9GuSSAI6dBxmUeMwobLKnZLiRsoblVFBALt0RQ9MBpME
+841jgLQIciU0GBP42yjviLPg9YzViYHag6ZwInzv4RpsiOo60EK1YTnBYnpKOZNKaiPVWmCdrT2
cuca9F4hVqkw91iLhIGQnAaRK4CaGDBgFeJ+NiilI5JApv2fy+PEStHQPKIT4mk7UGzdgEeI6Sra
VTeRnQfyNusVCl2HZ+9N9xbqWMVxZ7lhYJ1e/GwlRoiS835i4cUikgrApT7/Fmsdfdvpz5DkuUwX
hQzHosQxROXWWi1SgqIT5QezJmbN+rOUaxypNG76zEtRwkxGwJyM/XwEAyKTQ1xt0hQfjL54OLAv
D8tVu/TVfdbTXb1B+ta2rVeOSIY87jX+ZzaehoDIdMSy+YumvM6XawBJP0GDzCjX+QPBwONBqRDs
1bfwlB/uJazLgAFjAUZc83kEe7FkQgAWaqV9A4lxff6BiNjI7yEw07s3UeBzvlb8b2QWqR+6IIoi
FI+EYx8CvQTZgHyln3cptU3eHICY2kw45811kAl2opxpPCLQQDTbGUsvXfDSfc5F5EeN9YEZFWKe
cVPPmrv3r5lH5Px51PmFS+X+chkXxX1m+/A91iiexN0GH99EZTHgcdB0W8wLQfTNha727zxGfS/N
8HMCviI6vKgtdXbBzFn76U5LXLMrsBJ3/JYMfpnjgYpVVoiHyudsk4ZLLveUpMxc3KTXE05htU9S
+FppsB7q+qL35Y2f5PFcxS2IaskVnhuLZMVM5SoU/xSIKM5lrcUG9ER4I/7KVxTgDCjmqCys0nRo
CCV4lvQ6AADPTNQZF8jCk7v/S4wqUW8F/P5Jh2Z+SZITAVsDSQ2ObsbwHpmxfndDKcbAToGkAOHT
B1p03j8P+dmzvCtQqU796Vw3B3Lcj48+qV04xq142kKWL9ADB0zOP6yPUFPdrVBwqmE4z7urK4HI
6HU/dnZWRFW9toID+HvfBs3mysba2QeB2FJx71tKiwUddo0zN8AeJU2aYyAGyyC5WvTXzWfyBaE0
L/7XXNxKVq6oXjF2OdiQ9Z9tDsr9/eM+/j39dKXyH7FjbTI1Syk9UsLrQ9KcCkRvMHb8DBsMIgQn
WBkJ6F6/WZYBv12JWKwDmWYAu9OrZotWrfjvyJzTIf3vW23ZtmRBkQnNQ2YL6MMRd0qX+uTOceBp
WR/xYL+5IZ0whpJPFkoUYeTSiHNNGZ9RDyzqRZAFAyBjpnIb7MFRn3S+jDgbU62cowtpYCxMZokx
2jt8y3djML27x98fZPntEUPUkRK2UKm5ofr+/4rCZ22oJ1nWw6UcZj9rE+Q5txpcpCUdBwkAL3Hw
U5ujm+g1fH/B0SdlWtLWxVvD0VxZuOH3rqP84sv80dks35p4tUSC5Xap9WsnCE20WRRz0WN9dUT4
fEjzZAFrCqZxFAknp8WSmM3k7VxJZnlh1fNY5w8iDObPKUTQLiILiO+fh4X4AGxbyxur3Nm5VLtI
VzHikg8HQPLH0OfG+f4MpFp5pgn2UOZr6O/4TOrNQg6XtvoF3kaCYXbGjYcdZZ6tmePGAvVbAj8e
yZ3MlZ2xe9X+zqYhfdHwASGwrdfYLwKu+7F6fx6hAt+xdu7k5GpBFzhpeMQnqQuqA+rHMiaKB3LH
fjN71rNTqxvLRH12k3lGSKrAR5iiTDmDrt6+vCHZLfLkova+NmYviOO9mLjYDR35txziDOlJvbb7
6MgAnlPguryrrNhXtLlypAP4s5Yv6HTFx1ePPUq8Ji8Mn/kBFM2VJ/3THoIWxGKlh+I80QFv7bCH
M6/GIHfo61RWpqkTVlRMd1HvBR2L91HCLLociUUF5M2mi2pR0Hphrn7ZwzLDAqkgbwIlyd+8Puj2
rdEinINS8DaQyiGydaL507seZQC9nQM8zTE5znc/+TQfD2buiqNYITQVbgrIzAdwzAFeaivxTfjn
d1Ws+N/rWQkW2LSmj7BCYTsfH+qYtZEjYrAVbmnWvM01fihcPxLiX5h/R9ESVCP4Rg/3Dabz/+2W
txgTrIDAc2m0nIuWYTcUqLUVMzDdtm+NuvJccQ5i5JF51RsY9zk3XcAcGh317VBkgZfxIILnlI0r
k2RjMuJzWqnE2QUULm5vG8BWTv18K9eZPJsfN2YX/Sp4Pjobp8LwsTpieqzKCKW2XwIVF39fF7AB
ixOZ6iqwOQFkCH5XACWCSNYyM9s+E0Kc++8DqIGFX7zE83mmSlCn6Z0T9and5I4xDwmXOyGNM0+H
IR9HgDMgd2y/JU97G1v6IyhgKu/B6ylwFSzytfSwrDdkgG9WceG69bxHe7ccZbzscjpmdbtRdx8K
MOJ6V2p1VB7MhRIW9Oz819YW0Q4O5clbL6SvSPXtoYrcPi42Sz2A3lmv5HFmSSQ+pQ3+Spt70iX0
ZpyH6dFZ9MRlHpCD8iDiLbaue9YIF9aEVmTMsnbvPQnLfmgG+TqsbP9LQo9AmPidY3QZR37XvA18
4apNjgjNwNf4UVQQ4yVCUxX13YbsdbbOIfPC2MfQ8c80f8wkqWGwvQcqFkYldD3oMj3+IPLqmW+w
J9Wmd1EjwNHS2SaJR4vKBelG6J+KOGRUYSWUFr8/imp08BOKfvjMiOyVh23CJjOUE0R8J9GSIYKy
CPtQYIxPx+zmFpUBTZtNFWVqZ+Zuq8mFwvITFrQkFZy0mv+1NZuPLRkzgVUZbND6MIIoMpvwXs1X
fLos/q4tf+V/KV1TmnIpjJPFBSUwdAZrkjnO2QYfEPuCXIoCVTxIvZkwOepjN52jpR7zkSJrZUlG
P+PAhAbZ2VZGKKOovfdueRFZfg+h41SDyHhx/MlRDVl8da5+n08EJ9Xe7sFwGnNpkA09ZrhElWwZ
Mufa+Gg2RPXIxYFYw3bxDZ6Mb94YoTHVJf7BsVhFloMtryYCovuPsmsaUvnlkkjBRAmxMg+swB1P
0MiOTzqTCDzZIE4JQ38J9BLrnFu8khwIFaYU8mplis7Uw7D9oyRg1i/iKGFSLuZXWAfGb+ZBE8EV
hU2hzRTUKSQo9kMHmGQ/eREQq9p2USqz1iuGxozppJNcfgH7oMNV8IkD+VRZqG9M4bQkvT3RxCRR
eEwDb5xuS3SyZ6qpv4dwAcD+Cl885bD4OtDX9jh/FrX9usmomd+Eo1HJ9yANM1ALhB3v5gzaj1Wy
DtIzHjxZI8ibBslLubZ3/1dsrrVlsC0NZNcRFPqd4PHM9ansTNILlLaha3y/wddq4T1um3ihMYhr
9MfxJwYPT+v6AcKDsyEYaKgCdrVDO6sUfPtyZQdBeVbAD8GiPzDJ1ILERLd1bPumaKTpfaaAk4CF
WmOdbEbHy6TVPrqg+3GnpwcwCFP2GubYpWAjeJJCbVgUfkvZiNGsX2QlLY8B20Mh70TfhMnil6+6
rZ/1JD+Vv3jUm4VLMLbSqn2gZgLSh3HfrRB5422227t53P5Ls+ik8VKU0Rvvu2tVexttdKOqipye
r3ILribqr2FQ1yC1MVaPIoNzqaEMVCxfgmDH8Q93ITvHbiCpBggS+9kcV/GmaxEQ6UYASb8reb4/
7Wf39INDHyaZ+JO1Xh40HIzhKhVO246hOyB8c24s5IBp4/wjvSxQZWcTHbFoF0nZmoFiYCA227Ab
h5HbLZp6xrdBKHNkhnUbBugA0dKqJ5/KIXKM/+xgRIVss7srn3TiRrH4l8hfbbIdi/CyifndFQIW
zhiDmkNW8i629AzGOn1Avcekio3Ua9dz/36qI6w530su9fQVf4dC07YvqFXtm8GVPXb84ySUHf2l
G/H+kQ30FLfRNUo9ZkI4rM2T4hBZVlmyYNL++KY/ih7MoIeeBnuSfbBoQyQa5XrlMjPExJH0dLdb
iumsJ0MqwQXrKSSxdXGucEAhHQHkGjQeD4XH+Of+tv+gBjPtABMklrAG094U25Efeha8OITZq/x4
3+k4ZOQKOlFzHjhT74Z6yCrdD6YOIaYa2l9QBjHElN4l8sBX7UwVj3wNhu6zSCTNWh5tU22Pmr1D
89lAeWUAQIFe3QMwBQid52ztSuTnWXxpY/sY3+NXiL+cK/J2AiyO7mfLmIB6vhfUVwsBZTalhoxG
JOJCVmAdOlFfE77ldtpmFZlQLnYwls38rIQATFOxX9vgy+rbZkJX59TDMaQucg7IemoJUY8EPrMs
GpYGp8PVkx8lqvLHKhB0KNcP9uNUYnkNjC0ATTbT8/84/Ijgksq0xO7Ms8elRoFzZiNyp0I8804Y
MSztOGsx6ASDN8rueEBhTvVx38OnqCMfuq6aUIOnQMSGoBlvoVdsa9+ES4JSOv3IPK/6LupNN2wA
wEBNgCXd1+PyuhbvNCfwWAMznzguHcxqR/IZkppckZ91306GRTwx1+aOlvlgha0xiAQyrZgK5F+P
az5zakMh6N7TPQuxOUsRW8xTQj5AKFPt6ZkQALvD4tALndU6zBR0O6a/4CGGNh60EW6nZxa9IR7a
4CrwEM+TsbbRWkEUpcOYxjPTYjG/nzzzZNpPsU4E99OBAxKyPtDNyJrqFmp9/aL6lRg0mMzy2zXx
O7ipJS1SrPAv14LGAYagRBv4Psq8ft1Hy70HjzV5/bjhvHsL8E0PQUu7P+Iq16ubJTKZYXDflTsH
BzIkWcFY77JA8bef8UjWgMPd0NagbTcUUUP4Kw/lG0gZm7n8MmRtmg1zM7OkgQjeIH89W9R9A0j0
CUH/NRPLIgbsDWoR+N9/BGNBV4u/W0JKBXlerRbCp0bXidE11h4q8ue3LtNUVm4uIAiFiXJVQFQ1
dgurpDx2MHCX73EeFyX1WCIgjdsQBh7ySq+rpDx816Svj7FoL4sXL/8ySysSnCAEpE3O9MIbXf9L
ycXUr/e9EZ4z+qOZ/9qUZconcpRi+NG89jng1usWLqN6JjtxBCYnMrXy0Y1+S+kxnylbw6aFc4sy
0z5z2SDy/o624B23ZZmBsC4WEjwIxfYyQUZiw/Q9BoSjhPxZCTRKgbfq87E+OK+8nrFwOjdH97H/
snCM9oeUagvanKtOlspvKSr9yuOuWk7YSTFs5jLCDZarAiqgILlm+mw8mZ2WZ8wTdmfKnj2ayIF9
Z1OUBgWQZyLoECkuNbujR6D7cGhVcij7JZ37TadzR4jwRuKUHWWmWzmGHeX+dy1jqAIh6FvEgUmX
RyW1DEwh3k1PTukmjpsm8J7gHMpZzjoTnmEXLHfCBhXpNm6eBejGsJpbUF31HVIvE67MW3Y/l8yK
M/s09/oS6k+euIZ9kIWRXvRpo153pgaBpc5T1PtB0QRsE9kkYT0qQ1NM5kLTRGIfYAccQXqC0ab3
Dy6kDfjUNqPZZcI/265J7aVsPAFvgBkuL+A7i+sB3LMZhTloskVS/yAd7MjGAG7N5EcHrvJsQYCd
fb8HOOC8eqn+xkSvYJ4U+sTG2+pFlGwkO6EGAqx0alF1s0ubJVQFCDEYExoNP0BPgwPvmzEUaNqH
9rUCayipskpIMjUhQ5l0YWWjUZmukQS/d6Uh8CpqIrN31bzMMWAb2sD2YXnYuJ418xVTzpR6DWdz
H6MX9XDccqFs1QH5DdrdY1OuYO5Zp9t3Am3feKQmPqEnHWYMaH2Qy966JjyuFBDYurqzYLSf1oUA
WO5aKYQhY90IOphQ1EEdOHa4+zgOf8/UZfNZixrlUTtAgC+KHdPIlB5BQYeVkblDNrE/ZZnUsLq0
CstUgqwjUoMdo/+8uSgibvqlL+cfcsHHYl39mL7ZqxV42Hhu9BtTbVQcfiny54A9z8FjiDdEAz9E
FQLDnnXgB28FCMKrYeKo2rTccTA9KjmDPzI/xbW3PiWX1Cfj0GN7IC6T2lAIT3S4+J618YnCAXqj
uoWCvve2K3f6NaAYQ5CNZQN98GzF6KBspeK6qaEGHPtY5h5i0L+ODdSN84tnptc66UTX6mYk+OKC
v286btJyaRcBxgtzNAcpyyBU6vhEnyatu0073xa/cLEJ33bdHQfQG9p8nXdLVu9UaCAc5k7w9QHO
pg4UQkonvRcG3PYK/cvTnKIFeT44BXiLWJ3H1fxI2rB1WnoTYPQ0fjU/Rn2YCmBTj1MkydcaKnK1
DApTTIQvnH9Re2eCzixxyGhTinyZz9r2VkYfhVEkHR0qpKBpUE5LQx5LpKKgrkjYxFpjljx8Biao
yrrnjUE/SeVzJ8frPc9ei3P93BgHM65TtSQSpAbpm6+qWzaxXWwnQf6YnuhcH2Am5k+RIXVsnGvU
V2B8amNinzNlx0nnEANCXf5j7QjSb2U8ZsfhStFswv9Oz4nQMDe7yZ27Jdzq8gj2Q/LmNN+0yxbG
AdySUHdvqRHoej6YKJfuAcJN2iwjtQK/0DraAyzwVrY/hn2gjqinuceLGNOUMqvRCjrijhG8/65r
F7iIT5hgTso1mACV++cqEzh5h7mLUaTDvybeClBIY2K31pVapZr0NLiI2V41n+l1PQ5q+CS62Sdj
9BVV2wOybLokIHx7j0OQ9LwnZFqcA8MdJgP8Xs0VLXlTcLyj6oFVP/FsHRIh0BWEBxVsiskLJw63
K0+HhREmKDtLIS0gfzDDigpR7EUe51YTTXUfbULuYBq9KYe4cAQDaxZgSHTatVMXvVw/cMJlQglu
+Rj32rU17BEUA0Ll9yMm1SYHgqWNZ83A6ib0hM0jruFmi5eQp7erzf/15G0TE9cT7xGNy5lD2rTP
ykiTUcVSHLQXN6Gx4qmxc83MnduQqns6y4CJdGSiCr6UUKeqTi5NGV7YPh/8XnFRhYpwqslnGll3
mhCeDyj1U+qs9EleB4kI1+Hs5lby0xRfhX7h2u+HJmDMEGgnK+XlJ/zEm8tIVqhEbMZqGTeG7ZAs
0jofm+GxYjiAWwUQgTJ1rNMsiQKu9ve/UKKplsAqrT3HuRjzeFNUjRfvaSodhngUwmd2YBFgmQCe
soCmOuVVGc5f8OKrHYZ57deQWFXc1wG8MUB3YHK9Nw642Tr8mmlrpnz8mGQjKKVtfJRV4zP1JTbr
cZT2CNMyUTWG5VhT4157rcORRtdJykowXKCt/zrhCsysiIJumMTHWIAPrsl/kaLhmsaKe+jM5bm2
AdTwCdWRJJGZCspa0h+EExQ65U/p/2/mwxzbGyK39YGtrHb5bjImXFBbGn78WVMPJaO5J0HRsJ5I
zRpnoXS1oLFcXAEmQXkee8Z8Bdqv8HIUl/IHMAL0Lq8R4B9F8FDjKOaYIqOimL1ZFLdpqkI5y2sJ
6LeyvXNLdHO4D2iVGSYloTl/FOdTp9kSIBfqNx8VNtqRCJLwT4UVczK2ZsHBi0W+bLk48RnNdcQU
0DM6aRlvq1hNkUKah81HGK1VQe+oNyqKlAJ+/MDY1zOjkFVgMUUEZEIIsFzAc/CpmbRN4iqGunky
qEVj8Dv8lnpONu7hMNFs+D5Rtni9/RNEubLn95rz8MofLueBm6CBY7Dd1xMKCK45QKBtAEorz7Sz
GxoL+Qec1YBIgQFRApzAP6prwSNSY5H/6PUCVLkXrPX07vYosNFRB0Zvi21iVA38M/bx1fA2fqG5
siloAymFlGbSsOyGksNvubdlCO3fAYADXwDpFxWXbUVxY/Xa/JbyYwZBpUkqa1dI3MpeZZwVBVrM
KZxHp/Yl39OHUTJ4f4vzemIQvnxEBZkmo8W9h7L2FgnaIFOOpXTy2+l174G1x7qSNYsn2yV7em7O
vEJfZO8KZKG0pTRCfA9EnqHuyJz8dB6UyCfPtVf3EiH1303lCf7xzzsgw/gNPIM0qV8jLMh+pYNN
Lb/NRbEu+a8Dnxgahe/cAzjUWMAYcZVAPJsT6ZUb4b27gloCg+Z9VTgn5LSwmATHK+o6R7cd+9Pf
4fTBkyLOQ7NixdbdWB1cMEVEuPE+YRLQ6V1Tld+szh/zneqdtCHymnNH7ZsgnpFtMphupFtzPvmr
ZtKFakoM2OpcbKeNSGlU/BH6HWgIk7uLQrR2pq49ajlNZr95PKLRiR5hu2jaZvaSoz6NfJVSiAaH
70FE2huKBjL0uR36rTBIo5Km31Q01UOOkuMpvwLDwvOgO8WbyYgCesDRDqhUD37J9LePtyuhTr0l
zF8y+fAmVsqNSfttf4vPFnA0kl25Ly4wsDhUu7oxVuXqTl4P+ioCDnZzZ1vLrZ98XNp/HZrPHb0M
tj43eXxIKY4txgr6pNcrk6NUkNRox4GV84SidbpBl5u9ILyCAmw3nuejYcspwNIo3gqiAjKzZ+0H
LRjQhoJUEBUfIzSu07iV1HOUlblCaAdurSteTEx8PDBTSQQuP+7rLe/QobC5W5Vu9E9FhOe+Nxwr
HOghu/nXYimy4A/88A1QS97iXcnnt7+scgOGG5hZTCOt1AJFsHH8wUOuZbPHqH5aYrNmbDG/eCHI
DKSIqGl5WeVDku805AGWYu9XArsA5cHphjgDBuporFb45m52oXqjUiW5GUJVfEPkk1st8EtpdIye
CBOkaaN5BvSfVk2ndXTzllpc49+kg/ivDJWx9ynrH+76QBu8TQav3LecuMjGzptbTzpDrV2nXbA4
6fawwvgnXFvoVQO5cS5ya9uE0S4CoksyQtBi2VqBRQUk+DNwFcnPdeFdmYHd4PtV2SrT9A458RFa
04mnS/G7tYdlCGMooOtKpIFIedS9C8H9KHVbYdGkmqwyMyqv9lD/FcySB04a+4sqvuhnRjS8O7PP
/nhnx5f1xHb/WhuCobj9nOU4ej/dmQ7M243oa/kS8moer3f1nTqznn7Fd8G1/72mFWO/YZMeEY9n
8RWi/1kj7AnSfScmHuMnFfB+hGw/spr/h3gAHaTXjU89jVUrIQSLm0XsLNYulQB6URvR1qPke0LE
WOVXqECtH+m3YBCc21Mlnj6jBqMfxnaHOMc5a68YNC7nmozvmJDAyMZp+TAMw8APBVq3mKcY7VJu
3mbCMMU2f6ZKYSZnjajOGKypz+lK7BAldkh2fmb+jnm9Ey/Q8xKXq0QfrmhKQX9TdlWfesKpnyvT
a3KAMxDXPu6SdR4PUJHVjISvLnyoXqLF01aR1M30opwtooLXN0M4rkwSQ44xSed9cyBaFd+Ib4bW
t7GCncsaWnYvziKMiT2EmvkJJh9Qkkmlrlpz1tbYx1W16a8MqYP1EE6ia8BOAvdVGRxsm5TFBN38
AGElEd/Qkp9Y+TQaI7kC16e4EMnBCjB0A3xCu64ciB3yOfUhiKleg9vZN2KqiqGu/YOYS35kurSl
/ZLubSo2ZHhRR+GTHWKxxxeOjLJkaMtSV2lJs8NF63wYLStu68d62r4vtVzLNajh5WBmHIlRWAHH
Z3fdojPIosk4zF0IISyFjoK/FvKnN22SdpF9qRel+WpLFBc8paat8F80r3ZzcuIbUvfv+j/9H9C5
gsObFDCrjVikUFh3WzS4miaXbL89H9UdLGxzUbO7zUdkpKKTInagAyN/CWvKShIsOJzT61sVIRJw
aRj4/sWhA7EhaidEEt8CAk7vc9qZYxGojKZo7GOA4/LyZrIVEDbLJr2rWGwsr2FV2Qsu9ApOiNil
9/eKCsbJtckUDdysTqrDYWX27k3pFmcq0Vy/URYymuZeDPAE5EvuecQpZpLlnKlhtU3iWUlTR6Qi
cIEaWcu3tjVBIwLdnSP+mqK2yhn4LIyzPcgVHva2F0mXiOvEscHgYYVgAIee5VRM4xVq6ISPl6HU
5gMvSqn53oomStl/ISqjy4UtvL8vwIh2Y81woAqbvFPwg/RE9JKp/PPpqiTq1hPkTIfZKUjMM3tZ
JOL4+v/stlEtb2Y10dknPWAJuO4uER3ZObmMNECceFQqaMgZ3D0H3fmRlVZAtgW1+MmeQGb1Ha/G
8vQdrpo07BKP3z5ieU/dZKzxt0FtsruUirGJbBXG64GXwZLRwOT0hrR+rwhjZJ3dFUbde7b+sUDc
O/Q5ZQH/TvXWRuo4ysSmdzs9JySjj5g0WDA97kgvTQGuB60DlWUx9yNpKMBGMzxRRGIvvvCn+mb1
ps+yplmA4YzH0bsERUk2gM1QSs1UGYx5AQPfTJIm435MA8fNVTMMBbSVy7hOpFTeWVBRNd9vWuuj
jPiabU+E8J0r5759r/slpDsOrC9j/c6fgDAHPxLHDGicM/z7Uz/jH6wiy7tbX5TeJ/HhaMjjpLWR
2RyfG7YfUfmql/BXyV2P6sj9O2MHjs8zStO8yCq1sFN8CWtcmQWRPlDJowmTQdSN2xFyWDuMnYGY
jTtvvDEHmMgvb2hBPG5aASu4ts7+HiVgnYPzgtG9KcV89SfFnfMG7N/+YQ5IUcrMnSPsZ9jm11B4
JomPUZQfa6M6Fzhyad06erXTPKw82txlPZZ2rTf0bmbSbnSdGu2k4VxV8OSjsfRHhNGjwNX6jGlj
bD8Kovsch9hJVzRvlhn2AJbx2Cb3DmLk3rrzGtKtn56sxHsA45MMNGObbbQBb4R2nOUKcbpXwmh0
PkwHbZQIvYtfkMnFIcKApPsRBizpgZ5wkcYzERzBnJ429lPTmdTbFwXwdg+6gUkQ1CThpwRUPoPo
fh1Onp8tkICpTQZN1W5CJfKe4gVMrpVPmqXrny8nFyHe9/BawGrLrUoorGZ+v5B6QvtUAQexf+N/
6UGHb9aacnMmdoESlDIwIKrDx7RG8RCyw1WGPJ969KpcZiw4QR6M5BhC9/zE01ZW9hDReVczXcm2
3etWw5S9bprOu3AGbe2ZDJLloFHDufljpGUoVltJAIsftgblaVpU6aMYw/FnQzzMmucbVRQaosai
tjWpErT+9xOuEvqSBC4C+ZQjWaw+xqUR/ew0rUuzc4MQ4erBUd2uSSGO7OvV/9Ul76HNUhU9kMc5
jmTgbC+EBzfm9BZFFDU5D1lI0cFfVnObMhbS/gHrTi9btOlnL/Ks4OrRkjdipQJxlqwQae9JPafi
369vx6/r1g+GownvA5USdSXcJeUJgdHActf+kpdY642ZizsAPziBV6sIfaSrkimmTdmO1vhrYGLz
bkAIXd5fAazPa9Fg4E+b9779yb8/Pv0eaSnTxpsXvRJDByeXWNuXQuW4qfCxLGsVpTms1BSvO/aH
7GNtn0YwGH8xJ6t277E/1uGQ+K27ykThF3NrYBcSgPbaQPckLUkjqM7HozrUNLPPNql2ujiEoxHt
bWLiPAluxLjwWEV/J80SADjl2iBzHEejl2y6p7NUjjWKevL0LQ/DpB1yn0oj1cZaPWd0pviMrjVJ
cUChZWcfBhf7e9j5GcTugWXWrG+TWIFpALglcJ+gMcYvyqSqfbmW7UE3rIIdk/5iIVMkxzFSHhYf
Kyjn2PQJ2UA2dJDRQ3ZZPX/3yVbSltDueaLiIY2fLyR9AXthy905M43Wo94JHfwvfSFyJNZdQQ4d
sndj3nt1Yv/PbZbyb4fZZDrOVL3mzu4aYzlkRQP1Qad2UVAgiyCAPPIFp4cyFj+r2nBEtH0w1Crp
GWnOc56koTchoPCGSKIz8gfRB00Yq1dysVrg4aghl301THjL1XIJhHW/p2bQfaod+91VAJaE/LQa
L2pDyPSII2RWDBlqo0KSOEqQlpEUbiDDfkxp+SEQt1MtpCIVMpofvkfbY6cQYNe8Ztc1r2FPxGdv
1lQlleUuXfv2ulRR9nM/L/Pi4m8dYk88aCbutupYQfx5Gb4bNa2wxQ2+oYZyy+X+iPjVFwB/NzAh
xY0HiN23Z96GmFfjztJWEl6R3XDrAh+I9CNWRMCzbfYtQE+vOvP9cMrZoOzrAcG2KbAbfdL4Ka0r
tMEugjI1z+fykp/ew3x+onT0rzLMpGua20mVrOwGS1xCg+XmsIg9k/7sYcaV5KJBoZR/21Uu5tMR
Ckyyik7zkmAvOv1InAacCKdVDGby0d3lO//q+9YaoHC9CVtAarSbZCtn1sreH3KKCoGQGFKMxUw9
XfI8CrRQm9r5oPviozFYm6KfD4NSrWG+kJPei6FI13Iw3pqHclvVrSyCNJVPuXAgqRJXBlgPrPC6
E3r1Zsvb5Bk1jBrfNEOvIKrmfbnOHO7rDRumlpSGDqVd3FYz42Pu1FAz8YYj5S7vcMmhSHoCRKs9
t57EENthLYOiGc6SSiOfzvuvipLzBIh+q5K4mVZeNYL7253As1JPw0dfnCXUHNTzQm5Rczd2WXvE
FWZvQaqZ60wn1nZqYyO9z+LDUqIFkLDt6Z5Pwa4ugrw2aftvNGpMaX/4GLsPd0LJLPNoclS3oHAq
E7m0reP/YRF2fbN49rWM6+YGbxai95wyEqYRPVLNGzK0YWHFuaDyC9QXOqWFAQ+U7Y+wLawuntvW
sMFHcz/pUl/+/f0IYhLaXAlAFm4VXdl7cRWHg+mAf8pg8Q6duIr3UMMBUlIDfIsSrmkjEePjMObH
0oBhFXC+7OoMmZZO4UoI97w/XwW7HJIDH7YY4IyGGbwpg5JUzTfeNfG67kG47CMV7Bw1sO9jUrCI
wdycciImZp/CiS1p+igYu6fgvqCuMDYf73P3OftRvSKf8L3+sO6qSgzOz3/wGNyudAZRsxLxcZcJ
JIgPKF73zasHuPYSgxN2xq4jN8CvDvRhsDCwP/watwAYvHJt51+5zCE/MEt4CNNeDgYG38C3Um3f
j8l6yMszPc/0XYlVflL/7XG8c7lgDSMnGd/ng0HeMODqK+TlELTg/Ja1Que4QSHv8Yu0mBgQjbQQ
sjCj+jR1mVTnhaZbhTRc93AsEvFKYMmCodBbLg5Z0ngqEOeBi/BiQleuBUx/UIuUyHavlJ0BilvY
9wuLpJw9dJ7BqC/NXr4DzFP0pjr6R9u34Ue+P4x9yvYzmyvV6G1XqMOZwnJJqGkl+9hhQMK2Ya4Z
19D9bG/VhiJ7E8sJEImNoPYC1wF7wY/GhDVXiA2QmRyuCXE3jIgUHu51JYRyri19SpI2eE0awnk6
F76zEqE5pfPmYGsfv1cjze9tB42q8zUFViTjsYwmZNDecOvUHxO7l3y/U53LDUHL3zDOqJzV1F9g
HH8I204Q3ii5us6kNxht7PncYY1q2QRuqLVUi2qqcFWMoch1JpN9MJaP9g0YNTzWL093+x4vdeHm
Cae2/QN5SO050jATaWT4QG5sNT1FoOHqxHzluZc2y+XQ2K7/P2kmbJoNl7XZuVs4u9jlj6AdtA0V
8funUe+yPLe9xK8/+C+XmGPcv0Z8bYt8hvDfO4qChc/Ar66mGuWwv2P6uYijgoVqXIdPD+yqAb+p
0ZGWqKMFFAq1XVj6BupCPkwdDM3BD8xKMp9RKRp4ohVIcHU24YlxbBYavxeBzbyiJ/hbE85/tM0H
6HW3isgk7GlAIgato6iP77Mq2OHf/LcF1O2sWYmbvKSNG32MkMwuQ3UnCq9qG5m4oMxG1RgdP3AA
ziHm3byIex4e3W3mywQ2DbypwSsFXE9ChpawHFacLbz8+zazud/qbV/gYIEBOI5J7vwYqUcFkwwC
2OLswdI/mn02Le7hczxentzgGHk9FanvcVmIRohgYMljMeV9kkOQn4uB8QsNp0kLctb2hNYAK4fu
KbIQ0HRjDtA1gi1LiG4cVW75QrZz4Xy0RJ3TzCAE3AnN583TMSePZOHzsNByc87REuXcRoGJ1WKK
zloIeCP0KCdI1CQS2Gq/aWcm6DQTAl1jE78Yh4wCtGToM6Z6GUca6z6dVzQh6rAnUZQz1tUve1DB
SvKvwenDpnw6Tfe8T7OxntPXZEB9l1JbH5G/NV5LvmGPHimcUC5R9ymVjjuCjZZLWjuAjk3lj1pD
WwGuqhqV+Tb+zz1Bi36ckK+sUdbrRR1IYgC2we/za9EU8B+7addJa9z3NAwopxW1czALV2lKbcfO
ooBJABNwQKjjlik+aJ+/xzzud9CvyQPqTpcPCpqF1ua693HMFyX69ysKZ53kK0370xsHLcW2Gxxy
5VpghAEArm3ZGIc2nyGMdZKta3MkRfS2PJ7n/w4zqq4ks1TpKaYO6NDyRqP23aRmvyJdEORH66SF
hYbBVktHvqEUqDMCaqvtyXZ7NG3A3i8RDdsZq0cuuVgxO8QdXxvlpUxC5YxF6tRFpEQamq3AdKZX
1ob1MSXOq64teON/8a+rJUdoLScR4e6+m9tqMbK+c3MymKnnSy3BcfWkD23qFir2B7j8z+s+/WiY
vEoSQHnDZi3WH7t2aNlPPAJo0ZZyZsXD5qN+MxifHLUnBlDgVM/gzmUyf1R/w+gfS8QCNrdb4wu8
ym/RD8wLG90rNpiPn3TnSib8QyaJz8dBvaf1b+Q8pndEvOrzfEIj811gHH+CFrezLIUW8geNF4Zx
6HQUa13pEAN4FhMAVcCla3DNfCEP85qde+RecxfKv67SKhnxGoCYsN7dp5VFew291cPXUezPG68a
55tFcvYAiWjBn2PhfycZkCWuaHxHlTCfcIcX+2JyNbP4bh59XSojWzO87eP6do4Awuph48AGW6G8
koVPvmzoAd+IMG+diw9bw5dtPerBFJikQvqj+qX8GTaKxOL81D++eRDOk7gNgCbck3wLDIFQVFWS
Zw09dYnioE+5EDGZQSjAlwS8x+pSRMxzxR7VEvmg7Td6S9Xfn0KbC+CiNFKK7QUjwNJIHMDdfb6f
6BJSm5TT8jJkCep4pEnBrF/kTQJ7km9LGvf9EA8HHxKwN8oyGyKHtfZnMjSKnjt0ZWWcntk/G52+
p4GOYEdeLTybTfmimk+dNk71VjGyGnvxjGi5Rz9/Ff2Kz4vKPvDO01UUPG1wSopMx8O365SsxNnh
tXekChts9mswWeMkmPvMFOUhJM0+Cfa+x+WZCHYEVS1xFu6Pf9HdNLLfVGUqtzqKaWWt8Ji+mUVO
fEkO4YB2AcmL/Se+9Bjv1ydpoq/EyFaO5GPbhLY8ND4uifWJqC2xDiGqLk8dHy9cbmwbx27Yb46A
XOONKh7H3s8z6+O8+bk5YfXHCQkxBqgh0hMCnJF2zK0qcWQf/Tsv4za29D2c+ma8WSTBMHHOwr5o
qxkSUVCdkA/NaEvuY4FAsODu1zv/5g/mAwlOWfqveMheXZgknuDmcyGbPNWTS0X45mMRog1XNTNW
IQrLMKZGNrWYuibkrD9yogXIIbJyhnnOcPzOKJKrR47uwQj/KXY2OSaUuA/5eBEJKU3c1p8iX/D6
mvxaKcwaDe6YSOedp2JgdhnnNbamNoK7oXDpWJDln9uL35Lsk/RaFprtj3Uxaq8ODW5s9ZCWuFFZ
HrJQitKC59+rO8zfYIHS3PYJkAwfuScKmcut14l2O+kUnD/Fw+Q1olkrnU9SG9m2X/wBWsIl7j/C
MPt1AWAh1G0GIYQJGKXokYWDZXDqv0lndHm6QytFbliHE7VhBmzGQIpOrh/XMlvN/RAAsjw7BTMW
Es1B7PNoIO+NOlyxC9iRscayeAtHlWRJ/c+OIGmx42ni6WoiPamp6ONekBO4dNvyEaLDKB9v/boO
HndNvky10TNSajCY4Blexlf72YIEAL0HFVC7TUiwZMwVGleB6io2Dtl8vmg9NeeOYq22y8m0dc2i
7bGE7VofuG7mwk8sIxSoHZ0Gv5vCC4EEEsp0/UJpkQvSfDeQcq2lTzVnVc8O3z153mbOGqEdQm+U
mAQIE8Y/dCuklhzykin2BCr1FkbSmG9mH/Jp3q7cDIxc87aT/3wW8bYoSL9RAzUsentwDJtVtLbK
qzMA5ZD1uzXfKS+PlAR0juPt00uuDYeXs/JGTVRYgo3dnXAa1PkrYV+OhLyCs3HVmmZJjAUiDvMN
eEsJWWiFRKxlecTPcQ8fqyHxCf3RjnjQS4DFqx/NbPzIphF9S224QEMI4gYSrAEbLOR4udd8w5o+
d5RmG6KDaDMIcod5treKxvUbNY5q46/gb+AA9DWyq8ln4wd5zWkuAruen9RxPWZnciNP873rGtot
dmmaJ6D4xLVzR82KLKt22jnIv/ws9b9nTNJFZA+NScM9jIXJyAgMy5zWF1hu+H+YKBIW5v12ZUqq
nWE/uyGY5bZGgWu5nLdE9B3i5VTWN5pE0Abxn9AUUF9aTmF4gO4eD/MHqXS6wCGHtP9mr8AtUFuz
OH15cHhkBuKHTffz+CZdcBktV25ThHKId+8E8CVVCruYnnUGu2fd3gD+RgYiWkkJ3/WVUefjtTa/
6F0U1DIkl3cQ4yOTEcV69dptphfpgDeofJCh/q28vXBP+yOLeHLU68wu04S/DftTJhCovm55WK5V
XmkqxZh+ks6mYaUJhRFrQaB4/q1BCeHJAHcxCIB1k9lfkQ4hw9O4Fa3x4+iygYKr96ZL4I1h5P/w
piWIx4wdFrBk4gp2yKvjPfwgE+kycYi+egLpBuFRhavdQcPM6pkNufiHvdCp/xgl95LwawHp1Ili
7skzDxzf42lRw1AP//rh9CvL0ZzZzW7Eol3Lopepe9ct/Y1qaO+1oy+ecDsjCwtitOQMxOJCgRNm
//jOEYi8fIx1D5TXeB2vCbzyZMJK4vYTMXse2MdNEUBZBJ9eLFA10GVSIgySQrSY7iktoK4c6i9a
ZruS2/AfdJHvXUw0ru9xPm7SzoHDT5k518O4/ZP+3LGnKVZoCBm4OWP9jrvpI6DtgT3PbteLgolf
yhkJs6hqlICS9BFFxfZEBoV1yajHXRiE1S2Ho1SSgkyWbQjKJ+qxjelI/UffTlaQbq6ChI5Fky27
u/h9Is4QkEvVvp1MeFrCixaZ0g02BPiNXVPr7hr9gzzvotLcO/ElExbWxSkBQIGxw31u/gSuXaTk
wDBS4DtLMICMdEM5XPI0bY3MV1L0IirFfq5rDFokyH59MafHO76/lT1lvAczN4Fp3NVizx30fPSF
17IcnEmKtp1doqbIRdKAS+U5KeKLm1FKDUaxjqElpybt42ofusirfZTdY9KPYfy+3jTww8WNkI4L
oxJIFsWJbvZmRE2m4xC3pQhTgrnUFY6FRk/NViCOcE7uj1vofy7ICv2QkZCnd8oWFYSpKZtuEmvC
baT0lWAI6RhTiVZRf/5bEt9BmCmm2wiPNCYoL3JIh2dbMn3YnK/GEIJa4fDqyMfiuZoZBTXxNOtN
ZIkXlKJU2crdO5doJjDw7wUlb558M0BCVmhrr8AxnmDoW/Zyolh/j7xxjsAIMjECbObJQjY/qcpJ
lPf4slV75PSuLky2dNkR2KRWu14NAjoyHRwKTPWLSbtYe3NqXyeO9CHgBTxJgH4KwozDmmrXsI5B
s00yYJ7UkI4ONxLHtn0ZBKOW1lb/BgxV0SJridMubIZQLqjgdmUDPVoqNEfRRIIJt33Mqfr1qDjJ
+w2fj3PvTYZ6xZMgdc48hRaY3kflpoXmCYO6QeOF++Uk3hjtiCN5Zrd/USEM3/B8qzv2ftORmEPV
xMocPj5Kh4F7kjmEbpn6q1bMJxXIG9rKyH1R+uEip6n01KksXNP1F87db38WwfiwERG3UbJ1g5BY
5qtPlqxii8BZWZ+77RAh5q658eoEzvr/F/K2SHW0Bi9N1T0Fh2PKLA0c+54v7Y8td8Gjc77BsciJ
XkMjq6T28e0R6RYsgmCcQaHqfYdi1h2r0FuyoIPRYA5sjydBeOo6hpBByJmQKdYy1riO+BiO/mIq
gAHfl1JrxnTiRXHfELQ8NJqU4XIfHYVo2l7/KyRXB3QVDyePVj7rb1ggdJ5VWn3B9+gWI6ofZlN5
BgLpUQCjNcq5FPxwQ7XRUE4mttOn8Gws54uVbnUQ1ead1B6+QWVrZwqDVNYC3f0LvZ/CuVI7Uv/a
RRzfHeCNmH+cHShDqig4tAEpZPggBi/cJjrLrQ2cPD1HXtC55YCDxwMVQEgwLT2/hbek0kWxUEi9
yGPHwoNnGJHuZ8U1Ej41yyb7smAx5jGztoNQ7sPuRRjsuvTQUtWmG8DdJLxiarJdkf9oSx2PEcrl
GsLHc5ZbTMzeLmMwN2ZE252DokHKf/BSRpJiF2kfj6OyWv8mhADPHd9cf/0XJkZ0SxcqrTMR1w4V
VdZTTvzYHGr9P4igsgUmcOhKbEd5+YnfqqwymNrFiCKnUL6p5+/tVF7YiGsm2/+jZ8um1EZBOjPo
qOSyh6a9EVPlfK1yw+36bzS5gWEBMaypbBE7LVckOB1pNxM62Apv8dsCFEhKhg+8PT7umQJ04iZ5
SF4afqgdt4kLnIF8pvc8ZUkozew4zcVftiYbC7pdnlbWW2+AelnfvPuxf/K2VrbVL4PUjcDIiefC
GUbyXbBu6DrId8VwjW0ymlhZJXmho+fETQ0AjQkBBTiBF5COm5oCF3+3jGmw2RzrDI2V7BsnCnJ7
fJZCb2CXb0t4LGAzK/XgdNYsSDfEAmjDCtOPpFhd71TFGgwfo4bjpefqTdp2lm8yrUu0+i4GpgH1
4uaIhBddEUHGDUgJMIWVytruTQPuW8CyFf+R9qjcRA20NmREaYlOKCDX3dIcllDY1s74EhgjB1jX
CjAhe3+az8zM2litB8VQbF+YpMyuIuAniCzPKum50HZrRKs7NItV5B/FlUnapXE+BaGc0dD/TQZG
zui60sCfPrwuCrSaydS6NF51Pb2ZpSU8nzN+CvSg8jpCwWP5FPxDug5fg8M4mSNhf7G9eaKSY6B3
KzV5r/QI7vZ062NS7tvVO8aJXCNueCMSzMOMp4dlNo5D5gz3TI4wEqqmqz3Kp+PFNwDQ6MeCP63z
jzij1AzWEIKQPRbRzXyddXJ0YnGfbUSU/vrLQKduZR+txytN6qJTNlVrzed+Ck6mL/QQF05usXzg
FYaYHPxynz/oslVGhtKde4V51F/xCWqpPd7JpomV3FmajlzAyW93lSFSFukBtEOKWKou0JG+u2WQ
KTHKLIdV8KlV+iSg6i+GiXw3vKGFF1TFJNihI9gSBt3C12oZGW0j1hyaCbqqNVT3pQvxDQkiz+Ri
meGqwisuxLQDgfZTJSCUqVvH5gzqKA9A4/f10neNXzKX73gbfkCTpA17SsMK7OhsyeIPCBmGEqp8
MBWWdKhOCk0TExWTChDy4sUm9n7waOQQ0+Q5vD90T7Q/Q0hs8PRro22AcT5ApaccwQAv0Dm16LuN
2Wy4oK7zVGjfmAhnEg4A0uSyZXfwtkRh+Ihz971uzpsaE1AWibJ59qbx24h/5Dzw97eTV+c6uqNA
iIU6rRnjo01TBOQLeNvzi15hXnafZR6jLLucF4KT+8GLluboE9R4dKwn2kV0dKdkpqDxGYIQ0WSn
xKqZaZQT1xjenq6tlkOBlK25/aTgiB8a1YRdBN3MBQsIenUZqVhXrq+snGQNQX8PEGFARoJ/QIEF
gEeD+UFav/eZIbOoAQEb18EAVXFeB/ffThRhIfNf8EVMJ0yLCtaD4VsNNBP03Puz/avUaLqCDTgF
mP05MVlopMVQ0nIfts27OvPFGYuLoSOY/hVgdn6K9YJaaJIsqVc1vV1YAa0KObhVY9PP8iY127Af
WxTMKec7Q0RuRDvW3qZV8YH/GNO5sygpVMK5HwZog2TRzvjqbRRMP9qPFtzvh4c9CjPmaZx1082Q
aFrczD3ALRiyQyGM641TYUIYwcMmPx5yhMtPyYrVDFeh+fnuSuTavXVng3qgn5rnyGXAfmruDapS
tQZLdUrxk05O6dJfOMsnpmZzZPTdOwirKF1DYRwLLoVE7hvT041cAUVZTYwVoxLBMUBynYl7Owrq
qfl9q6BewiQHghz2lKZh+o7wWvkCBpsND/n8qFe3iKDDg0ME/awHmYeFIJ6eb1TreLXKYH+NPk4F
5PVdQAdLpgxeQ3Phcs4OG5rpGF8xLDz9MlXjjHJkLtBN1XM/5ckS9bghRz+5AQfu4EkrcErrux/q
QQWXq7xVQUfVwK3m2sUT87aiTv7ajflh2ly2upbY0worL5iT3/Jl3nsS7NqJ2Ilme/+vOP9EM0m7
7kvhS8AXych1r1Yk/Jw8VwFwnwz5/9Mk2hh5anrADMYxQ9iykCqc7VALCd17XaD06JVTFQprbHJR
V362eN3TmFvJI7hUiJIj4yJc3pJnEYmy3TmPSKpMRqxnqcxPk+vDfzGVOpK2153oVTN4yakgW01V
bbROZgMKIyPVLOaFOgwZjz7R9B2R2IPmhAnYKdLXfVNcTAbNkPOCPsYMxvGa7LS0RCUAaMLldBvN
X5KepEICsfdRMHIZSQcU8yIctweSCN/Ti8sPAaVwuLMVxLZaK7l1Xe71grLAURFvlD4aSqJgTB/h
Pavbz41gEzIpREIQpuliqwzA1kBsqF+rP6RpyhnIMSEXbmJPk9lyFBZSidQ6u4l67uWkUSe13WjO
Bt+I+ABLqELnc5KBY4wq2f+KD5acaIV2YEwV0AVHk159evs3nEoXg8/MN5NtbPiESGijJt8ndzNe
TRBfk36DYbK1jSKEidUUoqT7J2ivs6OiXHFNZTr+G7llaxRXP4Hfo2fuNwoXoE35pnBF0fBNo4fP
bbtml6A3RxNmJQe4kofygQ1ZDkmhtO0+81MLIr8U3Wtw3jPsGxT7ctkLKSwCzISo2OPKBj2639j/
gmFjSEcOq5bYIlYh9CEkkE3cBWrV2crh/0d4UMy4WvcZ3lG7C2Nd1iBRV+UZuzSkj+xlE9xiOdFf
0YVlzMInQWVqSLJw1mKibs9GF1yt2aBHN2AAMQfUzGOcKQi0dLJ6YuPFGM3FfmqHCrebsrZPR/+T
Ywr8ri2iFeKEumu/wxaEfwogVpVkBlDzknwuyr4Dsje8Gihnt6Ak7Zz7tXXHQkEWBpDsBbFIqsNU
tvJb0ghfsoG2gR8qpiT/HT7wcXUZ5RJBxMkwXea9mfPQR8NbNchPvMRc8WVn0Fv2WQ29j5djAC6x
kLVNx/IczHNe02G+Rewrk82HAlH9/SldV5wrZDracDVGbjkYilCeP/AdIphsCUwVRpJUWIMivhqi
mxnHMESD6b7kyL+TFc4oRFfpirLfnQXqIOjM0+Imw+t2SHvAJkcAdUL4YgggDNh1NhGWOoVJ7g/Q
bppQAbVL3CCnq3Hul6p1I19UxuNd2m2uwOfPp96ts6f+1NNzd+0/4EYrrbCl2CiWXADgZKsaFavC
oD7HChANeh1el5qAi+1OqKusbaNZKMnrdbY2JK8uKv08yHgVCfLVmcNW60ws2dNFQyEYYBVtAbfl
TjoXZM2KDtbyzNga4RGm5hc1NnWMzKx04ogpFeFe5olWBehxoKamo7P5iINHzCqzfQBZzNI0ZWKn
LD42pAs3AdyRUqz4Nd5gGf2lvsFw8HIlXQe8JTrG+kB4La4zxGLOhkcXFABCUDFHcrYJvvOgP7+l
f3gt0IBwpuUVGotyV9fAflg8HAZM6cm6LJGPC9I8RaGYf+OQkwM/fb4gaFL/o8x9ZuRtU7eS6z5S
k1Qt9wPq7kRZgrYBd3y//CWT25BjOKZMh9PJ1ADNJHDsJ+exeaoGqbwab82CNi+tEjYjyPe0Z0Oe
qerNgeC+CVBS6pJt/uKGjK/L6k5rd7/FJMTAVR6CBkrP9wx1T3sLSkHFhz5+bRx68tMZdsEXgwkZ
HC6+9RXGwjvxlv27R5p8WPcj3He7Xf61RBjgi57uHs8UfooR/sLTx4gga0RgoQMw1m3eZZTAFMhV
CGMCvl6LuwIY2rKsY7SdWLkX5Xz8veSU67qCyIa61OSL9BeeYaZ9AnUOQjQMID0FEDpB3S6XpCZQ
99d44BmeloEBoExBLJrycYjX7zEPsWBImtsaRs+d5A3I+SMGX3Fgr9UM2RliOeUrd9PHK6dJf3xV
3wdj5qUXIFwN9d9znuOimfAOlg/2PyVslccHSsCxygb27kCTzHGxWHYQLPkj0ryn+i9l1+8DVufH
t4tQnKRknC2tvLFHzmiUOkQwtCOhxJZwgsC7gTvErAT6a/qSkNn0a9Y3PWIKCTickW4dBY+OrEhV
hIuqOMe9OQLIEcm+1EQgypOVXjT0MI8wxU3O5hWttLooIThqfn/eFeqr64zlN9WxJM8M7z79N5PZ
Gt/M8GbxRfDOyuVzw8TF44UtYvIbuLZ5gUUD6ZoH14HEjtG1mAH0ACjoWUu3JtGaQ1TIpBs6PR5T
te9D9RqO76sEPaPiyU42RG65Eptv5O3qrbEjooTs8qR1lHt5DMw6O5zPvK0Rmwi3wh2kbolQaiAd
i91Mfy+qgXFA1asqY2q642CUuFojLDf6UnweXCQ3x7V+lanGaOO4+QVzawoPzkajvXeZ7EvxeCzZ
X6AMB4p3CAQ5+W+KthgryhR1jpCSnWFx1Hs0oAkHaA0mjpc+JU5ILLu/+oO7g0vxmG3wj+1p39GD
LfAd9t/88oYGIDFZpReTpI4ARb8cZE/4Mv8Qimb9VuCz+Ano3RLqFO/8bncrqSDpsB9HPiH8tUr+
voRfhS8b0psPF/D0fEakJpfJ8Mzu3HLQz+OIUYIIR7QihrcKc+37dyTW0NqLU/UqqwzPTvMJwAS4
8FPrLlG8oHm19c5/OxtJKHRrp6VerfQos+wR0D91Zsl0z0XgwJ+egyUirhef2hrinOjK+yZHqolC
vtF4QAJi2IRxapImQu4bfyHqP8W0Td7ATp+9bV8+3JUm58YlSYITNiKYEt8K4RNXo+R7CNsYEgpR
KPQn4YNaBtkciCiRvLg19rHBOSfoDl+sKESz+jyVyvma5/vJJUQIqIkSbdIxRlAb2ToYgZDZ+mlB
I5gyX2HGet4jCwJgEwhIBOKGz80syLBJFcLMAU/okiuwDGgRcVKiiBCDKQRF1V7NjQrh54S1/7t7
eBmgQBFff+aXfJzjXDlQOuOzTM7AwxdldAI+cQVp+Adc//NgyjzI1DF4gYeWAgjrRGzV6kL698bQ
y9jbIPUI+ITWv4vRag8qYOkvu3XWybpN1GaqqblO0ZlWb7Orv9GUnpuQoF+qJX/i+fiIjWy4TUTr
RlP76Cb8PvS1sLjwTMhS0Ob67cEzBbSyPOA8KkkVxF3RNVDlvNW2kEXmeVYJbZaVMkAyzTvnChDT
8MXRKac484XwV6MItyetsZmflxlxmHxZAH+rkF/wB0xGAmpv31flo1lLY44rPpb3qZ+8TwKXefPz
J5Ve490JzNd5brUAD4ZsOsV2NJHPP4aFTiUnVcmPEt2C7G4zjnAwz3g+2N4cbbGfF0DU6O1/2Fow
p0MGGCfA+1iyx+nxKJ4lqdgRMMDggJES0vI/Mhd4jMjB28Iq/jFeFzZ4K7Bb8wiHcEAoXQDAX6uy
Ol6BsXmWQHz446ucLWDT3qTFcxjt9NljbODgRehW90mRnERlwd1E+nruK7FcRUWi2pfrpfnT+edy
7aZOvZ04VoQQrp40awHnmP/agXVBWJWJI80QDgWPqH4ZRr+uSffN3kmoSKa7gAcnRGIbQIBUcxKe
q1Lx7364CUrhGGZEbZp5goDR+F36pGTt3/HPc467PxqaysATYX0Jw2N4GiQkyVh1seszktYsz3VF
aprq99jSDXElILClB6KYJf52op1bFWgB/thRL0klHj+hxoqbMXO1hguSmnfG5UkbA8bmiY3CTvCK
dnszv5Rxs6AA6u8y7/LMGnjNhDvzjQrFscEmp5zTKvlhcPEHsIFU/dH6EagNlAYL6VgWGPolkCZW
MLgBoVABLEVyPHQP1pd7tx1g0ooBJFi0w6dX8FrLIg4VMNjgI2x3MWIq+RXdroBvT88WmvJFhU6X
f1V7Oc8cWMzgupAGP0ZECpzRM17zZVXlY2St/RZOIvAnIL2Hj6+EpAtFcShej505cp7jWNQU0sWu
7rX+zFBQTRj3kw9FsMbbLwNJFt4VpO8fl6Jt2ZU1qy+yhYL89F78C2YUldqPQ8juylFTQYg5ea78
AJN4S+1hhpG5V+ANrQGgRKzHZzcr3GqGTfOxY1wwTSYfnClJaDgAQNiwZr5km8r9VHDxSlj/5CKI
rMxvyGTtfeu2yHqPq/WKHGptQwnN5TyzTV5OxGxYTjxXiMobnI32RkVhyLlVkI52JSMglVgipGOO
XBKkrl5IDOF4bhKMtZExUH3USVsDpc3pZRYLUBVSCyjjOpzhwEYlFgAd4fclFyWuphX75VP/SnCH
MhLMmb8OMe9m/+M7Ue3pQuOS8f5zQVqoD4sngGWoUm++j9vodzol4S1K+6lXLJYUuv1pjQ4Ae0jp
8Qoq//qi75TtZUKRR7fz9lo9dhAnUNeous9AIhC9Ysa9JUVa0ghNFEtyS7ow6+A4YlkpOnE4nfw0
gyp/CF+Ik4qgjGd1cC9YHu0F6dcBQ1SEtnL51iDDqOMfbIwzB8s8qnRdQ1eM8IiY3jxcr8B+Rvdb
qVHFFur7mATGI7b3qbTgb5xgjBLCQ31Sg4Wocxa/LLNWv4fvmqstMwHPRhliH80xP8pklH5TyleA
iOMTFJO0NDiAq6nH0iQc968zH/JWuRDieU4qCHnsxdl3Eh+9Cn4DmoMd4Su8z1XekVNitkC6aoPf
xWRXOMYDMdgfvpzZRYFQD7Oxo/mhRq+2DzyKskYdLF4vDf0+volgCW4FfpH19GW3cFhCQ5YdoyQV
Sur6A+PN1jb/stbhEBPYp+l3cNF8pBqUp+FjqX1+u9/Sgoucg+C9DPoMBXXp0kDm2qEdS2aM3ip9
r2utjjmamWCfTv+n3aA7ZU0BK/g0k5vfY92qJC0BU+idG8rKG9e22a0mzemkzhw4ykHBBLUu75Bb
+LHt0yf8btYTF0zdHKrIDzuN50eTPjujsLpStxVfH2va8LBpsibndBdITKlLiKD7Eiv1S9Dw0awP
b2gWCMvJw9wD+9curXtupDQ1s0+21OdT3DKCRwYRwlYM7ct/GfRVIAhzuSlY9hPY0egTVX3u5Nr4
H83dVlWqE8y1ydv33Ts24WtSBjOFFDQvcqyheP2Smn/3cLpqn/jfIZ3Dh3sErxoMC9jlcEfvdS+5
rlOOzV4N8uBetkTw4Tl+/pmxTKwtP8KL/fFMasuO4PHB53qiROkXc0EhjGytWzOr40tKcU2kM0J+
uuKX/FT/xfQ/vNBNEqsNW2hBL/ORInm1A+iBr2J0GMw9pgT+b+QKxPH3OdbXwpI0EjGY8MspOAw8
kc/5i8UqyQh5gLVXjN+1SK0868/xWlKS6g9XJUELahydwzcvrS/GYCR1RijP+2biSHPcX1b5Ua/J
H4AzdvYBj/bI/A7zYLEad1LWkeIQo0l4lbtezmCWaW3HQfs3ROu/H33qK5++2cqYCS26urYDwN79
TBrb/2dlwf6M7SPqL1q3uU3wR9jeSWeXoMotuOf+yLjnF6SXyapvEZwAM0zZjilHmgQQFQyW+HU3
eq5QPJYqcWRcAXgQNmMacIBPHEtfY2M6ZJ+bD4Jogl+hVjX2YyPqIb8VILC6Da0KxI68Kdx9vZjy
Qvp1lom1noBCaF78xYOITU4vyrpHfwlO+6CgaH2buIDlbeF6iv3lj6QUwS04wqdqM9blyjSSifd2
9wr2XeZl7OuIhX/hL+naQDvT1JoS/9O/mlniE0I4PBSkGwNelmPmBZONR3PD9mCbBHnZYuorlUtP
epao+8p+oj8dXW9fMr3Sr1vjgJuJNFe/67kgqBgtJpELQDSzEBpRY1JlWXBth+8Y1xaWGj+Pr7AM
KWcEbkxQGYokvTFf+7myLMIeAPEY9vnY4W2SSqchvEn1RN2EJa4xHxs10Yp2rAu44rTboWn7ydas
6SpKnR7k6hM2g2A4Tg7/zaRp2fhmNKeSlhaoaZOPMosNEWem8cmo+J//07gMoBXZ4ksfG8gLfVRP
2ukupnuGJC5rnNn1f/3xyhxb6mqXZiBIavDWUeNaPMZsbbtpiPl7Hz5rLoYVgP3yEVqNTuYBHF6V
3txDPPTtElJrGfcunatKS2abGt6NFICJfcYuzr57mjxRguagmgCtqTJCi+WyqVSxbLAjzs9gkK8v
bkWMX4w6CZrpGSveAt1myDGhjNHbBZ3lDRN89AbggiER+ESpY59bsBFGVgThT4MF42xm/5ARDy6M
gITPpMMud3WnYRopXtE97sOYnPpC1asuKocHGWlHma3iB7PlQ8xVK/1kEq1dKJyrbDEdlmit6SnQ
4LFgwCwSht2yfiYIhX1HIOL1dNeroklYxkXEBVgRAxW/UvA0Pt3dcKHKcq7dSbDKMSXxCItn+l0S
HAwhcRI1dzH9L9FsIAVX6tJyvKvCmMXeM791TEch52hl6rF3TGKiBg+WPbtQyGa2y2YIxAt/rsWy
Wg3x6siYCU9YgBgxvHBqov0IHRCb+0S6UresRoUJ45gE7aZB1mHlSOnaql3aTL0qqLaBkuJDMlz/
897Ma+eof0cTMC40ST0tsfMvaLNzaCCgBFK1IduZJ0LRnzGx09RBuZf0LKI0+Uh8Go4iMUi8QVj/
JRAsXUQUjFfl1SkiTCBltpM5WmRfdYd0YyHnp0ff2zH5ATFiMA2UY5l1veGJ6ZZLvLTOrLr7WkYO
NBMlO5N87MSNEVie42qHI+5M/hKfCDKBkSkKf8Z7A+JYi4HW/78EYw+Ou6JCCF3jmDnspvSmYbYx
RXSNJv3zslWLmV8fBAsGR7brnqRq3xV03d+dU4tlvFbNVCoOn82llVS/a2K/lpPK9QO3axmFdEk6
URaq9govTiOKq8jAc7ITmmTmEmfHQ6cElFATEFTtYGsPN2VildZ+Q+PdIu3Js798EWI+6xwDvSD2
RCc1//2fOlMeSVCTd73ssrdfd2gCl4q5klSJmknNEll1fZysDYyRXqhLjYOCSfqNf6OirlLOIjJv
8K7QyRgCbOWHILt8KtDhhQcanuRUeMLn649c8E0rqaxqtzZtECNXBgQlYVSbJVaYoJvJ8snBKTm1
blTvpAvWKkRGyvNoVWjIsFvOj+39hmDP3f+CHEloWNytXt9+ulNI+wB8HZN8iRpK/sVOOdF7qY2Z
N0xIrzyUBCrbYjG0c6SahgezvYv7mWLcDJrI+cES+9wYlz5qj92xltQFIne3mngZ/Zr6snnd3rJo
NalwUrpzQcS9nOOtCgRR6mtZVoEh4rrdk9aBPsMj+sY36JYFuEXCKKLZqJSy/JWpvdrp5g9q3ONC
sVAyKFOVrwC04a5NNo1eME0wNE/vyOnwE7mE1Y9sLYm8J4oohUFeyZZcNP1F2ekbqDdhbFFwO3bL
CUOnFeHXtrpmXRm8erMv3zzpDqet0lyRHL+478xSq6wvsSsvulWpbF3GGdlLfBJ+LkYAaZgeNWdK
eNqpOWXRTIzydN257W8UcGN+OV5VsnziZxEvy+0KcsCcnwZxG86/lIW8wZfthSoJt86bJJY9eGzp
3gjHXuMMJwovXkJhsUlX7/QQjZo8EWXE4r9j+TEmQoEMXPPWoFCo24WBzaD6rcMLr6PIC2XZ7W6k
kWon3tnNfDzzcaBbXxjh7gw/XEi2zH/8K+OGPniqhW8YY7+oKrSKJWdV7PFoSulAS8XabUrPC+Bx
qIzOqexz4HKkPNvILEdJuKZdmizI8kvxKu8wxzjrlLJnNaDJUiPh4zYY3pZ0iBmKLsL5hQVzTKyH
71ygo9zmpzcDNjQxHN8gjK4XqXamlKURA+36EP4xBsUYoowMN+xpDpBCgWdZxLv7h8/f0Q1nvFqb
eraMjDe3S+qDN7SqzSXySU/X/k5rMtVlFA/MPiITDKmZ7Wh9taxi9NIEiUH50GwK2iDMn19YLJJ2
ZX1NSdujFiwwWqnyaLdpFYHXhWdVqaB9xnh8ZRZKWZQ4qY0ihEioEBB7F/KV7wQoqexWQQq5lPUE
AKr2OiGDEPvQOv8SJYyfISK9ap5Yi8IECY+/oK7SJj//a8IfJg4xIB3oDGUHtuyf4KGezfkwH7gX
3Id+KbNuQYsUVbVYQ9TfAxb/tcbMiU7nBNGLs3iklsXom4NitIdyCc+jXgScM+kJ+esR+ccF45O4
X2QiqpfWZiW1OXrQhZE57YMSCzASgGfNlef/sNs0Pgs1SqeBgwRsnEd4OWIrc3J1ZvVkeviqKWs9
Di6thLKkDHSX194fud7b8GaPPaV1TjlmnUi/8dyanprUnc6JdOUFe62US8nxFq+7CfbrBCSWTx6y
QSz24NMj7L7+DR3apDu/qLqX8DEaM2VG3TnHBrP9XFlWxRyuUtxZjk/sfmP2AwI1aTGcTWFswtz1
Ytz2jJ/PbQubSZw5LFbLH9yC1XM7bjbzcbGw0ubDtazO+RWXZ3QLZMIWgGy5GO169Q8nDNvyXloH
jNC+6A3TTbKgPL4tsHf/YG47PT8j4zjmSGuCMlex3DYHnu++YdLB+GY5uR3rl8yu46K09JfORzYJ
MiibcWffH8jsBpm/Dx1PjpJTimznzMwK3u1dMxraqsU+p5Au3jVn0Wzw4E7NvCLMs5HgqMQGl3uF
MxucjtRp+0BZ4Ej4cT+U2WBFTrCs6RxjnX03+jRbf/CvAs5hgL5I77WhYgRepi5OKPvPJYXOr7sy
uZaw0Hj+lzfsin7Sz+1piKR6UI2vYi3fUEAXzLLDa9aOn7/htFLLnFlRdZ8WAHs7IhnVV3JG66P3
Asc8AYntHuP4BIyvEO0zYgbFDMHEBxwfCSC8Q4LMUWvRU7L5ZtQY4qdkLEXNNK24mqDw1vANPNWr
+iGjjxH4aHHuZeiZdpu1QbZZpuaFer0wpkdKRnSnftWLHU0nM0wieec7fUiSRZ6WZaeZ0s91lKLf
C94s1ljVslfgiVAvuajcPF/DbMHAAOXc7jZuQ8/+djMdDUarc/z48H/WjJNo8oDdaDh45iGBDm5/
ykA3IsoyjkyYSQSqnQjerZyoM3PyhOi+qBbwW+fy58MhX8J1ZNCYA4IOs8k1o9PMGLva2eYG5Ypo
KksTqdKxMppuxWlmIvSUx0wMLvU6mrQSGwjA5rn9dGbXWb3WoLHVUFOU94SMlvAYn6206XzJz4Lx
7zG2R2tIaAXP8bmoXB4vSKxWnQSEZioUN3uQPHeoPsfiD/HPjyH8ZNk4vO+Dn+/MVNssWDqFSk4R
x7paDOBl+UsxjB0YsuWFWjEufq3Od6pFUKMTiSKEMe+Z4KPwpLxDl42ueShDLSm5Lm68zlBDI8pE
K+0as/nMPco+x58+TXlnLl3L6hDTFJ1vjCUlMtqruClu6TUG7kG7VLd0CKqal1iNqbWLuSLyLKpx
VHlyJ9wo7aHs698XnHB/v/NLDDaxjnsIGI+kOoMTD0Kd7XMDrvwJ3MAJ8VlJe/3R2noN3dVHGqV1
jyMkm4xavzuObQC/AKhfgc40xE1k00o5inoO2O6XP9QGOJxOtT/iTrBKehuXvanUCJKgw4MbxiXa
Ai/TmRcTc3hZIyWBdgfIt3DS4v1nCbnZUEgo/dZFjEgphyWxyVqmzdFy4VEHuNFkBR46MNKVXRlQ
NTHmXLDkzQVM7kQxXHFq57+nJUh9RSxgEFdbjM+pguYe8pLbPfSDGKP8rBL6GLF+nmLHuEI3OpN+
p6vsVuhpwII6uAq76lMLEpG2B8ZHORTLxrD2h6R3eomdDt0tqZqNowaf/Qe6VoheAS1Shp8kA/Uc
m2WzpUmO1KWMn39gD8pXswLaMFLMwY9Vu+2vQTKuETRR8ntpRr9euALTf949292IgZ8wiOlt5Al8
dmVVv9DfLNtslJJV6qSCEMDOUUn9tUlMsXnBAeavp/pt2L7ivKHoDrvI79QsIXs60EGh+j2Qzx5D
Krt6p+dMv9tIExM+5IHNpUMnVKfEBaKtrkiM4iUU1PtUNucEcqj+uZrlJj+AanVAmO9szzOqexUf
E93+GlZX8b+EgnhJvkvMsICJiCpSvnb3wIV+uCMrFL8DaT6a9L0OPVPezujEvLyKWYDE3nLYMXwr
36dxChtEBuSXv9cOfiA4+zQ0QrOdtOQ9pI3WTPqe7IijSAekkVdQRdWuzgQVzpqDchGWr4PBRyJF
s7BZpA2IuaGtIRxefqqn52GVots676McA6F6fJzCYoFivfSs0eHMzy6iZoApYrmGRRXonB0rnY2J
oZ3Cdj2LsB7au6aDmiueQSE60zPbDdRo22nooNuVBTwXba+/7WvTiDLcpdUf2HRwRKYZa2uIAeYk
tJZstaWPwitOPnlkQiT/b6AUzwrP27JrNkopoK2A19mT8z69SGrchU0HQNn2Xa6uCDgMUG8p1cE7
Gpm0mYuqYEEEVDW0SvRPY0RUS92JtlY+5bc3z6fJ/SyBC1NRWPUurglzB+d6jiHfSrTG2PENahtN
CYn+PmbLrmkp0nq/+GyJYoNo/y1oNk+wG0oJtksL/tmOQG472PcOaKX8YeuXV9Ri9WrLM/2s50g5
3gnysxc8dEZybrruTXmyljNIV9hir9K+BDHOjw8iNrCKavyv/KgQck42qmTSXhfcLgz9OE4XgHny
r5gAZI/DlS7e/zcwWBGo6w5GR84GE6q259nCcPw1Jsre0/u95hV7m3Z0y7pw7zKrGeyVWMMBwhAr
DmQ5BwYjEMLpARAsJ7/lyacUt9w4Z+HHHSKVd0F3yhxrAGbG1un9q3njIhZINbFRHlYBeCoPx8j0
KLlMCZ4dbLvaT+fJ3jY7P/h7zsly4KskGqP1oTZhFewSmGe+p/0U2vvFb/uS35OAxREW+xUmqQDK
s56hsZLVvhzTiXlktWwENzrGcfTrRbZv9TeUWcDM9sNcPCdJ516lJPZvyPkw0/LOGOwrkkG19vMO
/vq8jUQWonlFsxhpvNKzCYSB1AC5TuPQtk+0Y38zNLaFvAGEHkKSJsdSxIno1luBv4mjcalNvwKJ
1O+YSvS4cikNJzc8mtvza+OCxF0+B+G+jaYT63/n2PK6uIF+neU6L2rdUzOPP2bvVzKjtsw0LbJp
Nnhsjbz92FuUJFTMJvKnluV/VxJI8hgD4BXV7nWaCYzr5fceuRpAoYpAzndNcymvpJkT45QYHsd+
H48uhjKaC7OBTn+/tCeSVuOwnxKO4uLUJaCTBo8mZMXcaKJlOrlBUgxFG3oO8UE5oXE+QN/Rftm5
c9QwWaxs03Y4Ve16d62nB2IaB24nXvnSTGlK0+QcRc8EIUecSpu15q3EtX5bqyS0iHqf5hwQOCtJ
aXNB5ifYxrmJV4XIyoZWKgQ+6Qs4bWUisrqSvY7Eul1fuZeLBeFzAzCT6RLUe4h/NMLFXVRiRekH
l3przefg2izUwUdQ2zJrrfKJ+m2aApYIqA/nDnfhU13iwjxzU0lfQrvxhkJ/bMqRltKhR2GCEeT+
uiqtqxx2UasPLhKuzEW7q2d6uXCPT/aHcUtaUG3xBkdOgTtbAJ/xxt+HHCxxfkuDHifkDQPSiOZp
v4b026kwzSJo0Ni/YS7ANXRhYbbIRQ+m/ymITkFu++UZOUEVwp5WX3dkiZWRy3ouz+NQ5swHdxjI
fuH9Vxt+EyWY+0E4uOhKaDnvQnHfpj4UQqqWinM8YmE7B4qbZOiO2a1JXIcd1nBBcJ7ZOyLoIZF6
vhLTc5EJjC2qDqUI8J4yGYriJ9BOmXqU5nb9IYwtQWDHPNGcyJwwXS0PH5JC53cPKArqgKfxsiNC
bQhhHFD/NSNZXhVktHv/DXa8wHQRKNXy2xJow5cG0tdz5mSTr3Gju9AJPjqL+O0O+JXMffXD2mzd
ineRedmonacD2/xOq+p6cNAFBHE1sBz3tL0aP6vySlPXkX3y99oaiBXzRYqx9sP3dduWiyga46X4
cLnLIQkuRpYyZzhmvLN/ERUbceh+gs06Kj0VT2sUUrhkkRo2nUkOQdSNNc6+Rpz+2cg/Zji3Tgeb
bKF0MN9iYhQoVh0r14CNM1fUDJpc3o2noEXbp/3FIMtAzyJ28Mt9JsuzDhx5nhcgh+zb04/oJmWc
AOHkT9F1hMrouILaodE+utDspCzaQ/zFeAOafoyFU4I+9OolxC82l16IqV1hPscvs6WgbVQuIpp9
tkyrlzaL49L9/7pNoSq56mUxRvtNK7fzU6OXkNfVeXUev0KHv6xz3L00eaCKstyYW7FOwP0SlH6w
93HwVpDcuyFWdzgdy07HbRCI7Pvdys1DnXipGkmpk7gnUezVOm8GAPRIgE9XrQCnhO6I66qqfvsq
2enfm+zQm7qbN80J16qnF7L0FoAejWSrdWck97DUMX5+YAAgl3TjOKXZmo2y7ncHxPRZ0noalJxd
FOlesmqZTYRyzS66ijFg+AxiigtUsMDBsWtUgQgWlb0EqVqfnMaZwm2EH3rWFsGJ381Vgfo5k891
8Kf+jHHE09Ic/bRp8m0QB/TUCx1whl17RIO4X5uvOXRmP4NWYqmII6aTC5ECR8KwYicWpsGlsStR
JAs32jC1jjPuxmBtLUbOnFXTsENCtw6wGuX0Yy9mJKCsoPU50zKbO2LYaavHnTz1NfdOuHuVDOll
n4+4rxSVrGiu8A5ov73nMzJWw86olbVU9tYi9KSnVS150UjUkqINOYqQz5du/qrRkRkN45zlGkxI
1pEWZczcWfR/0y5Ndb+H3m31Tv+jWZ+rkE6IXUuAqX+OaebBSnpi2PwhA6bv/nBj67UqSNHTojEm
OqDkC2bnjZvoknd/CU/NT8ZMgwUMPDTFJRpnUMHyLzrQh9qzVUCvakTe0FWIYQiCKOVl82j6W7ga
QF3GVpRNBevpAr4JcCZPwDPiNLJWMrEOmn0I+W0VUum0g71Z5IjfIMXoBAcSUoaTGQB/CHWXtLK4
9whe1D+3AWXSvXET3E+7pdP51xjncZVwJGYGf5la8DrI7gFGMvTpvMEksdDnR2ISVEBY+AXGsVgB
OapblBCNZAdO5i3tFGWm+GV1rbkNt3iBaav5TH0MYWlBVki/zexHp+/wVOOkn5rDLCflMM1WaUR1
YYzdZ2wvFo2iMyjHAwdK7KwWk+fsMx09Wv7CCqJymtheD8j3JCIqtVxLiRW7ISbtfk6iAUiBC9VW
RJqTXzOzzH0UwTR0Tj/IS8w4jVZRRmnHgbbA+vb8+rra2OD/X6k2R0bKf/NuTGQ9AE1DfYMpQIVm
ctb+fAi4pqff9NUwH74ts+suFPTiFA3+qi62KIMi0eforoaYH9Xc6iEh2I/xP5iEAfi7UQaErHoO
L+FNBSZ/vtOoPyVJtk0xq2y4Ksu76tmxEBjqoyyJ+Z5wJVRY6rJ8zqIpsd2iICSo4255dkWMl5BQ
JNh4+dYP8xgq0nH00pxf7sv9qehaYEvKiS2oERJi6jETIRXzBDDQ+QQj8JnslyA5R1ED4lfqL5pg
83+zzKcYdwzFo2jpzYJ6B1ThY8DOC44mpcHCDKSTKfcxDs66KS1sAWB78Bw2zgH8271nI6Po8GyL
Vf+WyH4o89xA8e8ldkiNx3kUAfSXu1sUQT0PjgjHcT539pqsHXQbeVT+7Igha/mS4YjMRI8YorbI
hULyXi+c/6b5S1KUdiMV3VXtjL/4369pcmnD4pm/c/P5GYe+IXlhufV/hE/zSjx6g6CXJNQEuyJC
AzEo1q3Y5YQiJhm/7YzYb+sjQWgXj+yXUeUvT/g4Hk8Vw2pYC3qnbcYNi34vkKahOhgS+eNUQk++
48yXetqTUB/7tNlkuF3NIJ7b83ysSJTN7aTVuu39xVlF5dTkFqfOlD07e/u4zaiftZDd/gBD/t17
cJbEHuEdW4PObl6RAsXTlFdJDdSD99DuV5uDsxpjBb2QEjur3zztWYRG0i1xkalseiAfKp2tOZdY
RkKVwTAqfjBDwfJKWAIfGhjo30QzOpKy/TNyP6+Btggzq+rPCS5mf5Q5TZYRgV48QR0wSPm5HTpM
bIB3EJhO9VG456o3DwifGKrFEpIk0tQEg3M7jGefsjeUkk58Md2yFkAUTp0hfWUGmszbfLS98C+u
E7zUO0jq+Mt8vCD9hacHb1/4qkBfND23e0RYueEUEBARRar9CnAFY7waEqSnB0bVcDBmLrOt65Oc
inlCTnJbYIM1SjKxjWwpfs/ufKdWEMSkb5/TfDsaEEIjlVmMURnflw+ShGv0Pc61ywCwq9xuWFE8
DhBCMZJgbjC3KOH7SAtz/ECg+fwbVXmsPDVkeN3TtBWjiyCJt6aIIACshKAZZc6FAPfVSD0Mp0Ks
rFGAhm8xBiO5c4c0XXch4xqBcrzUl66A9KKXakd2B23DUvp0PjrywkSD5cYlDaeAo5pzuF7eDs69
cqE+JdugCfZjl7onTnB3hRjBqFN6mbZPnfpkvHNvv9g+F2lML6dwptN/qS7rKyov/TXShgtJUfkO
b5VgoX6NY8UgvKgXmx1HjXVEPBDI3Prsh+Ly4tRriR5UOSuGs/8OUJl0siwkr1IkaR+Mid4H+nZF
NQpN7PFhHA+RERdtN2mQq0Lr6WHMy4fy5we8n6jWMM0ESd9Iw2aIr8oy3WEjZI3z5HzLlw6BUtZM
sXRi4FprGWDhYPI4Xc9pIo38lApw0xvcg+g8xJlXLsWtHw108K6qpzEedrCXi7+N1R8jdkcjJsa+
BSwf/8aLniAeVpcZyhxsxB9Ydvu7qp7nlzzXvYuMmcqOMyLgV57WPOvA73gYOGLSHOvxn6HidOa3
fItM2HCSSQaY1hKuQXXEqr1OSAfV/qcFdsvSBcn5KGhLPqwEMQtTScXdyPerpGxjgRCKtXzwgn3I
6BOrxbbnKNMvgWwxNZwg1uqaOTv38uJI0iReVq3wgHphnNJkYoLNtcVk5jMSy2z8clCNQxNyM0RO
/R8U9Y8z6yYN3pP2YjgVrGSFp75q9KgzsfD+uhphBrtY94VKT6QlCygEauXVvE7Lg8XOqS4TgWDG
bw7MpReF9rAFkPLtMo1mNICrwNCrG8NmEojJ+Rfat3d6YDr1+5XSOBtZDnquGqtcHVddnDJx1/5M
1g2QK0OMMrY1DX8pCrkxb03N1nuvORM8aZIlM4qRB/j3vXf8HQmLSgZrR4jBHWkvo6bk+wubL1vd
fah3amodnSbaHURMQ71t0UIZ88vOQ1H8/JN7CcUSNKVzYwZ5YBgR9QTWg+m0d9i48rvbJq4o+viU
WCrlApSYLvVcXCYaxNuifs3LUOGDG9rv/6bv5wdF05jSUkndaT/CtZQT/jJjEovldmOAFXjh0L7H
PgIeP281UrbJEwE55fdc1u41CrEttYgeap2LGHsmeddEAFxCGL/Octs/eoBia5ApdpLMoAr8rTqJ
7ee1hNBSly1Ha29SZ6Qo6bLD4Kot6D0B2wP6/mz/gW3Zf+3UU54lrBul9cgkyfAk9WQ3WGzjJiJL
5A4CUyV7h8UKnddCYVJYG1H7zSVQbg7yTwUuMDmdWAGdN5Lg3m+E8pTeaQH8eBno7vOoStkvHGXa
76yp4S1QdmCsHkZk/LgPoGwyeLvOancpI1B9fMrhGhPv+bWrhJlRV7/TEU6V+ybqrXYZPLWlJ29O
fLIZf1x5NRzyedYaK03KhNHmRaR8/vQWAoIv9W8nliblWWKHkV9zX5GvK/nAGyNKe8NKA/A3DhP+
awbfb4l0863X3XcNJFVyAG+hJVUJzcaclG52n9c6Dtq630EZSKkg0cwWbQjqU+9ZXIh94+atZ7Dq
H7VqStDY/Ir978VgfpMXxZ9WiGXwZfxve+OtJ1WsX4fqa9+Z/eQTpS0ibQ8MbLGJhfYqYE2jpJp2
aEFXyzd2xI1QKBU2F/su/gmQ4G5FSwhWpaUsHpCyOTcKcOOyjsiEAZ9xnkc1xhExoD/H79g+L8S+
o6PxD3af/Af/fvqt8LVeVOrWntYRaE47S1ffieKISw4ZttCfQ01ovQus6NIz4n6KWBrgYaQ0YfRb
ziIJvM0oH9stM2L/uZ/r6oCaheU9QC69pQAwmEMcYEiMxhEFnbK73ASPYIslgxIQl9DuP2MLYYn+
tO932vfyLdXmPux7BM3/avBfdMFbNTbLHQDmIcjgcgbVbyB+/k56pY73mh4ADfF4ZAuVrJ9fYfcC
ZMxFj/0nGUBiyOVcO824VZtlxUiUkGq/eQA4SfFuove5gBCx3PGoWHglvoAAsdQMJfEyZJK7i4bH
V2beDB5Jrl5f5oCcgehJ1H4Mo5rxqiYit1q+PkQ8of/9yMVtX5+W8TuLlIpCVE2QHVP/XOqtXNCA
XqwBxeNsKTSCMgglkmfJKBt/ksT8pDaWaMVw4iw8XOvICk3n+QRyWwro0H/4Z9lg5FHdGSBrR+hY
dgcx2OirT4cAfjTnOlyR24wUxFMoolYv192UJlnpEqA1gROTbtvSZDMjIq4NfCxW97+G6IUV02tq
P8t4PXQTIUvkV67lwP6U/QSIoSPB3/D8ZwpYC/W7QCYn36h8z97j/8vpHqLrC3RIREklj+URo2V8
PfbUd86aclNy2v0mpDf7d0ua/B/m5HGLn6EvemrmHOu1JjT6oIlvX6T9WGKR3Ki14NxGEbES+dpl
AcoEJRbOuV0+OTYzCX0wyhvou/0zDz1QqrANT4ud5XhUgOqAqswSPqPrAZ4JT/YfE6I4j3JLketO
sIDtv1+kBc+0TBLsYFOICJGdNY1ahBakE2/xw6v+Q8XmGz0d9WT8crX/o9a+WdexpGbFlOiFykIf
NkuDEZQijIlRr3W1Sqwg2PhWiy5nqI3w0xHalNd9Navy5SAlkd44HWlhQza/Gj7DltM+BPDCE67U
Wyspu7KmoSSdPt07kBGmDkKeZw7bvvnh70vkSh48uBfz3RknVcKUjXqFfsi3c77q1kX1rwzH8i7w
LrWzNDPT7TIta/3UU/nmQJTBysUbNUm1mP9s6TT2owtL5A75cxGxHIvymQrqHE3rTSVo9ceIUoiT
Fqj0JjGvtGifuiHF0xYiMvM/6WT2SQfBR7yiSs4RBR+dm9DOOu4NK3JUkVaeO9RupW5Yp6FIu2eU
G/8JLJWj5RK+vzRHp8BjabFlc5g1OmTqzd36XqRF7LyLGJuxQ4/UdAwmUw5SCxW/OqVg/aEfWRQW
qlkLyIw91QmzWSjSzliuMqW0r/6goAtjOXHU6OQR5F6oNf+NgBqXJzneEpFO+DV4dTw8xwrtx0Ez
5A4Qh8LKyLTkgT8XaLtdRIX8ALZMfgkLSZ61tnLshfPQNNZEmL61lcjnyr6NhwzmE7XUb4SFddW2
P97Ob2o3A06FD/QMWhDljXx2GYvO9jKJpThQla6P3KNnZj8tfCjZmB5gzXdXVzimM7fgnTT//imP
D+5E6eoNWXcOLyWV1tozEV9gGpQgzlQMKPTzzE8OJy8ftMcv9DJmuY0+jW9pq2JuhDRVIr2LzCD0
5E/DNYb55PCK7ql+cJmY+ICNAddgpJLloE5sK8U1ZQyPjgnY0TylZUb2JW+K+z6xId8KM4/nhuRi
S4rcNC8RgmkTSq6fp61hCrYUHdIp7Yhoq5HYv0k0443a12oUTDsh2Enz7M57XXhP5oHRa0dxWov8
q+npZKcPIa+lP0aU0a1fEw+Bdkxt2qbWNYjYlWoIhdWDBEd4yMFPFjS/WZVA7tbR5jKDwvrrt9GR
Fx/ZNO0QjCyGkT8Q7s3a1bgC7VYmGK1cO6JfufdUkDrVoMxzQgKkmmZCN3P6pRn+lyDR+DB61J9H
xHxJHvzwPldCTuoPQHjL9YrSgoC9jrhPzwJAHRgBhkBA5E6axHnkf4bky3tp3592aPOCFCgqySiO
hxYyYiKIQpl3/8tcHLh2JnuIt/dE+cJo1yWc1c3GjOov5UNCHoKhY8oegDQV4fp4ci3cozdQexvh
03HzHM5MqbbjCdZwYmpCSLkxy+RjD27tgVxS84ECGICDIqyzI0nZ+gGsI0sJQDh00q2rymilBGw2
/DEt056Q0txjZEnuafBeynJ+YCIyn0RebCkvUZg2IdC306Gwk9zGT1qXab6eBJQMKPPEzUgXuvPB
4KgUOT+RjTLHGGZxSWKWWhK1bOwNC6NcR1pzMOqi3gjTR5JdmKg//T9nGngjEi8XoFTdKr8MgStH
LyGs5xXZyHoVCe4Q008n36XD2Yy4w70n+mZhtEUhuZcg2iUazcmfvpyAjr9nMjkfxUDP81/2N4Iw
ObYPiuPeAhvFUfzeX82y5Cc+Rz1JwQ4PDi+InlP4e7WKxnoqJt6gIUg+lUMCa3YygdimcLD4WHZg
XJK/nbblBC44rLnOW2+SOuGCU2b94z0rqqu3xh5eTVQ9i9c4VP4gudGD+9DMV6qc1P+bjc0oZ1e5
ciOaNjg3k/k5E3DjatC6NcORWfkglFApt3sPkCZcgi3NKJqS+QysJrUXSYHq6aYIgd4KRYICEDfS
HqkOjcFDstdhSgygk8SuAiVYI8WEUHQ5PWILURpwiunjFC9JhawKAQfV1WebejwgyIF2Rv2vd2nB
Kgu6UJkdVGU8zJbAdgJuugyRUdnN77GvDlH8CIRe0T4TkZPUDkzoA8GqjLNrUh62CZosGqZGIuNn
CWLLlGCz2DmpcvrxQo/V2LM4RYbR+cAtnfvx4t+/qYyF3fl5paFsUmQOixxq9GyQ/2k+GzPu8Sk5
zK80W6CxlQ5WKZk7paZrVqqu9//OpTQBTWV7xGq6UrJIb2pw1VXWvgzYgZHanaXVTBJ92ZDbPlrN
ho/HtTK/3Xg/Rkk36NsuBZqcmo9Q8PGLWVrh0mOd3P0S62gAhmQuwKgd3Xc9b/O09mySob3b6F19
NjIp+CZztqyyaWtG0UhJT5WmOtw5KpqRtJd5SUhCCeffn0xKv5GgOdp93wq+tk+fp6ZQ9ly/kIdR
cmqoUrpdZZbdSyepvMfnb4VRTi9hVm+Hz96AsISvAEg5tOclgvIpQNPCeivP+eDxB7EENcPZYHWt
YRVGnwl8vSg+4ud7e+FA3xxgTqV06jYMf4ypB+jGSAILQp47Lu/jBxomf97VnThsD8blAcCoM1tf
Qp0QuHT4UHDpd8clBSCVwQlDAdWeiv0zfmq56G/JUGQOs3GlR2X3NY8z8KLBI2Cgvd6ZqmPjQ9lh
NVCINZLQT8KNoSsc/OAgM90TgZW0bLSbNJ9MOcO/uDiwiJpE9BQMfiRQYDpBd7CAwWB1kofrqAbW
dHP1OZJwULvQUb4VZxIJMkFUcCo0EfGo/OfnaiRJ5mOkO/z2HI7ByPSEercC7d0SxhWG4qrx5hLE
KSGxUiedPUlPOPnclWB1bwYM9KoWGX5BZ/jn73WQ2Fxtkp++yazriCmyvrEVLsVAmHNkVwYPUdJw
O1X60LYlrofzEO9m8XdY90MxRkqCyd9fB7KXIc2cgPL4Vr5Jd7i5AE+iwNbgT0PhCJgdAYPY2uPv
O/4RJbgVlF0ULIwdc9smpFnZwD5s4nAZTzo41Udr/Wd7xG8Crpb1HuGUnZ3iELZFttZQXaCHivXm
sXMX2gS9+o0vNc6CNFZggL8TlVuR7IczrXDGauv80jUGbcEG99O1JvhJdklrbcUez0TsajwE7th+
ICB2XWnqszrnG0XPnAzR5Duy/T3myjmhgrNPFoITD9b3Irw+IA8H+ZAi6pWsFiO9yC9xOSTdp42U
HWHqtV8D7xspIvxQu9MVmZ6wxSYG5hJW6iwxwi8X/eVORW6BE8m6oWoGjGq6CHxVO4kBDwxEkYSf
UWHHoC4oqoCqrZit8qcKOnaowgcEQ7Qb8RiDcgaA3kEXK5Wu11wtqfGClRkS/u+lBvetroOrUN4/
B2zOlFqw74orOrXU8AmoW+6F9sg4bPHYIt0dy0mQNiOGyD48u2SV1lINGXLR8IViOlJ4JNRo/Vl0
NAL3yE8zeOF1I5C1SAl+SSlWKHwiBAiwcD1TlWSJ01kC/pm20NkUOAuegsWMFCf/URcu87+3kMou
dVipYriNu4zVz3PeoSeFf8L8V9ukgqbdXlrIjt6aeDj7LVggq/xjzN/oEU9frroMvAceh4u1FfTm
sEszGzoF+EfYdygkp1UF0TpXEi7V848W2qvD2wVpSgF/kltLI0RrtiC2JpmGsHyFOBOVpHvsLlM3
UIW8qfZry0pYcdIODxqJ/xvCgxrj8lwBSW7ulo6WSCL9SIXkMe+ikfdb2XePhncMWixuFrPE7Hwm
0SRjy7bpj8tQqYO0KhjgviLZmJ2IDWyG5OaXtJn+gyA4O4o4x68zrSoGioLHLH2+3g9pjgKbbynS
R9cxSnk+4tPkp8ZuxGdNk8y5W7J+KaGkI6a5i63XuF8rsS2mJQ7KmgXkXgMCvlcr6/f6oJj4BRrx
Va7wJabHoewcrW0H0M/gcv7hX+h3qjkT8j/bVIqdGpIMnvAeNduM8Oznqhr3bktSWZ5f+bSnrK4s
jh6VHAV4KX0iHYZp7AmLR8ezf1gUbk9aPkPj/B6IE+9ErJgKB52IGt850qU+Ok22dcum3CBDnvue
AvgVDB3GLrtaseEWx+uqc2LJarn7IG/sBEshJv7iYsi42ioFL42X1mLSR0ZhzP7b2g3h7lX1mqAE
XUBGt63pRYX1YjNvcburRJAcbKRNez+BCjx79SxvgU+rRfEFye57w8p/Khmx0bUgfOwwLfJBvx2f
XAqPtbB2jhQlbeNU4OMSD0KSQB4KtxNldHEJswYq/MW7EnNXafZDCiowNt3v2xaSSmZIQrZFa/qz
cKJUe+5LElHf6CtZ+HGwT2KDmH34tTD0GL5hnJAqHRy3pxT19Ispw0XuEqOZZ3weddweYu9TlPc2
rIQHKeRriA/Svp4PVjV0lIyj8TWVHCCcEAvC5tFieiQtOnA5y4aqlxVXyqTS+ivpOtzlG1Q7IYOj
RJwDQzqtrs7xb6Zuot7M8s22MJRD5nKSAoINPJ0aUiEILzbpy540mtnCAhe/fg12IJKRd+Ld7HhZ
j9uUdXc1xDOsqg28pnyVTaqDlj43DzIe2efh5rb8G2P1EuIj3YY93DpOENsf8r44j+tBz2S1Df6+
b5tleEbQDJ/l9R6N8KA5p+tPM/dFRu979EDUFKH2uFIwgUNo6C+PmmkPJZ18vWS0t8/Lw2+Cxbw2
NZI/EfbmjlNkZ2KTIPmNG0NDqxCrvqGz/3CCwHS16AFMIQpUoSZc33uQCsm1hEe1QouDURXL8XZm
ei5w+Arf2tH0pj4UPlyGOtoHVh0nPC+HmZ0lRtFjW2bgohqne+Qt05fBjIwfQiOq97/xGqDVcutp
UgpFCgtJ8tc3mq0oCq0W+jXw/OtWWlBXqW987nzQ5lyxAcfd1fPivlwVuaCbMog9wEB0ep65/gqy
C6pTSVg1WHLG0mMG7JYESQQYkLJMYOjwUv4mdiIQ5h4sKiJDuIbLxUWjO4yzhVFUDiq6mlVMQH8S
7qChczZyV1KQOdpG9mfBifnWkrbq3BTGc7VyR0vLfsdp6BCyTKiKWcLZ+lE3nR5ttDfvCg8Cgy/G
qNtuJVZRABWtgiukYx5NXXDy1rhfs+xVsj1rOMo0hplBaT96SBAEps0QEABn8X51FQXY+1zkKgPr
FxaSym6B3gOEb5tqSs9EmNiYv/fLXqSS37LzOnMD9/S2yj6hQCVCbDFFGmB9UofKWmMEf4gczDnc
DaaTHBFylcsuRJb+wlpEzrRX6I2a0Bi9a7ZhQMGcBWH7yXVMfPt6NlVImbtz0uuoh/wIuhwEz55e
8l/YkGRppXHRJ1WoNsoX537v1BFku8nANdceoalatT2FGAH2VjtxpvgDF5Tq845N/0DnSHi3AqOU
PFLi43pF8AeyxNHhI5jFjToK5Li1919jBQr1bFrErhbYitrEFbtv0HefouN1v1uwqavU/yKsxMmX
57IB0C8JuzkXqF+MQOXzBUBnyomxPqTnW1VcdIv7wOq6SXKtslYDjY/tPZV6c3qqM0ON2BUFs0MI
qBsYm+c4tw2ss2nPyYkB+a1dXGrYpxz7V5+j0OOsx6/NVRhFq3zPwS6hJ2jWNCJU7lbw7PIL/xHH
7mY6vtv7b8iH97XMzgehQPyH+vr8ktygESiX/4y8E+wy7LM8Vb+ubOD/tX4D9MROY8sRR2eDYbj4
w/dNnvUImEuAijy1RcWrmzeX0l0yvT7dea0QNyiKu/2e6fj/5uW8MXxV/wvyMZ3MkgoIE2R9SuL8
T7vDV0YGfyke3eW0Igr/7EW2WfWG0D4t8El30ccGxLqZdFds2pkq8UNiypErbQXhphgMNB0cub4D
xcfRj0M3ItIDIQ8xzjb9CwP+d9XsDcTDI7NKTk5m5kE+nQdWmWwEhEZsruZ0ciFlihGR/qHnC0nP
Lv/gXQ+diIegU6XUjibuTmwuMMvfioVU5dD6tfa7XI1sZUECY3pORezXGviMVZ/4MUQx346d5UXJ
UmVlZmaBRWNH96NxlaP/wx3PAq3rIIN39FGv8FLbOMzthtNmaVMjAxn0QQOJ3Wd180ZKYU2lNN3o
hZM9MVA86AFLWzGU8ZhPQBc+eXQW+pXwAy0m6uICLqmiCx5SbalEkUpeN9Z5ExGD9L7r68fITW9X
i8gVdDriPIiCG1owwKrAdAIPJZnDbz2GwjUi2CCEe+/Mp+ytTQ5er2TAh8dXtvSBOzRy/5TTCgwN
OEPw0VxbdSOATttI3LWYlz1WuMl4BrVq9EMSVagb0K8ZZZLcfFyI200r1P8mMaNiDKcHbaXmRRKK
/B8RLIXsJatd6YGIhN+/q3yUYguWxCLHdHCCUK25jzhfPlI1Jg+YhPScQlHrg8sChGLuvsDJp+Ur
HdPOSesTvqBXEJh/levxoOX+wPQwXFM36o3cowdEAx4zHgGLMMSzW8v5yFUGP/imfdcC4sEpefam
SZjFQXiZYyS5NdQw92iD4sCAmfLJUpSefxJrv+b+c/A76UHS697dFMcDwkN7e4k+5j/VrVF8UB8p
VCv21pBbncEYDsmlOUkbAEQhT9vE4WBM6V8/hxHibRaXU0YDDbdAq2u6mcxbFCjcJvRyDv2GvboY
k611wI9Sp7ZGig6+GwEwWlT/dWi9Nu8JnPYcS68XkVVw+shqSUlOQRckPOeNbIR6XfAAUyf/hRz2
tsS7Vs+HefmqLdN8bM1Ot7Gb/TeUUy4m9smJ7KmbwmIYZ8DDutJoOSIhm89VqSrEDIgRZKdEP2Sl
jw9Uqv8nq0aT0V/fV1xy3EDttTeYhF1KhxqAzPive6rPYYo2t0P9Y9010kcvNYYjhkI5AsBm7+qc
fJqXk9gYknXHR0jiDI2xQLM6+eAOXL6G0cvOdUv80sjs377hCA6/YoRn0WlFSKW7pySHXV16Ohf0
kJzDc1+/J8BJAWXxPd5nFubmjNy+AMtdTLppVngSeHUhwx/4yB0gY5ROm4v1U8tqBhC1sUhzAZCk
TRiWo9qpLoBZ4felLepXz07QJIboRxi/9OE5NtpsFXjmwXNYdRLZVBIAZlpztxrEzvvOkK6TvF97
6kSklAuimy4vfA+z3EnkJqjLtDZrI+tu6qg2u96sDOSdwo4eqSbEVygEwoQoqLne4oC77Z9XWgzF
GTTOs+O2xr0dRMFC+Cg3mGELAb6lnNVSXckIYbQD2G8LIGGE0ilC/6NJy4tqlj6IAncRPXqQtgGm
5hM74kihKLb69MX0Myt4yxhoJVseDR7pEdbmRUko5wUyqhx8AM+cwMdysKj3Il+YBfTBHJebubxy
pxqcXAPYvJLh36csrqvFYroX0Yvbxv/P2Z1AZJS1FLrpEVOmSyRm1j/cf4+uCpSktV4jJ5TpLXMj
PNyCGJ9ULVtUAA191B0u7aeGTnF1ZYhtA2VVuTKd8bghPKKyXX5oxORWbHA4MQl4Jga/OhXYfcIO
MGZF3Vhb6QyXJWcooUYsr3Hq595VQwBWLccHwRxAbXCyf7gJieyPRcPN0yIbx8vc4SpbDbKScIfq
g1X+3Qe7IYJXQZRJIOSvToJzERg2UE6Im1DWhhDBX7Z+v1c5zTCUXMLmWuWNH+JxhTaryTfxuJ1o
UvWly/4dGbeCprNhGldyYy85LuVQdDkWYgDW28pZi2zHUJxKkJLtk+MvvaNbJ2S/J9zNfR0C/iYV
enfgIInVMVhpAi/PlfZDpuWGHzVPUple4qqxVThcoVfDq0ng806xRzOg0TUDfV7gU/6z3sD/eE+d
yZLyIjvfTGIXWaFr/7qgDq7xw7+aXUAeu1G02KLhnDjpkT/mMhNYPFjCKOVfBdIxdgThuwcGBdkT
gvgf5dgzPqBpcfU969/7MVHaoO3Db3yRcrAMLj12sdxDr/ZCle9WgWz3RRJ14sb82vczzSvwNcEr
IcFCzQc3F+qb+YzjlirTyATgBC4vV2su92zc00BE71hcuLEsweJTp9xBEv/sdOnEbGxDoJmVHCB9
tK6QrOaFE9c5tQB+Kncgudr7DA4oEcnpxbrh3tU3xjQcvmsUz7HOREDXCiTved/oaMUTj8g68s85
HQFOG2TzsJyEPU7yEay6WPJltVmuTufbJI+0TE6bhOit2EnSNtjyhryjtXHqlg6GgLWDvat1tlKZ
iu1sLC6JnOT3JyR9lmgz221i0zP1VF9lMuLDMkRw51W96pkOHRBEX2zvFsBinoNDY/OcXNOHFLD3
3dNsJTjlYUoVeIhigDbWEsWvIGOhhjItM1Z0w0nuagi4kpx7rnPVyEdIZ3qqy+/fm9BCMfl3uz4n
hu/HLmOMsYDNCBaqGi5WV45qmNon+NCb5ahTtnWc7JMF//LHOOJD2Oma1N5XApI0Djz2EDy385yw
HSYFE4i6Bp/pPDYQiJi2qFigXL8ZvvUkmLLwoLftblWRAyoh0ljikAKAdzt3fmV8ZzgV6uXRPDym
5VjRUAuah3nJG+Hg8WMiWmxiwG/eTQ7UnjlJCPmAKD+VxIucCl8VIMLUjzUYjIt8NBrcnFQmx4zd
hGabMjpCSB3UxpbB2FwDaVooGecUEkVqxsL9PX9ynMw9hZ1EmyW/TTa3SvFoeCOzmEdUJBal3xwn
yj90iA54CFOmYP5bi8EfQ4SZspFU5SBKZlDLYpfEX/hkY4VF7fYwOLlaWMpxbOB5Y0e24NJfxGc4
tik9reybSnWjYVXFxkhhXxS/dQ4RcPkiBt3sCkrPWehv5JEGBhhrbetqODpvnSmxBsltwZ1FEMU2
ySQ/i8xhfTJ69zM4OY06eDpX8oHRAogKRsHVooAxjQ8bODLT4bhuTTmlVJ00QakMR0chWzvD054U
STXiuaCQtUPjqBFFXPIqCirYlEDtmUMbm5t8MgUboJ5ar66v0xG1e1G8zKA6IqU+kJTbxklnG0vU
6wKPLevTDxgVV0xdo2YIjeSFq3zmvtp8mmBOJmA+W2KRAtO8GX64ZbCLfgS7LZTl/94e9TzvB1Hg
0m5VvU/xoc2lEMN3y4n5FNEzrxN8WipGycEfS4RL+5eUnkmjxQH6BNgNQL2riHQ7FkKIUanYV3XF
a9UlwZztvoW5wJEF7LOnHtVvgdXNXEJbxvmoqVdl1CP9dF9OveIuJ0voMgjtamYfqsE7k7jMd0oc
O/n1Js69Q7MedI8zsOebMbcnDI8ulGhaDXz/srOI1x8/iWYD+mAMngtyQMvUjgcb/gEBWm7yzZSl
edzq/13wdXV0bjCK3EfO69prKmiFDLYaCsKUSw0GjYA8xuLKhy14WU8EAq2EPBMK6BjCE0zEnqlA
bW3XH/SgpOJ44BBwmAdacYJFOdQK5cLsgVeIjIUV3/GfoGs7By7fmHuo4tR98n+jDrg4kM7PuLKE
zIBlWJocOeYERVQmxs4ls4MdJVZBcsltTr7RK2G4zju+ksNEKKeTz4+akpfenA83qY9fwFQsVuAP
362m9DrTL30NqrzObnX8wrwXihfkFntA/nZxPODG8vegNGc8IuEsoeR1lTF8wnotKdcgHklSWWNe
zzUGpCuGYWZ64mBnIdWmLvNECP5wod+RKuf9i3gQ7jv7DxMlfazpQ7pYH3xDzhfUZE1j2wHmy2/G
usL85Xh7Zf6Zy7P9DRDaIzWrlPQtsNLhv6+OCVlNEhUW1V5AAjxTmbU3YyWUMOMFVmlSPhPnjKjm
OlvuJ86P+RCXB55paJGbGaUx0cWj1Rsdpyn0y00MpPYKA/MayIBWijZMiy+Vlzyu/9nlKrikEyc9
IpG2tCWnBDSnJ5XeueEXe2V5SSOJykQHuVrlvvMMIFdbKUOEuD303nzYn8q3TcHbUa0UVK8eMZPb
siJNTjI/ipdPt9OayAzJ9DRTM35WJ84+d8Zr14XaFmiF4C65aI5YHPmhFc1vnWzEvfdLgPzyN+Bs
krkGa2FkaSzS+ZmvbsdvA9kqbYv/fbbnLOXfP9wsG3KsZOgVrwNoAGqlfgizw4CiOi+CBRsnq+eb
TvFHj9Uv8klikDKeWH3QyiVv+3By4bnOka5+qfjBkCphVoogkNHbsh16XAVDQAETmdlTqSYdNq4a
oN/JjHms3Yr1Y5eF7415wr3dxodhSJfKqN0UW/N/TzXVcYPhldzTaI3Ln/PxBgUw8uuiJ1F4VPMO
g79if4SO4zh9YnbV+29FwqOjEBlWdmfqWYdgfAZmjvkJSe+MdFHHMRBotWunkzGdtgmFmhYbS+Vv
EYx8+xpiPuwBvhCcSFw2cDQP+A3TogFP5Dq/mMVZjgchcdMpPKiYk9zlhbQ+AzxNvVhzCgQgvJxb
h6K5H0wOMVHiibiie6mOZ48wACu77kM717kDbHkxkxAvwYniEs10izBlYsXIyg1gRsBtmcZGbwvq
bWENeDi1s1CvehwXeXZ4FqqU8MZTHXbr0SrD61LhjYjO8U+mEgnAucvpuYUmGgI3MLu6e1Y4wB2g
A1rdpbfc8bLlugL5Ipf3K7941dgK5HcnhNDkttkTl4JK8//XsQuLMFxLYJs8mmAg78It7FTEl/Qf
E2jRR6v0vqxXI7h1qffbFSWOYowrlVPFmmX39Qxw4Vfwm8lLhjqqkam0sY1kFGQISKt9/o0A6NOi
SNO/UiAlaNIUdHivjbbzeXR5/rA0fu0/P5jjr1rYERHbTTR99ZjCftaxQLWvgkT+DO3eazU9Bhb9
+cM6H83c6NbmoUkxjSbS61Z8cBVje6PP2dSt5u5Xqxdaj6Nid9Og30UdXERMI9iGKGpO5BEEFvBd
0hHftTd3KvRQEf0bJOx0vAKEt+GdsepZlTzt/2FHJ2UwbDkDCrKsZlI1B+g+3Xl5CXWgi9CJFd/S
U65mbmx3xr+BlIllO+ARTyGNvPr4wH+sBLPN9+AUhKSHXFQMvKgP0mzTL+5MULszPBw6IePqviyj
51Sf7wCg4YvNhlRBxWzjMdEEZmwzhbJPFZ8AD2+AWsdKFgQqgg3OhrYFqpQPLJ3fygihl0OFXA11
JrtpdJYnsZ13HIgiieDjo6pDFBUkgexVgA4287WfwDD6G0OSwbq2HZPsHFKrbOhfSHzUmSi8u8f2
Ska40QCxPXrdnu/YpR7RC0DzznDJNLuScheLC+zl+ylCCw5flryI8WWPANYuRgR3NsTLPT+YJdHu
7DGdedHMJHyrxFWqL311zTX87E01RZ3MGoiOxqnOktWkbGN+CNfIPUbbXYR59LDAUkwzpbYwnw/e
ao/lPI+iNYJz+aPw0CrB9LFdPrcFu/uqPtNhsedCKDDoRcndNbnxL4YWlE8CW4HmHq1WmVccVZmN
JJwtNyKsgmcxp7OhzhrT9QwMjctVGtEEH/es/Zo4LA3EKatKGoqay1HupeW7XHluyM8ypfNf5VAZ
LUVgmiveH2LpKUU7PvEQ548Qvjf6lkJ5+wVeEF16FsfYptF4oUzLgKUt4v2utvRRnoekxg0Li6W9
LnsTM8xrLAeWVgpfqA1wzf3+fI4wzj4p92VIRHJW9m/1S9u+4Wb09tnXumLMhMB8sp31si8T85nT
nfYMF/stl+niHHA1YOBgoQ259cz0KwtmvbKXLjPFc9Zq6hnXXhI7F3ieq8oCS0aD6GWjDwvjMurk
W57mBWmBasHp7Cj6VDtE/KkO8Ga5XxJHQrlAx8bB6Y5PM1hWF3Kid6KBuGTsPXd81Nx613cpQTU2
JCmIdFKwqYV/3QWe0r+kN03gxXhE1oo+m82eT45ZvD+7nO9AlXDd2JOWLsTj468TgPaTlPf0eovo
aehA1tQTqDzVSqA3QuR1wUKrthj8/i9Wz58ghu2JGol9CS8zV+K2hVDNebexg+sUEHPVellYJA6/
j10SlNcKChTbeC0iHavjkDUIjvKrG2SwD3V3ajuWDWrc8j2rCfX6d8onyfAAQUK1oxDODp92uUl3
sn+qvS5nUPUW+Qtud5mjkes+bnLB+0lb3oRP+og8iqDyspceXp0OtO+Ac0RNXbsj78BSbrzUVuos
z6bV5sOWLMjta50SD5negeAM90hGftKat3yUp4b6HCcoG/+6Vprmrvxv4GggZY5HjLf+uKBVtiPV
s0cV3hqA5O4zTn4wHGzhog5Sjd5lr220ra32gakwNrG87oPray3qU67XEh4rzZoEDSIlLj8h2kTS
5Pg5BuF/RdzfA6meZvpe6+NEtaeVHyjb2K0ohbuHU/RiP5CCy6bTHkcllHe0n+LMSUjBBlFzYTFj
ee1kNY5n2Q/+4EPy+Nsj6rvMAkSkSFdga8g3MVazQqmhbbHxhbEgTZUCjhTtYW9ntX/oVx9jCgeN
lp/xtRXHXj6SHvvTSeCwDDfXPwRbmnmoZ071hiUP13c1/kpbu5S41uCD7ZTjVoWN7nXoiOAHkv5q
pyI7tNhPoDbjeNNO2NMqwR5XXreb4RWGWrbvYdKb3/MD2XbMGx7hHqSwZ5g6JAeRhA6VuBjjEMCT
tL6roPPrvlw/RobLzpVhEKIwx/J9Bxm2bXzd/1w1HtyBwnbDEAy1oPD9ev761aMQS7zzcGsBYvQx
0MEp6lbVP+iCvrOr+50VXNWb4jJYVsMCyZpVQTqW3I09rHf7179I1HhtwOkfGSUp5C+reV+81CG4
Ngdp8ydOJ10ZtiaN0Jqi13GDNxVK6bbKYT1PrtH8eln8Y+f9wt81mWQzbG2OhlMiEnht+pK5LJw4
YoARDi+uIA5iMVj0HSsWdvsJW3tV7MtQorh7gaT8piiQ9+8c66PqsvHdCFmGuFD71rpmFEIbrlMH
o9+zgjvyX3t5hwR7H+eqMjUqJri8xOZCtIRepHPsCDvNeOkDfKuNeZoMka659GKiiAn1BYme0UPc
uBODKSpw1Bq2AT0EGUrtYHQzmidO5n0ZytUH9ccYg1oBGZ15/9ca1rlc/jAqcgEB962BspCQysC+
FnaArUTRVA1dn8/ootHk9tg+XJ4NeAV27F8NvJywXEEf1G3qB5uvT/MszhRFtHmBlkS1k1Ue0M12
wQ2nhIeEdUoEaU4amb6EtsuI5WseIzH2z+8TBk4ws1RVfOx/YcBfTJeeLjdWcYI3EP+OrmXjUZWY
/sEsOb2HlmOztXeGv2TCFctp6odUofntabKAiiofLVVN6BGbWkIyUE9BjiS9w8ML8KcQ8QmYFSRu
QFGOCbBvOkm0fPp+I1RRm1soaNMFhkFsYNjWcmZ0Z8XDW+7r09VZBIOXhTbfblIzzuHLuzsKH2Uk
43WyFbhtmufXkeR+4D2MwcoNJFPeR0KkDecVI+3JqKtpfkcOQEkrL77xiIemjKPlZOfglQ3sHxVy
dJM6mObLGtIh+K8RVn+HEqSkhNfCQulYHi0rjthzF2dNDqQbX2d1Zu2P6BkVEWDSFuWZSQuZKv0x
SukU+5+sq89B9qIZxDylJrWinY8Do1y2Q5JupwrFIwa+eH8QJWTJVEej8YsitSwFLoqpWrQjMrK8
faD0l762Ok7nYOXW8v7le5whExOD2RtHD2L0IjB1T0iXCW+DE2mJ7MzW1qZP0g9PpMJZRtcZX+kz
eSTV+jaqlA3YNLQSfggoX/WJ3roofiAqJ+BsZ2EjDDPMADQfxpimPDE7HxyoXFr7dDegFv0fbhMj
TjyG8UWyXaozAsz8wNLXjKFCDofyKJm06bHOgADEkFogTEb2PcjBeE74TkLuuj5Y7DHzmAg2MbwF
wWWrn7sCKzYhB38gQaoasDo85kG3rFIxCSNoEksBeemx8wUcaxe6i3t/B6myjcplL+OccYpphv3p
bT8TeajQPvUP6TJIKPSHyMdNmf5ji91YNFW+VV0oBt9DTP3ry/vfxjMWfchhaqW0lPRwEEnDgM+i
Vj/tKjZNzwEJz1g70rJ7VEDJU9jx28cXphO5Dsg1432B8lZCsTtnEiiRhsFEcfKqeCuTQm9Ftvxi
Oz5TtwV+QPUcf7uzutN2sT9UuFrj0zSGARQcIeanCXyTdRjIC7D0bINFBkBgNK5TA0XJNqoAdE9j
3iHnD8QPNGvrFqkY49CYDtWY1QBbzM0UVMc9afhcCT+AKZoVLA5+kJHGlqttjkE4TM4yiuDh04It
zmFYngx/DzHCyLCbuI4J+Ntf0YpSh1BU4ewbI60AU6/JytT6sV6A7Yp/VuUCKnzV4ztQkZPVbGo7
HnLvDYOtdmzYaqefrcFOyIUY78iY2lQbXS+T2o7yX1Kzzj+4eUpbbIfumZudJJ7F+Wvo31s9/oLO
0JTg3S/09u36HHD11uuHZhxrl9LdfZo2i5a+GDhtTU6Mjit1rrta1QC/IYkRC8jo3ZvQ/PJPv9jJ
8/G3y7zz1bats3uDZ8opBHfkL6tAIHCNGMDwyIQSRzfF/REIZVyQqM7iV9SgShJY7ZKFClNY2k7T
LEDQ1aZyDR3z8nnbbOdjMBHlBc1bGUN4B0auJz+7O3U09gbM5IRppQDt269KKvLD1gWGgoYMHt2w
csNeTtAw+Ez20m25rxtuv4894LOk4HzsIVcwi4fF8p3PtH+5x+zNVHifFJr6QmSLQPCg/BgKMctR
I9Cjxlk+lm8VeGDQFC2kCSgSCe21xjMHC6IW435ut1PBHrTP0OdslExBAfoH+b5Jyxbnn61zRF3W
F4Jnjmg3TgCEVgI9gbMVDlT6Hoecwy8Knxc2JECAwFCA6t7d4VLikMyA5rKlXFa/vQxpXoxTPCuf
mWzxDDFIn0PnuJCvaZjvholaW0L3xQ2L2IWHob/y4dELbG0LVBJbe8DdA4RZUkfxxl+AlMyRYoDs
7qp5vCjOYhS3/M/JnUuRXuUyOa/8BOnGUBvjDMj1dRtf4EB91wxxUlqz4kPCzhdc9NIOFRf0qccq
C0PD03MNo6ltreBIJLujsaoPHlJV8pb7MLKKuhHMTnY+OVQvXbc6kEcLybbFYj87bCCrgUKVHNW2
Iemp5v7rPfHgJbOZvdDv5WeLyNnDnA3HkQt3qfAaMyO1zhTgD0DATqHjmth3GmHZs6c4B4zl+RQZ
JuIseLTT+FGbJJiXKwnyf6tI5eeEq03dims+ttwgejWHzso4LtED0PQMZ9OwK6Bl/f0O0Hf2T02l
FPZKMxd/a4gGHJ0KLpCj3nR/egid/Z6LA9rr31OsE7F8PshO5aQ+degwrmAqUERV7sVnxqJmw0GC
aMi2cO8EZg4mUKvXCAVmz2yZc4XPjqIs/CjDtRaW45fxhcEHF7Ofe2QlQFMo0n9jWRwMfxorw0WO
uQTp/QruA9CmyCrFc3iT6pSY7ijeZqgIu+EqYR94F22LH2IzAUBAP1ByBkiVWbb8fpaLIJmmForZ
NpSFQieX6yHP/0OxQRdOJXa9tIzpvMYLyK+SvA5+e5T1FAiRfvio1j4luuDXzkgL+/0JsBYkFTX4
5N+G9y2ZJNi+zR4OOxr8vZLyv9UhryPORFLfGGfN+U84H0Cf27Aop6mCYbk3j3bawcn5i/sn+83/
+RMvufK6uoVun1+oCyDtOcOg/yGCbNX1bfxURJ9HLwBn5CV73UwkGDqSFz4udgyuZCl740C0exwb
JHzxHQO1vJGALulajgkfwbR+Ma43n+sC+zPO03AK/dRebYgeMsKXqVhuQr9IO0/JsPIXo6gtJx5f
VXSzI2yB9GbBz3TGS4jn0OCwltobJ03+E4XrDksehY8k4/PjZzvpjEa/Ivfd2Ddjuljjx6UpcIG2
tBmwaXK9xLUL0TIQZIXAgBxbsL1+kUUBBcPlWpkTJURwPF/7/0zNN1eKT5GC2zzetrkArOjxvIx2
F4difeD/7OdYPPjDiAfOYJ9+hhHjcGh6NTtnwj7aUsbeRf/o/lv8jHidLD5cm7LLjsctonB0YpY8
agF7HBdj5gnoZDBQ5HyYmJ9yjY9xVTLTmljOV/GdIa+3sJ4hpVJ7V+rCKQxjCl3o+HkzUV0ACAZf
7dNGPvKXLC7a07yUlCUmcQ8u2fHHcDU/6sMhHOnL/wpEAI3CWTvHrZ7XpwdiUdIlo6W7grMM4OgX
LOS5ML22bwN/iTcs3kEncDLjDnZQIQh/HAxMcIaeRAm3aqwiQlpt4lo9A6Ja1Sb7oVuTzIiDlBa8
DWpqHNmE8kZtO+rMqj4QD+LYYPjlpRiR692WjFrKygdq7IdSHh3Y0mKgCwU99P9x4l+D9a60hcQc
7URmdWIJYW7eKAPCzw788BnA9SEAWZnlCXegHXZ+kFoolgtCEt19XkZTLlJi3rvhE6HJLfeMBX5J
+XFtyfkE5sR28/4cTlaqQVvgxOVzQJqMe8BLDwgy3BUDtKygAPgNNg1v8+vAkUQhQd6pIjT1CWmG
9byZ2nZx/7oAJEIU+g93ikXOEvIdMb2djewgXRmErMfZNJgLTHqO9sYRcpohfH9fXveW9ZXq4uEj
oGCIwBVg3AVfGt/VUqdSyaqJ9q892WVUWIOd61tvIymOrNpnevvjyqQTJHaLlIC0Ko1masrTmAA+
NLflsEPA0iTfZ4MLZLr0lRzyKmsTdy3oIWin5AMrchiCSo1cwQ+5FyS5Vm2IFtFfgG6quyrHEPeM
0Z8dZquktCzIEhuxQrBek1ykvfySDgfHMP7lN6qCZRMkULSCB6YfTxJNp8qh2tpy2pC1c3Na+pTA
mPKqq/nDbY6QQV2QohIu1at7IgJ8tcVBTjiPghKW8aJcRn5hoVHy5Ggmj2f415nye/z0376UtnFc
n+i5CsS6Kkk86bugxMmmVM6rfPzZ/4NUOeE6j2lWpmlhzZhIqlzNbMmKJVCccpG/YJWynaeoxi3I
GAcuz/wppMjKeTrRjeg4iXyYJiBJ1yLjovIOeGvRInp+d5rv6VNwD6k3YPcVVdQQEF0Jpz5YCyZF
osubvrIN5Ff2PX/THhj/Oqe60VkkgfZ3aNXvyLi/sfN+h70w7t5tBibGo6aEZSLJ8LSyV88+nPHQ
gjTyKCzq19tscmjhJfJwgGB0fKhJteQdpcG8xmZmExULZ5FrI+8oblhSFMRQ+aRfPCK6sYMi9Emt
EKtVHT4j8BMWtVwlaGTVpy6CGJu+9L2kr1NNWcIEbTkZKKH0wHHIiR1bsCHICEehyRRrdr6d4L8Q
KZkZrkezXde1ZlUayjOqBzd6vLOTdoA7nRw1/VkdXVLr3pfVzAQ+8vrnPTAehlha9jflTKaFsJ0Y
CCXG/82ocBPDoHuK03LqoOP71L/yqlh6V0JFON6k/lmaHAPmzembPsSaObu9rMz/i1Rs0CUNAxwe
n7s7zlnAvLDJuYQ5RbLYoaRs9qfwN5JQ96JLaT7HnH6FNp2wH3d6hfX5U5GdvGgkHiCRDCiRwUJA
gTpA7P+rFiNQUYrbgAsi26fptmtv5LBpg8NuhO/grfKwb0AQ8QuJtyKw7fN7PO8bKgmVRqZgCrq9
LxAwQMJDDl+zV43CR9DigPcaeirNWTnslU0N86Ubq9BgioB+zOvIy8aHDcVmCm6FjxTMTHpryW7e
rmsJJz6xwL/WAb3tCLApEaxHJGTQprq3gyR7kHrwpZaANFeOnCZeUIi9V141aTa1fFKgdYsN+xkv
0QS0aC1sV5EMsxRm7jhriy8o6dnDNamP+avyuFWYfO07rPQqs4YsMJaJC+R+sJ3C4PAlwMopeGjx
9MBAGcSJpHG6TwepMIL56sidBjy8FiCjHTN/OvjPsJRV8Yx94glIurcFkAUOJH+yATnuLx6rbw9d
Esbqf5EWfK7/EMCxGV65bQv099PodFy78GaGpPObNT60Va1B4xqhvtzqG+gYpWTNULFdYESQBl3T
vm0x72ONO1rzb2Ql41XFxPIXBpY/kw0CRqgG/LvYAS9h1ywp8EJVhbzJEgM8901NhX9QqRbxlUYE
GX1r2CTj58Eo3jlbNheVIbqOdz4jfK0FmhgolW75UxWFvas8gykHv+J57kNUcuKIwGIdUGeQyAPj
M0s2V4xChnFmWLMojtDqR5lUDoK3pMHK0MkrQCwLZ5m8be1uHy7YQU9LY69s8IjBVROFK28kIkuM
V6s0ONQyPPG9HklNmCf3r91zywZc2JrwOWtr72blGqJv7/r3KO7YbsaazxpS6rTNwfS9O1XuNLo4
yg5YgwQMOMn/uLMLh/kPakrZJ8OE0OEmWnWKdhg52JceoJdEKQdVWI+C4MFXoVOyIwW3FNQaeYtx
jFOI6rHtEDUeKGlQg7vNg1tXoET1dt/8KOnrj665K4LHqKmdILcTYKVlSE8chDHI1eRW5TIgEDWg
Vt75NXT5bU0akQxMJ/0DNzSl7nlZz4T6HPCK2NMJ7CAAgDLRGo9yy6ZYB4Mfuay8prKhaQi+K9lS
81fAA1FgYSTXMrLW3Yy1GpgpiFGUBgkAPW+R81PDxhz98glfMwJZIFaxZZG3jIpAeqWKpaJz1rSY
/1BMrLINVnRa2wSrswKP2q3A5sZJicL8+EKyUWTjbiX3o6ZEfGJNSxBK2DeftlauTalV80mg5LfX
eQOvSxvR+ce77oNYN1cnZYku99STlQmo6ydvmTxkyUlkvg/d/QmmjZidFGRh2EThn8JA4HigV5Fi
cBP7709e1kjN75Mq1T4KW+/hFYM1/w4B7Ngd3PMzvVVDCtsau4J4dnjFwTDhMsqjKlkE37xb+pF/
6NOnyypSsOn/vuqTeUfiJktDPSSL8zoid7UrxV4pa7HoIJKNM6TDynzeoYDqugv/q99GECp5wHKg
R0/BQ4SQjP8N5qj1BvBh+48eLrFAJbownYf7pUq8LuRhwK9iINrCuyFuxOxaWQgQRyHQzEBkIJAD
MH7uz923WHUQYFKW9iZ7UfRvQCjhx7HvnV+2tNOKQok9KyW5bXlUT58JH3GdhQg99Zu82eiZD5na
PIVvBnmHTrinlR5fFwgVi3gTwvi1LYAXN1zxBTyqeiytQVuna+JRVi8F0IjADI2huPpkfEKlEbvI
/3+wkbycnBmxxZopj0ucqDh5klKsEpaIkqsaP3mfWwWtk/nLB3aFz9fo6eetCryuwVAsajLOILHs
/pa4+V1MGtEW47mxoBvLS7R59JWtnakKMJV9A5zSWkGrXmh+5VTcv8z94ZYVoZy7FuDoUQSHEyDa
9+kZ3b5WyeUiabd6DQR8MkkWdo09MJgTty38VlloR7o1a2J3K0lyZcP7EBrNjF//hH1ClwpT+Bq4
cIQK+5NXk8ddgA2ns6GiPoSqZZR5WBZ3BFgM45od0HrA53IiDFCLdLJA6Aed6s0/PkgMoP336DcX
q2l8XlkOj9/bSv2d6rP0yvkvKMKv3c2lUCyJcNc0RO1mIZKJeFb3f7G9fcVyPVDu0eBkEAGyteDv
Q/yKcq5NM2vpVU7hmqL01YAXu5ftpkgpqaSiLLRAGycvPtAIWGcX1zQYE9QFtPy9cA3h6XMLWL3+
8bS2luaBXjc4pmJD0e/JJ+qRJIz0qlTpYWb4uqzkhBhBYTfcEBfiv5gTHy7NHFcwGyLADzQfRrpP
hlM+f41lXhfVma9O4jvv2UVfWJg6hH/jMvIT1ZTdLtPzzQFM9aX7hyuzn4mcQKkLCSXG4NO4lfxV
fBoQ5luLrwdHv0/VBjZGf0Ehk52A07uf4aHZYNQJ25ll8j5oYcjcanowTbV3REuQ9ORrHelSlWBc
dODTiV/x0mqr+p0QdWYUSIaAFd/9SOt3wQmW2i5mCwr6ZNghCygVpecXFhSmhiKR/MuXVaQNuHvm
9eGMxlJp+tYxvQcQZ2Ek3tDjkemZBXJBbfYEAyT4uTenBDj9ES4Gxwy4WP9R0V0Ud8M+fgzJ2DIV
8EyBIppBgxu/22ERWm62+cAxZ2ymPn3UvkYqnMM9JtbDjd4Ew5g2yKS7AXzAvLQz0Nnkpccmmg07
xY7/nZf906GJuIB+M9lVCe18088b9ij8rkZdvQ+u5KcQUR/oRw45c++pvIKhCtNLthDd7v06424A
3wdqMWT2FG5rGdIo/6Lc5Z0g/K14B7uacZ10E8f5tFD8B6b1jahzW+s83+ydPGKd2Kcs/mO9c5C8
ysyhtHLtvm98XHQyV6TNHD7PymWYD5iij1j1rnAgzgoUPUkCDM963gOSgvEIopTYhc1K+34tHDzP
c1tHYCX7AzJz9t6oUDzS0PUG2BcqgJiPolrVGiWWbF1TALmBn8nP+4P4JM58xdgSc3xdx9ttE7rQ
JVQWCr9WB+yiD9/mV2N8IEDO86bLYOYWrpaIJRO7D9TxsVMHJHZH22jZTOydAwsbhn7VybBJOleR
/Jhrap1GMNo+c236DLE3LXe2en2UxN8BNldKQxOTZetxlVTqHhIWrMXiCZC6ldn89rfFelHKvOlz
eXnWByhRYFacuwlRQUDZP16L2VQOrxwN0YRt4uzWnnn9PQZhTDOivi01r9hmPEald8xtFbkXCeoc
IX+FOz7bzFjCa1dI0PqRheUtmx6E+4YexxAMIMUrwX3FAFhL8/09HHdL7KUjpxTq/BziGwUphQEy
McSZuXjLo/XXQ/1Ljys6u/FAlOAonNG/zNBf3qc6JCBliAfcl+lFiTleElVfOysk4YZU9rqvXmTR
WoHjnXxN63iWfVVPOQ8yp2GfkH+W/YyUPJnX9w7Q17rOXvPeaJwn24lHVpaUe9XCp3MZAs8QZWzZ
PFGpR9AWBy/RrhUoiMu0knVB4pzMoUEVkuLQE8Sb8nGRy1Xvl3BABIHWjp72yQ0iTemvwvc6fNI3
+N1QLeyTfhRLabGGYKJh5OOvnbe5dNir+ysqWXg0ODCEREO0zvGK5NUQjg1ytk51v67mBPtAKn0Q
8tPDrbDCz2XSTu2uqRdSxY19Spm7wkp0aRw89ja+XKwStpuo7xXLqJUQiPjKVohvRZV88Qt0W+pC
VnJLHOyNGYLy4hNjGBUMgEqUOR4Cz3AolVADPwpjQ0TLPXiw08qAJGjU/U4OAW/cNXwavDEvYB8p
xtakDTC8EMy3RyCDgZ256afbld5HnVF1snPs0mI+06K2JoZIBXP277wEuQzWNRluB3UvTM1i8Zqz
3ekqWnNN5wQXqV9r/4a2Bt2ewTk/bYW5FLh9+PEObofqnXZp5vvO2Q4Xnz5vRgB6P9unYs3JMIEF
i0r/smodoGKBaACaZT86Ndp7Jv5/4ZceEJ+fywm9gcLMirUL3+KeQz3K0zXRVSBg5j7dw1HYCWML
LZ5Sm97Mj0lOtMDCe3ebE/qD4kM3Fe4XDsY3eitgWkxixM9eYZVHeJ08OAVe5IRWQDInt0tNnc9m
zoJVwGqoMPaT8eifiQNfjnwGm03IU2MV20RejsGFx7IWRKp0RB8RRkxZm+6XTb2I1Eik2oymNbkF
HdeAdViRwOB5U08viewNDBdrCm8SFLcZAUh9++Y1MfU5SiiGSiK29NjrNoXx9xXiQ4U7g1peTUwq
OfRRGdsDTOFvgcZdQ4NnNbhi52AtZfwxy1rqQhr5fRa5SXCHcR6dzTQEr8iEicTTsuyjsTpBbtpD
T8sA/5Fd4YIYNEgvhsklmz5ANJaTfGs37fFomGWIy2QwMmNMVplcktuqLT5rPpQy4B3kFGeMwjJ2
nw8AQXD3k7HVXMEH10YzAsJ4KppvRd+/dUzuTLqK9o7oveujdxGCzxhxwEW2Qu9wLa5uYr43tHlG
e8Qh92Vu0wtsS9J3TPMP+nxZYvWeokIfRXZX5ueVuhgiyn3GRsTgd5ma8sJJY3jscVH91XuyTNM5
xQPUSfUV+DAkbIAT3MxTPi7i76/MDACknZH6VBAhSPfXaYX0GprSnfSw98fU1ofcov5cm9CaER/l
dBPEVLrRk0ZXcCKm9JNR4uW/ZwEJv0bA93Hjoqom3AVQfPcvZE3OIh5Eh9akjPI1RLBbHeVTdSM6
KYyQ6r9JP/gPlBJ7FbfmKffXtrZzZFkYI5VVVZwKHrexcQaZs6nkdQrBimZzomiwsLnrNxP5xzba
VC3o77YdByYOOZW+xfUEtDYfU2tscUqxSvb8EehVXP7LaFadHzspwWcLRXbr7tudSJ+1buCRLPfW
NS2acK4/ChoX2uS0ZaRr5sd0eZq5IVQJeqrVWOEu6xfKrYUOaLAE+q4LC1OJcmqXanbTwpNd/v7j
ByHEAu6BuzW99Uo7PhwAHyvwdLBjTqjucB2fjgVy0yK2gKh9DPZuYtl6HSGb7mhJYxJrqzXZgxi1
jWMxJTCzT+Ga16abWYkHSrFquiNQoe2IHTW0uUkXMOh3c9JtjavS0Lc7yQwWVPPf+6FLHVk7lLgi
adQIOVq9X9ZimGHPNThVkfuFAmFd+DB4EQakJWu728OajjJOLOp3GqkkHae7KIxBwjLRtMJ/xkO+
OpzfraMnNVQUYoraUVPgCI5JSn574xJLluWISa/Gl8RW64Ub0CmzQlDUCWA44AeUQAe0miMkHeYu
6lypQczrSwD0z/xOPZlIjoxT2DL6ex4/p7iXnfDbEnVoE3e9Wf3ASNtthel/hs32VlMgvaCj2ZAG
4IdEXFiSYKn149MsPuZkS+H+Fa4iO9I8hxv8oYkspzM4G/7G56LVHGx1C4XQ/tNxndpzHlN68UPv
tVOlGMC4F2x4aohvHNrt/g65Ne5hsk/XLOPQItQElTv8azmvaKA7BddisGVqIRzwNfHakvmGkMwg
gHlHYr08IijKNx/eYkSNUoJT/+MqFgapeHZOst//8iVNP6gLEwuByBjo3SVjURB5z+OunSmGBx3s
2i+bXBRyi2xG8uCrPhCzv4MtzjnMrZi0E2VOBroRPvxUruybg8Qf/rH+tubwdGqFHdMi2qwwTJt5
BoLcykLk11XUreJsfSBY1bZpwqOhxaWyG+X7M5rrB+M7KV+2oWUpARMsRbHB8UKIgWTufWBps4+Z
OVX0c2CAp4eakKjmolEbx/uQ+moMH7/o1/nGPtLIR0222j3L5bz0OXcOna459KaOPpxVfPE3rJp4
pKJq8R1bXawhmd+IKqLMKUPfFzFj+je3L/Y5Uwccx+8rgzSKUZGqnQjIKwBxK/VPtFqO3YGChCIW
EJgLV2y7ULFuOV1b15uh2SKSVWIsRbjHoLGXQAp6XUCVV0bGUF+I7EtypMrfmWqA2O82ST+HGY5I
H4H1V6/wdNvg5znN2hbHzbL3C8K8zNXM/Prl9kAmpeCeKjoNdXbSofkyd2zMZCjUQNXc+tw89ECZ
MVvZpBkzaX5HGB9PuytslxfN/NnGW0GKsdQP0j6fWSQYRXuFzHhK3eHnxDnjvv4zdbgA61PcQPWc
DUWmEYSiof1re26dHDrVxLpYeCYefZIz3ha/SnM8qNJ+yAS8S+mc40HwxR9R/tjT7LgO2bUr/5VS
SoHH4ctivn3ehG/n1SuPV63290NRAec0CWfN+XhVF5pk3vFY9kTvZWsGZdwbREWPeqSlSInaITPj
q0lmKuIRE0j69Koe4EuzDCZgx4cLwjrKCqVXKnoOZeqe2mMNJVxDdRC9DrioGYVKD58kt1Ffusk3
DqLKN3PRHfT2r5sBiJQFJi0jqbyofMnz/aT8WmW+2+CMGRSY1W7uTI5/XZoIwu6+wYjuLwMVEWCS
12hOjSI9EUIIR68BQ1IG3eUZYklEScMhixxNDhama0K0BboBfKItgcL+ksAA3c7AvvvCkqq2K698
x1jYXMsJO3cWyKcRsLt8ACwusmDS9f/mre8vMBpNk9OefvylHqrPRyjgCGLn6vPL/KsY/yJ8PAlF
hV4h68+J8W2slghK2lYErBuO+08YKbyXjKy93XnIogZlOWqdgccmdsNxBRdcRdAqP/RsT8AZoIh8
3pTmUeFsy1aoweZWv1uTSwnxRI9F0OIip0k3hoKfZxvhqSB/XOpk//71PxvbdHBnXrjBAsFCiS9M
psyHSynderNiX0tcwJmYhtQXSRq+cyDZL5NUv/l6lUqjoaJaevWJaKVaQ9FJEXzhw9XK5Dket6l8
2WjBFpKIBZEbVimxeNWN2NaAZee0BJC6Av+jh3u3x7ID+N01WQAT4Jb+qqCIJ2vY4az5MIheU/rv
RL8XDs7gurM50+IxMu9s+UgYFZS+17EhUTgLgnfxpnY9mU/devX3LFqVqCE6yXNnvpYHQPlp/dpn
0EydPF3bOTpJ/J4PnDXgKlr2RpjcjBe4Q0v+OXinKuYkIUnkIDEv4eG5s9WmvGFQIRdt4OBNd9Vl
U7Aa2HqLIR/gL1UWV157iNYY1Lole7d+3WbPWdDGhfmQJOsxfQx5r7jrPqRn0Cro8S163r0pEljz
9yu9I5trgV5ayz5kQBO5BFAtTDCpa42Vr8GgfNfugXQjKrod0Nev7zIlkO5gerpB9h8S5qaBBf1o
/5EuGgvJ/P+T6PTXS+MVibTrvcQJGDO7b5IzjLDBUOmOn73lolo8OoEPgafNlnYbZp+PpxUIYdBi
O3sRQl8Ru11AWDrQzbiI4l64kBolk/lCyUD9E5OClWLvUXcZXfslVAhLn6kpNh6vmU8hAX3wCQMD
A2FUXulq3HxgXviKSCM+8FUQbilK3WPlF5I/MU1BFchI6bx2iu+MbWUJP/e8bNqcqJOSHX/xNuP0
U2jRQxxesSBMg5AdBfQjtxzl1nVQ9MC7Nu/VntiyGeDidhSpyTdsuNGG98PxnMXLYFCc+/YBOX1B
EU/y0Fr+MEsgROtPEIQCpCXDzzDIpVYSikNPLWeh9ZAORIs7ytTN6FlpOwRmNiMQJi2XaK4ifyE8
0tY/8tcDsYo6zzq+nG6TpncGpQ7ykr4xcDqx2w1nwoMGzgYKT1GPS7+Su9Rg7ol7a5lLeww46R0Y
ifH+D8D1l+2OtCu2RtV5lF8WIlx9QCWgb9xTgiE05OWQgu3Ycj7WEoyAnSrLPi4+ym0fC8UHX+rR
4hkgq6rVQOBPnXW9XbqJWYxLh0zm11LimkLbtgJ2wpowEx1pGINbSG6pm6OpFVoF7WL5CfT+bS0G
YMklTAE3wGuywB9vrz5BT3ah411j3GtGtpS8WQWWjMMz8JxFOINGn7MmmOwtXSfBuzEKWSwQ0UzB
ngmyrfP4QeL9KY4wkW7Qms34KikDO8kf36JR4eq2M58l0NPpJfzZ2JUrJByY2xfBH3v3umYQKXm7
jX9orjHJiWLRXUHbBJA0wElaiqIatK+n7D7KGVj6kqLFeP9DKwD2NAZClp+24VHySvoxt3YvlvL+
w5uCES5YHEzxthQKIzxxyjxA9GyWwtwcg3dRPJS3pBqc90jg3AghROw/Rv1JqgPXLDW4MeU8dC9K
PlsJ7Zbq08ewOr1RVhNFJUf94FXho8ppGxmfdaCdgW3xOD0Z8pj8hwEuMeiJXEaEXDpbgZNCIt5E
GQM759+IX3IXbZZ+LLuvWw9Z0zJbA0JHwzi3xqW44LBch2ouV1w51g9UcKYaqYRlbMbQuUpQ46dr
tPkWGen3O2Wlz8QKFwwuBNEVv4TK+U/6NB2TeC1/R9iTE5dEb4QHSsVkWSu/q5A7ledkEBp7rX9X
gOU9xIjGQvplJeD+8XKSNAy9eUHDn6g0tEdFqSgET/+t4EFNptJUBW5/tNMrfylrHogIfenlZR9j
ZueGNFhK6CggP87HdTSlwlcUNco6seox6ruXFqCASvh1bfLf99BKdh/x0fSeHDgN7ypZz81ggvCy
EzOJaxL9rO1w6NOdzu8MHAVlhPvw5IyGx4UCB+mcDDbxVGxF/MhUgPWJwjCs8E9thSBBXEWeGRxR
UmbWQVuE6I8kGzRTlO9wif5zA/Ma9I6aHQSdml7NGJDAY7ev8PSEc8L/+iGA4mFKkucbidbfWIgk
o/V/7UvCjXqFR48ek3svsp4l0jAkqqILerGOk2HxmWhl4Hxgt1IXwxUiOd1wBl198AGOKT6Tlq83
+Ogkbe9f3k/g1YE0jjiOtahTKRB+3lc+yQQzMoFzqr8vOG/FDMWBsduHpOhfGyoIL5KV7BFXJ3bm
mgrk4OzM0MiVdvXB4z7Tulb6DrIkgp497Vq+98XXyg+2VuG8SNBqqW1kwpYl8We+FIow76OTV5at
waxOQ+K8snGPq0AijFVnRWbfG/zfaJsSQybpkeQF8m9iPKA3gM/tZJE0HcmKcUueQInTeo+9sPit
uIVVnJSLoCPs+jRV3MPn8kv+YjOX1vu6s4WBavYyln3cJI0Mauij7AkyIe+nGTrhYRMeQQJMhehy
JjrxtSoXjDpnpuW2VGNqoG2WOtkRS+h37GeYYV7a4ObLIAu0yDUZNc2oj0UpjCkMe44TXRkJ1Ga7
CUSx2uwbUmYlY4CXnDFknYA+rKPCFzbroGYd8n9ebRSf9mA4TCshaCF43jUIxjnYeL6gUPnYEJ8r
bviMXDWYrUyJUz8fPVPbmB2P23aetsFQuEy0sbZBRfg0wbzyZytK8Rf4m4FrE76rztfosuddZtbD
ay8ZYaNfyloUvz9RtCzZnhoF9NjxecgWJ1HktdOada1l8XhqFgd9TgcnZLxgyc8dTS2RLBDLSI/1
eTQi7zn0Ajtubi/vbHQx8ItlQo/VsyARnw9D/Fbr6km4FNuXghPsG2y7DtdbY5HtQBBPJT7jhWOR
sj7QFRlwxiFydG8+K7zqZE04S9LRdoy0jd/joDdyId925OAux2cmjJO1K/w7g3gNr/BNwuwa+Nqg
NA6S1nXJTTyx7K6wDNK4jtx2kea28GEJ7YxLddofEh3+EDx2Og3T5elhserC9DedDHr8PexCaILY
uHZpiPw/GcUBB8dP/2crWD+yAePIcQ4qchbisZRRdRDYbeSco24xTtpkElVz/CnmboBprZxkPtvI
fZicEmzxR+XFGa81L0W5dMURY4jglEmYvMyDP5rgMHHbFIPeM9hCqtRvKSRSgZ4Q/hlbaO0jk55Q
ZAKYJ9mDwtT8xLcnNmTMMKQq01KrLWbHXJj04LJieIBvMdGkJPtYSpshvhox3hiBtOzijZnG4CtY
oCx+jMfDqtK3YU9AXLKYMfmZLaNoKCtavh/pxcC9GWLctCfF30dO4m+3rdMEPX4tEvEKV7e6aYw9
AVI0U2zDw0WLO/kXE/C76wyvB+8iG0CcpaDFaCwE6M9vOAaUZD9I/NwFrcCSQyWZ1oR7JeMlAFGK
u8es77bGnXLnxfQCihG0nVZlXbw6+7oR2NfrH5bZIhbvXb3Dyq7nv/7NVuNcd/skFz/8Kb6oEgg7
5/+0tHDp8gWqX5Xvt6aTtKoj8RZDyadfB9BQ+h8BIldnQfHv6ynkKCTcP042OycqMQYeUycLtdRK
hsTly+wTQjl7VIkCQhWNLPXgSWbippl1iWMdBSVrQlAOGH/JysIlHKjTFRGwsVw3E7+g1QGV4olK
IUUCeVvviBwyNMUBli8Oj+W6OAFvG+Sia+mgTSPWuvqN4r3AkPhyLfa/ckF3HQ6H2vM9xis2l8Pq
JPFKAf+MMVUWty/pXQeSzgaqAN5CPLOh3lTnVcQSgoxfRhvF89pE8VMdkJzCTmF6kDTvk3/w2gWX
3O1xSF7qeUbdLG2GUeMjfkjFNh810ST0XJcfFuEBdV1bqeKkV6GJTkltm4s4JhT9sxV8hH/08aBV
oDuPg32UI2ulf5eCXwk0LpvnlZ2H8SU82VHfSFxCEFH0V1HMKzCiL8s3M9OnhmypFA8hxpAIhTg2
L38srawVLyCjb+zBCTcJBKwYI01aIDoS7ONE0uLr6TLc3mbjpCNCTVGrMvhBV6QgKUDjUkr4n2G3
bHWSOYEQ+lFo37PAfXNSNAc6mAegCTMm8+FCtDixRXd4W7UqYfmFfLemrd+Ha36DnZCLzunWkzD2
i9p6F7Vqbssmx68i0FvDDA0AiDZs4qu2mqc4W/lTkf4a8E33VOZMAWNBP1AIIlAaQtrww/G8+5HF
Mo5DaCQO3XUdmbe2d5Gh7zIZWgpKW6FUp16I0BRkmX6n75pPGoQMMlbQHb/0o4AuyV3g5RE5ThFo
71B3pJ+E8qAyIOZqB54579u0mK5oxIHsV3L6CkAvifypLZc0YAmAXbAX9yCzL6YbscSBqOQ3trtD
hky0N5rldIG9Zi6hBOXQJcPmY3SEcebdN2wo6st3pTVc41TOSHm9DZyi0dO1Uw3vYMbJIOGL0Em2
PS8P2BD7Er+e49w8efxRsduPBvPZ+62mm/THoSMQHe/NbhqFmdBF7XBuj3MaHWOdAaU+YQMn6x9s
yGDvUqev2eKHDtIZ7waKf+efK4AH2kcGIf5S9QUThBmXBlFzMlPt7FTz+vwBW4eTou1AS62IX908
qhCLOsarofvbAO+xeCQuXAPqjEbitpAwnLdITBRX6Hp3Jq9pBaEkIGkxLPO0ZEPcpHBhiIvzeFfv
sQUBE4C26cgE8Wzu7nOMak3Y5+82WIbHNFhlW8/YOn8WU/9xG5xom6+HO2l5DTk+GN5EPZaPrd/m
4oXRPKB5YJRshnUw/M/XYBB6Weobsg1RgPsDyHm4ryolUjSh5tXeQBAtmxJAyB35tfYbmXg6NI4s
QeZsZagvZIFkpONJ4fIVvl2eGypdKPUPZUGZ4BUlkcEPKsDYKgS/2ICJTf1xOMdLQumwvw3khICO
3hr2YEL1JeHe5I6SJhEijIK9boPn0iy8bI6aD9aFHr1CfR13mcAvLTm5z917k3Jwz2jpRiCopgPd
dgEhzEaU8J76OTDzfxKnjt5Kqx6oA4iJB86DnuugA9jSAffPD/TTtTf1XgEvtbizxPAJAuR4tJS9
uEfC/vNYOhVvvEs+rS3tHyFn0KYtAJifS1eQabWE3zHoZaD+9WPptDjJTb2lG4NSBIyMZRk5Wupc
GsKA17q8RGB3xPhXkMENq2VSguPFjVW6f+wKeIkUAVxk2s7r6cwr/6TQ6Yw+Ue97Y73qu0F2YJ5b
rtBZWT0PWt07z2uYN9H6gBLY3+uXgAEHtApcKyHq2qvoqvWA7gfQAdhJRv0qoO9vEVFVykaImqvk
MOgL0/CLXM4d1M32DjBI4Kl4lAXiq0kzScJujRUwzzUdAZNKB4jaQJky24NHbdKScMgp0zYDu4KD
Es+0STyqWTTf+RotlMj2mv3FqPwQJF83TdWzGE2iO0woXdT+qhdX852SoOtPnx7G/XVZE3jlUOEX
wZjJyKBQN8TSi15C53S+VjvlANNgUygGkAkY8S0oLGccY2oKjoUO2Gk8ZfES9Nv2BQSYR0hMQq4y
u8eCyKpGS0yGXarXEphF04SgO6G8fGmK7IN8l4Ki2/srTiiD+COmTkd3t0WNDmn5RvaySOrmjLO3
K5JLcuxYke7sajBaqTIzejJJwqOaCFBu3NT0JRwzf6eOH1rmagDAl6LsYr6HfQX0vjVz8hNdeMdc
DrUjnlA5gKv6Y+ZRQ5u3H5EhHAARLeW2R+/to9gcw0iSfn/2gzbwpWBa6/cnsvAT/ULD1scq4THt
IBHU0T6RsPZ45ILEfDGR9vd/I71Ji3/QchavdzFuNXBAtpZuACNpC2wNHNZXQT9VwbGD+y6M4foR
nD+XKLASsSLVv3G9zQz2CnslsnRA53Qh+Fj/luT8IYtnH8mpfZ5lOGjdeKWdkRBGQ2PsuyWD/pin
N8hKxj09HwXoWdiQScVLpsSNjzTH5LB8jxB4/M3vrDhaf7gnjv4/rqpgsvnJSV+2Js9R3xq3az59
xCuRGkCm58QtYuAKvD0QvwyybX5225zGcrxZWYRjsbXyXI12EVSB9KNbAc9laZHdPTSILj/ieeOM
3IKKWAkpF7mP7svZ+62uHh88QlUjMbWL9WK5EaSlVtdnTYGlJMVmTTpfwnlZ3+ppP84+IDj5VYDv
wJU3FAcKFFRoKNDjGiS1ixpv+hLqZNBu0ICdEN/JAe5XvNw7g8+9AFZwiURjKEDpkdGUwjtUdBIM
GipqeGkqGMXfixSg2cc0VKQunR2hJI4Kw4/jyjSriK6sBQCExO30xOtVpVR/TBgkIWLbP7UmSYrR
mPwxGAOE+zraQvu0o57ZC/RM6n2WGLVjOIYWErhWldgHkruWGWPPe9To+JkQE/zWon21qh2MsDpD
dRjwgeNy/QxuRchP7U1eVWX3ZlIRu8NHODkvnaeTSJx0SD9pkWKDQ/puQWsUkbTkDIjv2AO0Ei4h
ySy4m6fFivVC977REHwklyAfzCXWs/Hv/DRywcCvmsUKmsLfAelyW8MKIqviaIZlwVd/i6M1+1sf
SkqVPeI6bsVVLAaKdUwdUJmTkmXoUdbSo8rktI0eI2DVYlbhPweynYWxd43Yr9fDKM6Qn+hSmkDB
vvx4b5n9aNM0Q+KZbAB7SE8SgrWFKH8ISn+nBaYzfC+gecte6fdy8Z9tLvUhQtfrClJ/AzY5os1D
WNihAcflfdizAXGJqYAd/cKMFlFqIHOUwdCQYZqcUPTvTVp3jsKIyXm127dVCx2oG4QKvDOh+EG+
MsHLt8Hy12krDip5YDrEyO22ITsiH1wfx64hp5MQcyKIACKU355iHTEPu05ehJY69kkEm8w45dTh
FS2+go+J+soTiQo3fWsHx91AbO8P8bNLcGwS+eXGGFCZbAvSKt76Dlm721Cs2vGUeGfQY731gSKg
+e6UVTeLhqojp9kxUsIpRybmrW6wgyFWco2Zc8HhjjNMFAIqtgSoTAx5fGgZ1zxRaYCwFI8pB0WR
UNBYZFl20kAUT3PvznoDyhn2iMDDFFWuZu0l0f/uGfaOgD/JrWK4zkLhnNy7CO34VS0cR6E6Xc6j
+m1zWvYJ2LX1PVMsL9wXwyOXqL+u6qnvLdHntNlKZ7poUrj99pymTSLxl3U84r91mWCBJpFpAoS/
ba1tIQOBZ4ITWba5lxqOep5VBBk/kV+QezzE3ZXHmPs9glbd5koRGmzIX5NlkhmQLMQQqmqSSi75
17L19ZCV6fX6dX4hOKEQwsjNOQXkADOBiKM7dHrgVYpg/i3D3Dq/w8ZI9qaVOxyGK9u8Erpx75Ax
XwLBn0JP7l17fP3ONQsMCNc1oLcjRifd3DKPL7pzHg1fVW4poiYnmkUQuHhmm/jFUvIblWte2crx
O5Kqsfcc6q9MGGlMK9VHhW2aaS2LczNIPSgcoWQwymbwNQDIIgmxBL2d2Ltr7M/ZZE0oj4SjVtao
svUoC1NQxEgNuN6SDFthRJcn8niZ6moX3fTU0Yd72cTS/rRadv1QddWjDzgLQIwSHK1qpiL3kC5Y
AhtJIA9whwb96fTkDV2u523y5sa4X3sx8GwiGIjcAhLYw3k2Lctd8kAodh7n//RQFGTSRkdNJnGQ
1ab58f/ZMTH0txK484fykxLmWvLIeV4h1VOTB3uGr5ED/1FRC6D+RelS38Zlj3jIcsw3C9+WfLti
AKHXIeKQ+pvSQYF8U6Y0lQBU9t3VvXNDh5ANeJGll5y6z9I8CJAxQqrImbf81nGOdE9XlZ6xhtgw
VoQZmixjsr0WnIfRfSWebtyo11p1UyhF0fLK8aFzxlj3p6BC4v404p0Lpf7IP8TN07IPbufcodua
iP3ozWELfa+rLJQzd2xuvM3TVi4pWkeUke6ah/4dPQTDWUHz6zQnfExkGSWp9b3KGMkanyDqKXdv
lT1avHrOywPWwzEVj1/bKVZTxeSugB44EjUemGefsQ/3YNBxQtaT1uBxZql1KV4lu7ji2ObIVuLS
KW6fn9Ms3TmwCIkhh6yukwOMrWpPynuTjVpOMOQUYD3tdzT+zUyL6PjpGWFBW8IQbF2aYtYz3MGt
Px8uQqqWVD0SDkdv+iotDUEdb6IuuFshjCJtOMJ56a8VSJQ2nlqmHwKZxOHsz0hpKylY1Aeq3VOH
28ty+CXFP/O6G+5dlVRwMuKIAhWYUK8Z/7cPRCJMChjjtNedQZieOPqw0N1dPkL7k5hFYQw+edR4
0Oi/M4zYYgVBdHFPiDL733F7ZntUJAvkbNsN8Sdc57/TN8+/WQ4oZDMlyddG2eeQ2tYlfc1kuHIU
KIpoOICD8s+jnDsBofVPj2DZQxmQw2RF5xP8oH6PTo3Mxo928psgvnv5jktUVorxi8OadmTiUhtC
7k3WXY/FvNb2WrQFOy63KKkGkUhbt6mkWd9gHkRQIONWFwkHP9VPRQ52Q530L0CqBg0CYNrdtUry
uYK7gI9nBnIF5Qvpeh4JGUVbQwnBx8vM4Kr/BAfO5o5DC05GHqyDYahfHnPHArKkHFSeihdctPew
7GHQh+qgpv8EXS9k8id/vEDDbY7hXwgS2Ggv0LJLaMtDh5bpb7XRbaR5KjxhTdogMz1KU1XwpeqW
TAA61okRavlB/jQK1bf8DsGP/AVFIqM8qi1LNsLw1E975mn06uK4KViLDstwG/qymhCZ+jXd6SH3
BX/Zzf4pSQ5bLuDl75mi5c4vcvJKn5BpTILaixVxljU/lNNRiwayCKielhSUmTtHiYfh3fJYucJD
s29Tl8mwFaMu2Hbx51sDSA0kMRNIlbW6LCvM6GQueA2ulo3KNAt/0+WImVFiqYxtqNECz4Rb98OZ
lmMSYX2fTBqfPUK8ef+cw1MP7dICeL4QH1K5OsxhRRhxQy3HK73KuBUmLyjpyIXyRCturtpnq+en
5Tpdi2hndfcfCwAkbTKeh/R5EqmKP0xoC2MfCx2+m9QkM5AbTlcHJyE96RQge2Rq6GcOzwbqWeZ8
itff1isJhXoDhMua6M7F0i/F9sv4JBrSy2zP2IJ2qAQlonOORYVfxbEOGz66gCsvJimyFqTouZRx
PTi5SMWYd7mCDpCtIJpckhZ+CgxaK0374KDTNhg1qOoY0rYsjYMVtjO7NWP9P0TMWZSqleY12t93
bR/4DxMFsSo7jSUivUp3EENZhiAclgqBcYKrNTJbdG2raHV37K2Q5+vMIPR3sKqgh9+Eoc+zzF/2
h8S5I42I4ZJNVhrNBecaC3UaMo3gx0jZfhG513h5aVZIKk0Mihd0K/dYJRCUVySJ2EZZjVKgPD+7
+4h3QqqXQWUtLATaCukCxFz6Ban4/xUhoi4RSXz8m9FWFXrDgLCAF24S25nPpteDntnL8uC/evUH
gtN6kks+9p4PsPNoP/FQ+X8WUOokP1a8bQQ5r/otwoic3n1KdYubwMuHpT5ZOUauFLlm8OTMwMY8
33llxVPuSy7icsMr66UNr0MxqrnQMkXlmVeoEwI4BASWoJbL6kZ7DoeNNnJFb1Q8fCcmT2lOLlyq
xRAtV9HlP6ylJnIo5QIFQCrKGrIDv1eMFlWYy9KMLC8Jg7pB7UxLm8E2kGvq15CYP3SPl7zWWcKb
0vtjV8pY+M1qVpaE8zllzXbokKk3fRW0vM6zXKr910SQ94n8C3+/5Vr/wadsX0d5V9akB0vzG/0w
axr70DrM3OMt2REqnoS0x36RK5Dtun3jTREaLa350PYXpxnNtVmo/NTutefdKsc2mRlRJAlrKcqC
XA0TkfcRJ5Kfaq4QDV+Qmwu+7qHC6aKCA5iiJGJSq3kf6lG6Whd6dpqs62mr4BPvgcquUuYdw8J2
puhbET/Kr33DR8JBErEIolMQwJQ0KkdXiRwW0p42uAGUf5MnKy5FNaSnSXXejwAQbiS7TC3w9R0L
B+oFN6e5YLKnaXC4qeT1g6R1TaNh/wI+nr9qIR92CoIUjK9YgJReRfOv4avu+90+lM3ZKtIIV6Xv
/B1aHjO6S7r9bAVYdZ1wFdhRyrrb1zAnJ+jOxgA9NmwG9eDuszSJZpTwo2hdSTNOWjXzwihlJoZh
dEFJG6pA31kRUAR5aNh/SVWylgjt9/8KO9JhuZoDQGQchmpSu6NXsP3trtw5cTYXYjJ73Rifdw+k
nEaKaRxXSfRcFIncwYrmwT4IxAWWVwj5toSiyJTxdakYKVvs+44J81gPowAtjq7Jrynsyeyt+9tN
ae1m/C3X1efoBQZAPutS3BH5wFj+wdrklGgmY+7zxE2tdgRiUT5M2yrXkcw9lzuxfYQRRg/Ta8UL
GLAnEmMbxq2iSt4wgkTt0HbWPJy1Syx5PM/MGS/HUntlR5VXxUubYqCYOn0baDjg87NOzBbP0pEJ
slcsV9cRBkFEvMUd/O5jZydvs4dDIsvlIe05Qf4J2XtTRymlNuxhuPaKs5jdwysjmxoeDN8OpN17
4uq3y8XdP5fQ8rtaE8003MPz+3BcfENqWGYr1JlgR7bvjNNZWgjr/0KyGNKVpNQ/xA/tBz6I1XW8
ifLDwwiUHsh+sDqjASLCglfHL6Q56T3tBNAolXxjZBNRZxvMidMoq1HQ7vX0ptgdsJnwmWofXkXf
Hc+d6t5UXvEF/4vPjCCwE9auKx2ByCq23LJafW/q61FWbCtN8or9v8iMH1VDWQkKTVuJEGemXcAD
59mv7L7ydTIR83iDhucvCoiy37zDjwymMH5S6Eh6RPnz6wGjk9svqosahihVgityB1lvl179NwcJ
uIDKm9UZNDQh5W3EPnY1F6TMFoXyKxcg4iWi0AWl5raB7BOfxmPWXG9E63qW1Q2I3hXJq3sHeZmx
me416F1WmghUNNTOjmCcQMexO/WhX9UARmlqJbfgR7sRYCZOnsH2R8XJuIuPgtcfizCjnQGwcj4y
07gnq9+J3IVIVpW/frxn2wnqewWmeK/FgQISyp3XrzURthZQOzWc1Lj07y/dWhSDt4tYRhzSz8By
5uvnkm2Mlw6fnI1CG9WDuw1bMdB7x4FC3R8Z/4nRIq0WvSYkpBNUVCs2UoG4r6TXFHqLokUo87jv
+B029T6LrkYCUaqy1v6Mc+9xa3Y7+k3RyCqfnH8MVcwaxNHATB8uDf2TTuvSZu3bo15W4SR8bG7f
HjgamPoLtAYHpGPC7PcY7WahqdCJA1YBs+cke1C5FORfavBrwc1jjSIPHimmGqwv8ess8pwZV1wc
Gogmpj2C9U/5TcqiWhLC20eq/PX7CED4f18gZMMiKgHCP0y+IlJVFkVYyxkicKhC9g/WYoqd6mGS
zu7xQ0awr7JHFwYO2Clvd1OcDP5pYOyjuctlabQQvMJDMsrYogf3VygbaCAkuIcEz14qxnJHWq+Z
yKbeYPX5QBMW/T0xhiuWKivNiCM2bHE9cH7CuBMSWXTSNW/iCz/G746rmChy6wSo2im8BWSRrzq+
8OoXsQND8Y1u3AOxH5eC+HJQVJLhRtTY+uyPLZYrijFQ+4lLlsdJpfyNgngKOHrJmzanCReuqVo0
UN+rXBUaEhJWZLs9JYzinOU61fbRX4HqIph7fb1q9/tomRugZUC6hR7sDuMu9GJdUVVyWMFY1cBv
CDYFWv5uYgF/+zD5Laywn5RDLzbDUKb46XY/Ih+ke4COm1FTR9Yvb7zea67YppFOrTmBZf0h76r+
O+XC8vaVAX0nyTN33epg7jJoh9YGhCjnPkt/cZMZH/LkOIvohiyC3Emg/30rl0IVn8flK4A4O9mz
gAwnIp+J0rjxTpuBR51oneqJJFe0SaBudEDvFTrd7tjDjFNU7JpAuqYxR0erkEPIoi0CWPKQUR+y
Ryphi6GVFSEHIrXUIDHJzccSjT/UY4EX0Dt3mQ7rP3xCCGC9v4xSsUjfo8eVF2UAeclwk4RyGfA6
Dz2qKMLzi44NZCUfyv8XOmltAzx77ui0ex+N7UQYm5LJhLUlN8tOp7rTP5BX0pTl1cVRXbh3w4J3
4TzAxSAZiLrokT4Cd20QNqfVrzN9eYwfIpuv8MSb8X5L3EdIIdsPPV560A2/E3QX4nO+bE9H5obb
LALRojGfYjARockl8PUXAK24KNQEb5HOi2cfn36lwgbWeCGFfY+67O9nbbi87fLH96wLwTuy1iaU
Udm0+6mPVtjlQBw2Yv2WNBKdvY2MqTgRt3XAPdkasTCDpWd36igzLS9/tOf1L8bqEgR9IjPQV+Rb
ZL7YumXwshlislykVh9FC5SvqThKi1bg5XhoesmLieXB89JYtD8ssrVwvbSlMRcw2+i23d9l9HYR
ooCdHAnOhJXbsSdpsi+u7uPdCb49K8tiZMSScXZIWvSZ4hNc7EsnLcBRrIyTNb164b/G6rZ1+rmC
oc8T0tr+QMLFtYILQLLUXwM+1DPA+QNsBR3SS8XyxC1p9l5z7AlRGwIQsIRIYxoQ9iB6tdwMCFn6
6drq2wJWjAqAAlioi7tJchI1Mr6UJSlt0jaJxP/txC9m3yfisRXfgygubAWZ8Vk3gUBXpqWJTsJR
XxdsaB/JbsHMhS1zdK1eLirSbUPOTBJJNpOGswbllY8MUl4aTZJQdBA7+48MmzeWn9Ne1ZbIOUP3
/JNgbBjjGWv57u0Ipzg7+qazCoUwaYsbY44EC6gYfbMuDbuS0unYYa9RypCBJeEvN9sLYMV5/jzh
6EK/drGB2rOx67j2WFWSbEmTZ2fAdRtM+PibqQh0d894uokdN9GgRlM3GqZRfHdjmhAEmjM08+Ot
Xel62DHiyAwSqFUotWK6XPUo9Ezq47g7iimihxhxlGJ2IYl8dQ18d5kTgdrEYcnBeO/9g91CK1v9
ORKGLYfO1NMnperDvz28gmuuBleLo8JQDAeNZxMAyB7/P6z0oqsMavPU0DBFjE8OfhUbPOLXdgWA
5iJAlLpxTiW/GZgG9lKv6l8GIgxpKa+psNvLIkoJGo8F6gmMWDud3sbL351tCQK7YJJmPHivpfbM
3Dy6GZbBQC/epiwD8S+N7+IKfz2O8ainhaH57jmASW02rcMFKW1PCur7tLsyOqtto7mDCIfR/0ng
ViQyJ91hOKWYtgxeR78XrzPkgkdw3i08p64e4+iuIkks0hLyW43tnep4KhMU5pifFgYZs6P19ZZ/
vF6DJtAWc49gZffUtytVThbihuriwbIYhpn3B0UuGRdW7Yvvyn/7PUILXJ5LC4JHxol4wAZ6zAAV
W6yHecv10O00uo8aIrxCQLLxEHBMCOgIF9hR+rMmPtKEEd01eikDpeKkE9vMOLAtGXnsgjpfrat2
wo5fWJFPT8WpqslJmwv3brybfA9BOXUVmn7kr5jb34YOUjqD3lsD/Ro54sMtOXgrVw99pM3B7UT/
KMZvhsRi7xL8jEDSng8wqiAnKJIbbqTK+OEFYJdsZsjKh4G6jy1LfefJ+hKCLRvoI4PDbWtUGk/4
QN7LpQhxiIxhPZrn4CFPTNBg+CXf1y5TAD52RnqB77Z8mrRRDe69ejWLs6Vy4a4Y/KSqjjTs2aqe
GcizUKKT4eXKPKRIePf8t7JBN7dnJEEZriqHBGiTKqlXZzit5tj4PbDzDeW0on8n8GKXlDNyLDTy
6viCAEpB5SccXl5xzTK0ewamIHyc8WNBNOOF5ioHC+UfA/HBpjohRRdbD1KL4jio9LTLUGtj5jB/
ICoGau16SkxIPHv2UY6v0b8CNKXgtq3WbjolGSMp70adJQ+oWtP0Byf5drDBXdOsXzYdgRkHrOr5
WxMI31psXvGq5rAM6fQ9RvsyvkXbhxoTc0fcUVT74CxYIEaczneYRWQ+1LVjAyszuuu/zp74KLA3
s6fP6VUJaYiItpKQI7hiQakDJfgrXm2R0dIBAre2pIxoNHR/8UE+d1ZSBgc0qG5UZ1+jc+cYc823
3mwiwKxQbnqho6J7u09MXceMKzz1M3W1XtJ7UvbiAxpyVztuSB7ULsc/nzT/xOQeV68LejKLsmrJ
O1GldF+sqFrJkymFfmNq9YH/C1s/540s/diDblkxxtlDyXB3rXsWzqzzcv06L1+w2VH7qfoHQdnc
R6XBORY5di+2o+4GTmCs+1f5w4lO0OXMOZYppijfOGyCsgCD7zYKTOIu4pSnLPWepJu2Qts40Q3g
CbOi94D0NiAANM7A47Jehdy0HVbpi8CE6GQZC1/Y6AZnGVaYRRM2HNyTpOn91lXjJ+iS8r2R3RZg
ffaDpjLb5Hyls2FSmwQEjwXJUm2QcxK/xrxfjSMVwfO7XIJgFX8pb1eOxOvGinA4/kXXZ54g/Qex
SviRbxCoelotG//anZHc92qSJyImBXoeCCtoXrgijah6+FXeB2vvDEYQD6teNtGRiEy3h+yYvFsE
Iy0/nd3ZkEs9AUDU2IgP/YqznlWrkOk9PrkXHScpijPfBuoi4z2s92lr5oCHTBBDQu1F4GAl36T1
jiQMxWpRTERJU5yGxq/kGWpEJVt/aGelxGYtGipVx3FgtdPfd1xHpjHh17l/7IZNQHMWL9tFm8O5
nYIOmQtfiICBTQGUqnUMaJkK4N0F/h9X+AMt7pQExYhLgOQrXzM+sYeu0XDDmAgrFoGVUIs67fVn
CeB2WKzJxcQYLz9H4T/b1ImneMIMX3Vf+FrinFgAxPTPJWquEbBY82afs7ibfSy1e6W41YAEuIOg
LQxwGr12/pfL6Y6agpnIWAj7y58C6yikeaZXyP6+IPL+x8ORzPMzbiBA2QE86RTQEq6OzotWocBv
V916Dx5xI2Yx12KrCwVF/uzryu1+P5JxdGLWHiFyDLTGbKmWSkvWwcPwnuk1AWhnBtyKMS0/w6oL
DmGz7dt2/eYmLktbNN/pNrV6+rlqPSbxmnCeX1ihsQYWuC+E1a8kJzn5qCeDkwqt4NaKASfJAbUW
TH1c4z/OTbaOjarGPFfhBkAtZgNOuawbln1TvSkdFSjsSkCc3kR++TOeWbn238Cktum+EmxahwVv
mrzWKv1LWkNtpgMe0nXgA7A5y0+im1GDI4DEdrNp0fRvEeY0i/raX+Rj9aMWj6XQHeaR4UIy3BbL
K94ivwGgg2rwAja3JaytF4Z5i8M662BotjCJV4s+6VsioHvRGoX3nWUO6XFVOMIzLsxFvrDpbwjB
P7wZ0TEaC7AN1D0r/gqzCH39Is7S7t9mVNWgeKQvS+tv6G+UFHbKIRbuDpzcEsDesW3q9puoGxlb
G0g4l26Dd4b8w0ng+VORRbRGl54HWJEOyaCwDkY82jbx5OneMN54wCM9cjmAf65sW+W0todi72+9
0XotIX18GzogVHRW/nbp28GUcGe4kkWe3uzHIsNIIlICxFqAos4OTFm8GoCWCxHxwWaSbehUPNSi
Tj0ZXaq45M2LQ1Af67XHF5B73539BSZgx4AkTq7vVEOQMhS8FojTzzY0c9Dt07NqLdQ7xPZMBjRt
r9JUWt0ko8+hJLmfAgwhm6+UXY+GZyz+peDK8w/E+ATJGYSYlUhPP37Xy5zI4837hmS3Bo8UEh2P
4gXoNHjsZi76l7rJEBmcfa4aoKDVYN9D79CbQXkgv4A9FU3wrGKmpv1wUGvDF3aaJsY45URQDfgb
9Pxq4SwYfy3rRyox2HnphdggzP6DlC9cWEy74twjy5it+CEaXo8uLXbPqsWdyzpIowp7VyZ8wpKH
s7jPnLkTXsKyeRLb6G2lIcquRFkSF3qvBBv5kJtwv1kpf3rcbUnXXCkocjwSqcECRzlTGMuFB5nA
s7LwcuGLREiA71cjn77lg6R1bPYfuFFyU8qQdPopNhIeqStz7jRPtWgq/yiolZ0AQ68zsFF8VxMZ
V9rouNj2DhauM7W/BLNe20M5Q7nhLzdvJ7U5j0iCMtRtFCHgepbLWVD4kQRCjfp+Ii9X+ejsXV4i
dWcJVwUz1dm8ID7SB5eGzOyQnbj9C+JdslkIjXEFjEQEib2sdT3anadOxrCmfxpCloSMzEI2Ggy3
heprlAfGnJETQH7vW76AW4XLaJG1H3FnZuE6ntDVbJKwGr0YONFm1FNHgli7+/clhwAeMp7FqrFA
UpPS0IcvCPmK8zR5oIfJarB45C7TUA2Pk9RwnZCE1hwitR99ZmFnwf3thprpLBGDE872hSi4cDjl
mXstdFt/WRmY79A1YwfTU9GUYAjpwVXxApZcrWcaMHfdgKHqm5Y8rW37BhdZtCrSTTuE9IyIK13x
VfAhMtToeZSl91cNrWDp2qrcMLT2eRBqeGGQ5kt66nGAZEd1zU5/bGrjU8FfTfzkrOU34zBmCQbj
ZdNVL/LMrAWuSP1Omk6ATL1afqrh/OAfWEmlq1+0hKvgK1PqGKmsMJN3QK/tGmQoha6wcVfGd6kV
+gTebXSskIO8YEKVYGXWBcQAxgasrKikE0uVyC1UzgPAFeoYk9VUbXJhtuhG1YkLoGFdrXT7qfzM
33tD4ciYki38jcvSNGmU694hr71tO3sV8Dtvd1wro5qvtF1WPGOk4RegaoHcqeE+b8ttuWVOr4ij
TJKW3COnqzkKza7Wam0e6vaMq1tW/OOuGsF5EZP0OCQ0/tt7u7FTWCXETkFogLK9Gh2ruuKQT3Ua
cxaP03ZV2iXNsvtX7Z/oZKmptNvT5Xtr+n+mcKLcbaPJrCcMerYp+f2ryKCttwQEfT98Pe26Q4tm
m9+ixaTc526pZLwhjvxuWbvUROayDjZtJ63jg+Fd/PUp3RzhJ2zSCcvlq+VhNR1acAyhgmYpHc7f
NYXfk2bsYuX9naP8qRc2FrAuvRDgaXX7aR65DjTPAOjFzHR1Pc4oqnOwoOroiMfnHNwMzB1AV0hy
zY6X2OL+avEdlr/NSo4lgo2Aq0WKDWPHwhgBZ/wpPBexUCR3ecGG03VBgGz5x1bLmUHvq2ds3vUh
NQ2pCavTdCSGBmhfrs0Ku6HlXpldHe2yF4N1gS9L8pt6Ysj9iG2yOnKm3dIHxI0bTWUY9M0s/E2j
nuCOsurAaw5FabMJY5i7oPRC6i/9CLsP+fOTL5fwWDaoLVeiegDrKTfb22dkprEKuGDKzdsMhzUY
9G9YKTgqsljFmC1q3MUvwkAr/4vmg50K8GR7VzNS8wX6mpN39qoc8lF1VtnO/FXa3JhVefqP4ZmF
4VFHVrHYWmohAvavd4vHbIg08yufnx6cCsEYvddzqqgzoGzC9Ysyo6t60Zpwo1xvV8fbg8nfhrkI
/GKhkOf6iLUc/18ocWHIZaAr2x0hxOtIOuLeT6j3aZQ98ZY/2z98Kb9lOzvmuoqDjm7d83U392Mr
ih6fcWruG/JnTY1goKf7+OGK0uno6ChJ8hqt1zQlUqreLidxyJPep0g09O2we7Yvu//DGLqRgN4w
fmLMpF87EgfpCjsQF9JHeN/a1CG1Lc+l+Ql+3fr5lYW34uVPlNSzp4yElMYW3BR+Lf0KxJU7AxMn
pHd5zUPxuxiB5L2SX59HpsgzmU4ltnlh5Eq9PZ2m5JVIQ2PPievNr7ZFQmKJfjUkk0JPy8CjqRXp
WTA6E8UKxTq43Wtd6WmfEoyLMYYeMypPAVJWHmb92VEuGf6V8XigV4IAEH4FnGDMGTFFTqly8nUE
w226zq6fmyuc7vwKnI84xcRf4edDKmfTkn6yXiSIcn5n9H2iSrSR/+R9UKM7mL6CHL2gcPXSbe4f
e/wus00UJHPFAZVjO/wCtYLbXxbV6OG7vHPfuovs61UmVj+VDewYZegyVJ2GlRK9sSsPWRPnyH/B
3PcNXjHeeaWp12VkfrAwfpJ80ldGBlYHxTlDCMzqAe/35gnSxAgcGWuSd2RAJ1sC5iJlNwGBXSyu
phvETbNhdBT/is3rQq3immC9MpbQyNrrW89CEGpd08mr1G6aS9Yn5L1K06ZLJeFPMzM3qFvt+6d9
TW417GMzVBq0n+kruh2qxi/ht6Vm8u7Lr0QKPJueuQju7C+XrLPvq5gboMYMfwAPRCXthEPEaW2k
0CyciMkBJGxailFAHYgUd4m2eoA5DEKp9gcnAnNDX3Nx44aoew0pVxcMsz5xmMbVKmLCdCJjqOdS
1TTKN+xZ6oiwdpRCO81ls6JxhIt/TEfnNxIOpWnIJeZ2I/6u/jTdRooY/QyYA7uFMAl1x418muv+
1B+LH2LZPKQOHHSkD7VsWa7KNzGkTcDxT9gHrtg4DlK2HWqMLqeaWqz3HEfzK5PFJB004GWgKwK5
h3+g0KgBJ9QxmV04HkvKrtAUbGtlBYmrik9m3hT5VQkvAB8hA1p+lFDh4oTqPO7vrEcLVxa/wJjE
VTBj9o8BSGiOc8Uco6q01gwvHIJsexQi4T96azlvqweppE+c2vQhHWta1t64uf2Xrwn7B1TRdacF
LZvDpwHPVag5AbamjaDDjhU3LV5b/1yWsyQaUy+EMdnGBA7jZBaRL3LeXLzYtCNGwHqYxumui05O
GXOVb56ffUI5qn5r1gkxeLId1R0nONZ6LlyXOsmhcgsz13jsPYn7MiRFs70uzfiskrv7mMwmikWK
Vr5R3W5qYSllyd8wohlOQFKZXLU/mMCFnA/MJBYdAs//gyMy4oyj/pOjInd2pYqWaHnKdX/crCDQ
iDEA8HuEgMe+UtmpF97kthUGk9O2JL7E+jSbcvrx2TOo/XvfQXOKJbzFf0L74XOEJKzHd/p2/NA9
2mXIRkup9cbNoZYjjrgcRO4++VD0PLi8Am3rOkbT6IPbFGKyu7ZCAkGvU8oQkvaBC7w/CIaIaKK9
u95QkGtXhzqGSTsgCD5c1s2ZZpc6yuWq0DYW9b7wCPd3CW5BRMXPE7ZQ8CHWKS0SKZFY2FdsEiaH
yKHo4DcmXgTIycMBO/pKykWRVpv0p2LVphfvpNe5J4si4mspKajMzn4MfVPc0Ca36IteQF7MSbB/
+CE25GR21zqWcoSD1OeewiV2k97hcb26LGQJtzP6RVHhgxrjCdbRPLHo1VIyf+D0O0CYzDzZy2q0
c+4y5NpudJ8ru7xSclRRVbQqBep24JXk35I53lQwaJCQqZX9oN4QiWGgBr6m5eQ/VFdnT28piRqk
M+Q7ym0reROtKKbO+k+rco61pfHSteKUia2vjvk5YiPVIbNISkxLCoN5X+WyEBHYkB+GdZ+zt+lV
SJOWIZfAKiPu+NNAPtpBFAItvuoqNYiU6dZIWxxYqowDH+d9xXZiPp3kbGVUezXPtpvooQ+axBjK
vWtLfhI+7c7MQA64gQU98y7YFtzxM+a4CME1hcm0NFUnuCyZelz/7ZlpuPx5VkF7ey5V1TqNIN4M
oi1cygGHrVnbzajSgWVOYG/e+Qkf5UyN77SANMI8b7KrR3QfY+DUbspdxUyn3BXthrKWvsFefF/z
2WYI1ertDyDaUfKhGwPoVFogEv8OqmiVAGydPNF+LfStV0TO4SClNMNsb/EBRSG4L220BSOkaP2U
SVoeWJq7kzyCbSKfCGFEDYz6nthELhGyf7irDX75uoaxD8x+2Gq8Vqwi5AWtWNEB1YFzyBlg+55P
bgrpBv/yvnR3NQIpI4DMsZVm5yGmDXKjDgVOh0MUeIf8sNM9k597hrzqRvTkIW8EpMCGScMwtmC2
2qQht5zRBqQqNUFusr3jchKmh6JuAG5xo+r23z5P3FRRctlmfEib6EnvSzP+IDZx/imlDPFVLs9J
PZHnLgMOK0/Ze29u3JpKjWNKiVrs4FHrdj73202yF1udg21HsRWb2K1fTF2kHpvk8HswBsgRRbOl
QDKVODc37zII8jtZ0dQVwFxBxpD62+oDGgqrOQzSNKW7k73w558bmbXhuBNZcid2iBkN7Uu1sV8P
0V4Ll/fll8M7NS1Uqx9OXXNLJziq3V183ps2sLeM3xYGYTWzyeuVE4kKDUjlnY8QMcks57Pl3lZn
gJXlEv/BCwaMHhCuR5X1RrTypr8n+q+sJRZiJgi9HQbq16DpKYNceQlvGjqhBeO4r+S5Yk0l1s7x
WJAu1ph3PS5BN1e7NMvp9oFkgmnMYCVQGCD4AkyKlqjCmHdIrb9qyhTiyLBT61YOCih3b+tvgHyL
OXmeN7yf+jmGmfyYEDzJX0/iEl1sMQ4HrcmyaPQXMJ/DDsOxsuYix7IBVtPwJxE72d4S7R3ncDtY
N1usA6GjzM+cXc9wFsjqPwQV0CeSc+tc9EEfeyW4f9/eSxFupNZG0wvef4UnAnfoOtPlCZb5qo7x
9u8fhoFOktHvyW9p8j8zVn09DYb9TseMteKOMOTfbeLGF/Kf8SBrzNXf2C5yr9LCnhS05p7vMHop
7YiazcMTeHyVXhfRx7rbqdPT+hbk5g3llgPLUmd//FWeL389Q/TKEbOfu+CL9+Z8/gutUxt4ISsL
kHHlJV1+Ko12QmzNJhHo6RZqxfxRkzSzYFXP4hqBn6L10aE+mQM+h+JGAOeTJnpBNql7YMGiEM7E
yJAe4WE6MndlYeJVnaYq7eKTb+LRCQKbmeTOhVrOL9V80YW+rGPIkaRkcX7gxbw+GQ55Rpo4eovX
o8MIgNzIdQc69F9tjwUruYD5lauV5KV6yGhgPksx+2z4LVgkbVqi/Pr71jFRXfdiglliPqF6fe37
hVjuHVKKN/RH6yY+tCLIzdsC6LoK1BhXpcB2FGl8xHMa0j8Sn3PJb3kd9n30apxdwObeGSxxGVkO
bGIaHpmN/nKje7C2k1T8W+PCYU9D1lA94hSccCnpuqaApvelNJJ/ZAWhX0+ZRNJnLnRCZkDYof8+
SZWPQrztkFOgtoDDNyc0AX3w2j1h19OC8YcvtGdcMIE7Aq5ghJMtlF9i1HFG7sHN4GCLKiCYb13d
R5FoAzdbAL9rhFD5NgGDHWpdmgQIbrURczUafG0MgRD0HNLONUs82zDU3vX1HTH5Ejz8kdcsJgV0
LZeY6XSKfuiZ1SVlRuf3iMVGSD0GNiQ7J/Or8FegSw97qP4UufWkLTyyLikjoFSxEqCQESKSU5KC
VBsqP8tRlddB+HQDNcAjOf+kcoNqt/2Q2OQYsAcbj6RUoUqHAg3pFBFA8aznq1a3ZgSGW5glYFl9
9qdTdmdPVHWZHprqfFlcMldh5z+PX67+8f+fe2gk6TFsnCpiijAs8nDoXq3D86Pv3BDhoqstcJwC
BuCTx42n8frSkk89KkOltLJv7parsYZLBC+QDx4MQDbLULAlo3w0pkiLVC45BeJLdcN/7RhaYSMo
/jH94+2WnkkI4dVBPtC1nkUNmNP+7waifz8qn9eCXJvfj9zAPwfdTXJXq99t5O8Sz13CIj8r+6D6
FNA2Pzp58DE0rXFu7WrCIL628Ox1OutdAQgQnIZzRmSuWmxsT2sDlvbVvWJsGWelOA0g+H2rpi6o
/zpgMtdB5G27g6iwUmxPvVafDcBgvRxb0vPUj3++QMbGWgSKQZxLQoqcgGZGRJDFWaoovWPyVub0
Y+9rcjNMBhRc+ivBpG8W3JAqtdUp1tHLDFTChCe6B04muHyn0JPRnXB7PTgJDFtY/keQ4mGeNTEU
QqkoyDnjjm4xI1icPC1/YIsEwbdWbOxmCNVQ/4E8U5rBxKGu3lluJQjH2kBTJ9i5gQaxgwc9XIFf
NMtVq+nlor4AMj6JxjCIKsCF3J6UYWDeIqmJieHQ0y4uSToi9rYeL0lRGruEB831VRZisBFLqOzy
tsbyCGlwngqjlXnt9jV1W9ZQpZffZmSTKiA780uVOFlhp830GNZXDE1HcjRIpahi2zKg3gZ8aJwW
ord3xPo6mjkrktBt4mK0rS0rtYr+I5ZkIq7awmAJSKrp0AqsX+qE7QheMsRbgSkfUzMYUQk+M1Id
gkKfR7bhnPZ+5mHyvZRTmTiUbZ3dCiOEjvkO/mUjS8okRZPssqBdMgOax9T7Wv8apsdgpzriXurE
47/Dj12o4QybCTpUwoTfCHcg/oMv9wJA2xFkOi40YBxhqQ2hFloqPSZX40XcczYCG3KGG2Kyma5+
nfBEKbf6o/cgylZvyLg73Z1vqj3f06c2zGv/NhmT0ifSjALmdhhydiyBZ3y6yHJZ3iv3lx3fM8Em
ZZFNLC0iNCfYN2D8N+Nfp32ujvM0IuV6x9NRmNi5dfIIMs/EkSWiztU7nsWk++dkIM+MO/UrvTIw
MxykVOcPJbo9cFAqM+Ne+iKU6hmJGRPOiMnogctImOP4HaTFYIXdSWNRmtyp0k+hIHmj2ka9JF6/
b7/0uHGoXM74xd+9GzM7Wm69gt8HqdRzb0kn8UxgKTPcnHaC4ocT0PeMYP7dAgzPACKTPN4nIWYU
OBpqQJqvrHWDFbIDgbp+MV9Dz+RpI5HilObsMCxyqmkcqwf/EWpsArL3JbnmreYLrAwWElglnlOm
UUZooaMKZjXBQkUOb/IjtDQF6nz3ANCRfhQrynSJbx366gHiabG7mwCu5HLGqi1FgArMCYs48F4h
L7dWha+LKWY1xmnrorn7Zrt6gcEvuMhs+VLWU9Han0wu2eztGRLqg/wNepDccpTJHEUP/K0VABvY
SU0dZt7E/+uIohYCqGaHUCul8JX6+sR7oqtArnE+HtURRyXTjDfYlMQItUbbRASHDC7lLhS8R+65
87xb2+QZIvfBoMRTqWObZKw6qwPa+KONstOcoUss5W6n9kwc84gqbLdunC1BEyLAahhGE5AfmImC
5WR7MAfOqa5Hr210PArNWwDljJ6a+lD+T9zL1YFMm5g/viWhUoE8U4HNXj903hRZd1R5CzrZKCYV
zRKkaKTJ11LFMBn6xdqXX+3ADTgpEeSgfCaVuGjrQL5B93xBvM1CLp0mO27OLG58NF9bm5eRKcOM
XnR2csGTTIzLHFGqiicrCVJT4cawTNunqVDlhbLHJ8hAJfir0CpF4kAQWmCCp+xoD/mvs4rHS8xj
uO8Kyl/nQ+v+SvocS86cxn3fxOrSrEcFUFg/ochq0YrwYJHxBIYNa7NtL6VANMvwf8YCNIZgnotg
OqZtN+WWIAJT3bcWtgxP0+we82hiLKTh5dKuI8h2f4u0SyaH06QFfz9HhyJTJOT2uVE2acuZpNw7
RhJcTDBIIU4H0foqDOFF5nrTPLEo2mnWeah+sCa2O6/+I3xDo/Ke/AFvlxy1uU1lpouyyCIwy2Pi
uXYTO89fB/y7L7j7PJ/zq5qu+y3ZAJFluRK/zs9aav3gU4edmepVG0z7A2pAkaLCVxcitiRnFUn+
iCdPwmogQlXos4c2GGyfOSIs4tVKcz3gPyPBfsE7Y2/mr2vQceUSZ1eqvnhU3HzInIyOK2GteXfI
Rqu00w6bMAl9+mmLlXzoWjaGyPJmivZJnqMnf0w3Rn2/Vju+G/ZdSTUJz+97SLwZLTiizII6/dlX
PXWTi64n7a0EOaQuGXVEvtBWIjnE/PgvTR+efapO3TbXzFQC5aT2NhDrXnRN/MpBIJh/VRaVqFEF
uS6C+PFPvohtCPELxR22vQdbgRBxZQV2/QWaKMBPg/SzuCTGlbdrIaHrT+GPb08ZNDjSRFUWqap1
5h/v7TM+2C+vfe3eSgKFfvjBO7cn81h2RFeBva3Dto+qXAG1vkTHAjgsIJh+qELVgOFiCU0Gbytr
hnqfy3jOcs7dc7i3UW2pgmN8SrZlC2/BbibSNh6vSlu8YeBKHUizmgJ1jriO61/E7rjrLpp/CoI1
gupxCOUqr0A41rxz6yWvJRBhSMmveZtGe6sMZa/XveuOAIVMnQRLJY4AhLyYI8nih90tu7AL+KKi
OYonsxKHTUHQDYRVfsBOJvLpBpmZo/yn9A0nc1oFu6PsHyAYwebe8BtTJ1yLoXwnigMLpzQ9TSwE
tHskv8hg8bEdlxYWVtdW1WO1pefHMmH6U0Xif2ndg1buozoNtw6qJPJ6jfNf8EyUgIOgBaq5PGI6
uIRBc+66WbbSD7x3nSejE8x2xul12OiQdYQNaIqbUkrenTPRW5vPxRKDpu4mhTXeYSHoH2m55kYM
8DPQmhEQUIfIz4tBFbwj1+wfmPEL2LpDEvnE8NNwOoOHYZaldhUJyLBerCDTZe3XDXsLeG/dhTFQ
aH8252CEsh7DCDxuMuSO4R4dp2LHkVhqde8cU0ukgJLTJK4yd4uJweJ92VHu50JWRfB93D9CHRN2
37KzO+raPldltIQzgoC2bSK95+IF0GCosR7z9yjaSyx2IQazBaPtq/+pR6yw8Fotcv3QxuF/LOTa
7fSuf05GfVjWierbkysxgVUO3HrT3QQMFjahDLQ1+eczWHGBDZIH8cDjjjGuAU8qzFex85waOIec
7nIkolETgliBK/p39ImpjYPKOAUE3iYjP7vKxZ/t5eUzvsCpX83/Qval5F3kbxgDBzYCicIZBFQo
v0SDdrsK/hCeyNeufYcGihTq+LEwkYDnHaYIWAS9fL/lQaRHC0BP+pEez+CoeYvLe85lKKr8SNUu
HPePYbgSVKui9IZxFjg3ezQe1pKqnmJVob6g+i6YNaQGqeb5MWGMXB6aCVPiHSLEHqcZYHmbypuQ
Dys/nT47mRIEBv+9wkxIm7u8G5YL0bxbwSS2jsfhefKBoG7mpxAvBiNEk25XDGCmbWFOrCdLf/D8
YzBA2oHs+PWDHVeuPkqhGNCTvlX7TkPEUqP1e3t5vxBAdV7B4v+RDesfzjn7fEyN9zePAhnVdXUR
h/UfArgU1G7ivpDlf/pNfje2pe/xTCXZmZ78SUTgsm+rxRmSL+CxaEemeN3xGl9VW/c6a/QTTATa
nrVitR+nFI/6XfP4WLQRy+u/b8xu6689fpavYkiOOFg4PnWD3GxAuqTW0PW1ipHTzkt1iEuFZRZ/
mTfCZOtd69x+vE7MJFR4bwZoTZCNZH86XUe5b9Odioqc0Tyl53FxHf22Ytpeu/Ap/yh2eQDLwQY7
Nk07klQSoPnusSrKU9v+QsrxI8sUaUiQEc9xMKvuXggxgH/O5ydFfbJnuJKAtQNGFLv5Jxqaskup
7NLZuRL3z8/Ebn0hFQIWFrxh8IRf/ftykMMRzYnxSHJZ5tvaTIXwe86koIb7hMWOqO9PCnMzQJKC
8LYxreyrIyVzO84/T7iVJHxM7R++3VpX7GdzCPs/luG9Dg1gh8OG2qUcjXOmx//NMEbktbWPo4cu
cFdFrNAQxhJ8UHZhKjuB3tEV25akT9vqXDfkDSCCi/3EaKD5zeA5dzKkYuAI0YtjVbWe6Ds2Ynx5
MuODCgSBk0veRfNgtjBdnWE6YG/1EX6J+CMMNrr8xjmWgl6kUk6c7v8x4h0WNb6LykSjrYkd7Y8T
FBWnYNGbboX5wj0p3ePaeKsQ8kL6BQVXZug6UFQkH9QAYEUWDxocQLDSqeGplevAAL9bGY/8NuBM
/X8bzB98DjcAx2kkIS+Pt6g/hgZPMxUwlBfQ/Y4yvhzX2ATofdQev/3RbIrd+7koTlLkPbkt2iie
Gi3p7Xr6mH+q9jvVKNFI5Ks4zGLcHJqQd79jG52iB9dW1U6day2bajRJB5PGwgVQxF1uwjLNPcY9
ivXM7embfXX9GYaOixsHyxFrv7036p8B8X33P2F3jqlERplT3KCAoEFOtC3OxbcbwM4d5UzOYG/Y
Dsr1w5MXpLpBj6U+nxGHJK9HO0zlTBDqMIfyfPvv2Sz4rSG07Hd0erkwXqBMlVU87U3Ev0UaMGwt
G+ZA1akXf5u29mcXz/iDjOvEnp3ptne3c11fD/vRvxdR/wZIlJ5AjsMdiObwlpZTrCLWMeuUUka9
twHl7Avoj78UJrFxSzpzJ7Drfv2ar1nIKQvyRcP7ysvSuqoEgjabcKw3vj80YWuJ9rNBkYGbZ7iN
DR5nnN+wvyklbSxT97355wgayQwjjyr6I/e9dfM4X5XGm00t9OAB9SBJFLW+etWGFn9MIpvqTZvV
4pyJDH41fKIrHR04w7Ro9GouRrLa3ByBDL5QvbMTexg/hwsIro7XMMCPGgaun45E8X/PiTvtHCe0
8slFEtg7VifiPiVi0idet2v93uBmvQozyu1qWFjZxsR0drClcEhL2HXowWW936Mm6UK4eXHXc82L
u6rgfKXfTWQnvX+IWxgTAUcjiJ+T/nrXQ1FxPOiYiHLlezXaGX6BlKFlWkp4CssvQIfSQ+T+iQwM
zPKIqlI743c8od+sZAGkmBbZp7FhlFQ+M5URTs67+VzYUnUwPSoaO2PYigmAh846U88EngvP2LE/
B5rwnRNLccRjE3FT34pBJBfQ41X9T0U1zPBBHQdCk2VWqdPmiX/HJbDHld0RHUv7OkmFuI++tEPE
hIZsmOIJpNZRpxPLaKJR1wJK1I6PxS8CWnMmJyVu0wWGBxJxPFZaflqmQqa6yAwUnHfIhKG/V+rx
q8OsnlNiqBfN7SKKOHrDW/QQTbecOe71gCBbVXRjZLgh9tW9vm8xwDyOD3kYvJTSPojKMu87AtME
BwSx6Kdl34hqexPvuhmTSMNlL11CKm4+p0wtKCYWPrl+QuLKsULN66tAw0jC4UzAYzFkJiLvK0EA
q6mOPn7Ttb5S9YoZIgFO3rAIOBky8hD1TIKloE8fjPplTGxOUGaWvuPsrftHv49tfgJ5Leu1+odG
WRvx6mxVoON29qZNTpfcgX6IDO5VB9mVEzMec01oI0LIrmHMblY2fclMcpN7Egdl2zMPFGDi26RS
ShSfZ8pbPD+Qda8Jlb4aVx6JyOaRNWuLCt7jNrvzRBc/nXpL/eb9wkSygyeq4iL/um1V7wpEDAbt
xrpl4LNgDpjxVKT2Zfk0CwGNrQPcOOHQQkgs1Y4FfHLNl6uWU8HpJ6+fg23Lzb+nEANCmOguDHmw
of0HnTzjY6LwZECjov5QV2hRHcUrYbhaCobtyt/3xEcxGZEicv15TDVn98kAhZB8Og1IoeJbFBXw
VW0xk7u3virxQitw9qcrl8x3lOwlOIuDLea4Ec7iiRiPAHicGWT1Br79zRjzYKbFY9ugUzglyXY0
EFUYrrk5j5piX232v5jgaTPD3aV+xYyW4J89yvZShV5kA/DXhFUHR4IsCWSO8vt2zqQFBzLjku/8
KWSDvUWOHiBt57fF06Z25LWhJyKbNqJhZmJFBJRc0koOXf2kbSBV5urtsTQpFhhNtDsvfO7oCKqE
k735OfJr6GIP8qcTwBOTYGrX1b0fsWG7Ma3//cEQQSESIvdEOOtLZWcgIR33BreGtRoEqlQU8UOw
/GnHWzZA5NbhvAqGATsoqyO7hFZXSaMrqcLn5+MXy/rlnOwFkQ/jAmGKZnW0JkyDwczzQfW7gJWI
OHhJXDqafr7TeYoOKxPqZ6Ei2gvMwIR1h5TruCNQvLq0Rkfv/NQRRJWlcbrdKGp4bcsDsHo9bSSA
LX+dsDIgeg8yMU445h82hnNibd5cTKJga1ATwH5MjoDnWkshJIj0Q7nNtVogH6387kb+RbsxAxPD
/Ewwrn8G14QvCsCNqY65BhxIeB/bPUNLa15off8n8OHFJKfGGyHKCr0UcfsEYRAgkZ8x65UExkLf
esxOSghP5oPl1zz2HH5mF9XeIq3l3LWWwiiw7Wlm2QLZO47Y+cBWeP4vgm1CWJ4zs3/+hlpUt/zC
R7BVkeRPSDkW9lMvWRYXIJ+TLQivvSE9o+36dgXTc6kts6wPg6a1s+qRdyMU5e5223rnChHcM9Hd
esdYczR8GID2o3zVQXoAa7aPi+Z1V+JlN0ouRlovWn8GLHUhX5NfaHdkUSI6kmMoxS5nxG7rJsHH
TDz1u+wGgg3CysKZ4yAnJtGoGljy+vQREX1rP8o9EgUo+mG841TbK4bDHjMXhJA4Fmtdmkxl6yFd
9Twm+t0uUVLBcKeLB7LAfnWeOWFm6Wm2PveGKtC1CoqbtSbgwRe93OUl/5cXUIHreZXYF+Ad2KVE
+5cLW0Qy6bFLzoDRjRQ/YbOzKehZOqgo/tKeCqFm9BzVO4vHRPdUm0B5vzXIHFnWe4HjqoOsIo/D
pspSLSEjYJXutn/ln/jdaSNC85U04SRbxlUJGxqVJ14jS3ZQDIRlVVpTxe8StB0xYXUwfwkoPiay
UCDnUsI0WBusRe9vTYD0WKbm1a/N73+AxOgtepJjykXVTsS6DEVQUQbexRxjx0zs+l/iulEb80v8
wH/v+zWx3he545B5fL0WcOhTbKo0k+nL1Jrb9w1Lto7cSHcX4Eig/19skmX2jNYmWl88IzwsqxHE
H6WwIDCD21fF7D41uPXqNDszc2cX/hmTIrZsfpP1qgF+pBAmGg6/SrHQPqjpiuG/rUDfQ+A5EIzF
rJcnsIhBd62WqvQwVWv/FySfyCIFg0zlo/PT54CS8Ex74pO3ujyfz0SeezeYvLwvl2gWqXIsUs6F
cDJSf9oBN4NG/5jalWoxnvyjDeyzEz9D7aMS9UdQew2TIyYz2O1ARyXITAA8Yyo45t7kccvajDgr
U2+L5LFvaK28hfcnok8YlugvYntpqSjS15sWNynRFdAGH5GRCe2vPGWDclrWg3NdCQ/R1esBuHyH
iioWo7MEq5i+F4Dqu/QWbfTxpWFrDRce5hkbgRVGobXL2Az5ZiJX85EoeGiprn6a+ZsSIqFXJC8m
mdLpmglEHafgZ0cCjFhLrV0eYJDdOr6ofnsebpX75GXK4w3jZ6whrPb1HEn3+cmVwvnVKawRm8o7
X4+kMYRvQKsS8FOIqugBeP07rT7eumbNYuAntX9bJorJya2C5akBkCOEI3BDnijfSR1NnKDZwOGw
Re7mPNlXmVcFXKr/+iPW8/1eX99i2DDnoyt3lfYQsWCSKYZuhhhPW0AInQwL9YkiMflKc0+cNv93
WiXYuJERKO0nIoYMHzxabt/37kGxxCEwm7T6yeyIp7REj0+q+8ImNS/6nmz9JAAWno1CzdsrMOYR
9/hb6XUjqwapv48OSwscFEruCFqKo88IUdH6OVjl771qcQkQyU8cvnNi4nQRuvOTV5G7Nvmh+stz
Fr+wek6G4ZbamJ0C7NoJRgHpz3vFezzvcA/i4H1d1OkyrJVKdtjCoZuAjN4q+0TUUamEBs0qTxGu
le3q7zUYm0o5xs0Q/SkXr7tQXtWiWTYPtZ8Q+kIxMhaRyd8vd9VI3u2LVSkhw1qA4WEnpl/+vKz1
pNtVac8HjH+sSmLMop/BhAtVblqxG1wtiKRSEorw5BXYzBfawEaumy/Gcgp3fYtdy1BoHarzmWPf
QQIwz2WKqtQ97RsVdEEKivlLemwlw2/BU3NPVi6ONj1HEv5NI5pzk81jxV4OJFFyqdsuFjm5r+uF
Aap9NNqXHbDLqOmz07dypCNJQEu795Q8IRmL7cGB+ZfgCSb0mCmnH/dU4Oev30fbw4xxeg7Xf81f
D6NwvOiib0ZIXbDzs7jkHcdbzLhqTPiNUd7ChRF5zypZWso9SEEotN1dw+51HDpsObNlMxZeGTnv
RA5ALMWC1yIAtnFbrdGTlf83N7tgn4EZBtg0xalEeoY9nIc1u0cOv9/ekwQikWC9WV+twO9lxM3R
vDzNRYqzFBxku24eV0AEpRWOokoXVa43AIUyrWoWSU7yPY9KQT4s5UhMgS0QJiLNrYPAhDAvHk5A
SIB2Xb8W6inQosmMmlGNa0WR4GAk5yGQzwszOxu4Ss0HiMWKaMCAMBk85HIswVXh1YA81wgYji9Z
FrVoM7IxoEsKfvnPsXGR/mLyNQqneHnZJt/OAxl/SSJxhZn0HgIxtqi8v1jVZXOK4/vMg29WryMz
qEDHliu+J1Ti2f2eM9JLlIMupRFAIZBlVqxrQxbOvfrp5yYgZAq8yptjkQ/an6UzhlSA+/pNnA3t
lKgOfYFpnAq13LiPoNlcyflWN2TCCdfhcEF344yfAutohuK+OonPT+jxpQSTa7V31EU42MqNrbzO
A4DdKh3QYVuI64irSk+YSlU16oc516aKYc4mC+zptlxVuvK5NyxTZnlWtsy6Y+xooyYHDshJ9NeA
+FSw7c27qneIgDTQtjRDjxi9K4z5ofW33B/EjX7L6RN3pypjaB2Pdn2VmPcvnom1OD4o6fcF3ErT
GghtDfmSt4DOisA4z+B3gzquCbb3zNzwEQtji+bNCjGJSiJYrLkaLhoas4tLklFBH+vPdr1jV04y
i4/w3iy6dcVZwMM55R3UeTdMaWBa+FpsmysfYcpZzlAbl2pN+V8vsst1RTGaG3drLOl6kg0j5glh
q52DT1v5MEUMULgln/iVG+Gk/OvbIhs3zwtvbMW/i5nOxI/zCzpIWQQl5GDA0UJh5RXq+bPY/YJk
Y+Q/f1sHkv8V+jtY8gN0eHr/70MuHoaPEvs77ykaQq6T6nju3FahxxKhu7XY+Il0zrFNjHs2bm04
10ImBF+6MRZAqlWODjNxh6JqI316i87bjRWlaiIT4d1xNoSdlJqEbkK5jBejOTkrQdJPAIlNr/f8
4Yh8/PUKTbihXeATrP9gAXKwKdQlE7Vl4i1GNShR+/S1jBJs+GinFvmEq/zD+h3goBtbqdFXV7Qg
7r639pZciIuViqEZXxHYq7rX3f25JqGOaeRAtAknGVIH/9g17KK9U7MJrvoJSo/XbUbeI2PCftbt
l0y232gTHsVV3xWyRqJvsIESg1qjDkWz2v8wL3sCctDFhm+zLLAQEoMcLQ3sFT0WeutYpU90cD1f
qvFzE+mZN2iIsdtAN1qBKA4ylcxteeRxodP73ulM4maAMnrGnOm+gjMpnSScrWFv/hoo/7TpHLlV
Tbbk14xGYTKLdEvV464ocxO3Li+rlki6psnnTZwCdMIAegyOkfVN8AX19HcsdZXzIuQpGMLOl4SF
bj6g8Q8iu0Nzl224GzxkTxkoxJBFL+gFR5aWCGRmOELbJ1OH5dmME/JfzihawuaTJK1TzFfFUjWE
Yz3skx1LQi4lsKEQVgPwyT7xYp8EQtmLMK3IKsKgkkqMSi2MCzD6dl7zxUjCzy+g6UJ2SSChllB3
AlgQb3AxsD6dAyzCT5MeVg9BNqPVOs5gZZxD+xMeDzKfW3+s8U4bl7HktgDjZGmscFfB/sl/YVZm
ff9PAwkj1kSIk59eQgZs+8pe9CHJGw5q9TxlUUuq2sGUpHHSFTdXRLx8vyeYnaMaHwiv+z3RXVCo
xeUC5aFIg3883xTgmkJohHdSBpDKRd3wdnxSrvkWS0RiTEuJjjhdDpE94QSbqVIoqejgnKuzdIve
/OzquNjQ+vBFYoGfBAY7s07d+rrJklYl6fBKX9dnZKnjNGRLFd+QvwyC9vxOemxaaquKCtyLm9TP
EFUtdxE0ak9DQmuCHnreQLXKYhI7+wSBCiqVGcoK2C2QTF2MjjvMG4rZXv8wITlNbLblPNiHlesr
AhhcdIomQUeWa40xP5rWAYU1FmjKHEBVS/N630A0d63plNq2iurm5ssxYeuxf76DVzeGCR9J0/Au
5Dtf6ktGkFLXK8C5fNdbwoeRWq4JLGDOmMA2HA+yboeb1WUSFormhQnYSG5i9el69MnLK5G6Ug4h
PLIJdHMyvaSxvpeAi0+90G5KEu1LJB1yynkE+dhXrXnKFst7atWyS8KDs+GHOOwMgN0CtrOLg4fy
/CrYky1qoAD4JoOFZqRAaBRtXDK0YcmKa512RYnO/ptZSKKRjccN4JXcmUfHq+IPl5pZERG3Zy89
+ZZmKZcAkxXXAETtuyf8iFM42T+VQFtWuD3FV1aSr1G5JW9iWbuw7JsCNOn8d4WmrBsANb1GCQfW
u6p9/TXefcLMnKKGPs7kbUq7z5BdjrORKlL6kdf4i3xfJX6/xaBnT1nf+PJktHBEkEQaGdIdCpFT
c9ffSnafi1ozlC2nVvlT0z1CIXoj73O2r3LGbPF3pAAKfV1Lq9GzPl1KzCvmxW45/iyk4vM1E21G
GaFQ3w6isNhFGs3CYKrlpCG/+5WnUMVjD/w6XGkwE7rqKM9oa/V2mYuFj5qg1yV8p6LvfUwbP1W7
oMz/7jpga4kJiJkse3xPlS/Nr84Kd1D4U5IlrAR+rWVUhshP7B7vnBlUnWGdLVUejk+S1L1heGEO
1R7AFWFUspks3Ol0/qTYG6ZCSq3a0CLKPQJs1e4Z4zBun8A8uumJxi+JqF+gnbTWxE/ZDVFxHsQ7
BkO0FFU+MysKztzbBGfUGBm7wCR/Zjq2lL0P3/thn2okmtSN28b3ZDwOPE+TaVH6hl1+ttTqLs89
NnfnTmqqPofvUs38Wp6zklhv7xlkt5QV+itJPvHJkm7mAyqrrCddRly36wC3cq7RzX2+m12KqHxA
QfrjVDVTkqjL6qGUeRwabPTrlmtaRdJCokntsKG8N/RAvj4ONyv7dTFunMR4cDWugZb3aPib8+1f
J9V3GbphuUDaoUJ8BK6G6IJrsje5g1P1XLg/D85YMuDdbma1OlGAuZmNTkRn02thwsk2aAi2O++p
ZIG4OYXqGauYN7Z5mob7v5Pz5U9+kFT7K5AEPe5I0/VX687jGZGKegDc6DsZ75jaJKPRDHTQOFHL
KdlxHqt5RHuEcvEZ5ho6e+VpnC6nOfBsWOM7Js0unHPgrg/UY6WF4HB0s6dPGFLO1ixd6XVpig/i
/+0qhbx47faGnL4ELhxsslIbYYwTYSjZDPPYRQ2xgv3Otk/cjXq7ETtajdUrv6M+0Wum7I4U2Euk
D8/TMVSgIKXA+00iVkKSA+21Cs/ezh1ZKsConavx2LBYMoaGbDuxiyPkfk5eu/deVumYx7HQUS3F
fDg/srcWhhfbcv50sY4PpfXkcLtXwdaLv8UyNPFeCoc368bQrIwqeCx2XbYabQf02o3tqX9YtHuT
8bBpG+9fhrILqEhVMuA8vSoNQwWccGMh9BmpTO4YePuIKjJ4qPWBch4+SbrRAVcoBVfzhTjtXDHc
SlMSUgmjPWy3xRevjAS+zpcrGgYYqkvu4FMnOJafASu4fS6DRDnmSp9VcS1Q6OCqtuqiHDF46A2X
9J7D7Es7zdQk1fkgN6cOYhHbrU2hxb6zQer4R+hd0rnGzuigh2kukc7fJRn8jHbT0vVAZGIJHyap
bAV/CgXWvc3LELxYYofLDWXXg1aNWdRhFoPr1ndHwVc9B+IG3Cz+OHK2yRuJbbvdOZyal9mgnBOO
qtnczTI+uLnIy8oG/ukVw5D0cYuwRZnJb+Wc1w+ud1hxN1LzhQJaXSpIG9il+JbvQCpoDayS4S/h
AfKmAPtBSmXTdT97wYT5MiL2enaOzCaMlWsHRHKxtVhe7j38/Vh0asiJy9ps3q4SKrE6Q6uWGFQa
pwAcgMneLD3Z4UhCurSinv2kiSYtyUk7SPsB/EschC2lssGHvPHwPkV3g+ylctC4OpMp++lGjC2N
Z/knAgWQW1eWedRhRU0JEMMf+b9dqsD+ce+9CFYr9iBlza2koyPhKrG1VXO47i2ZSCdcjZcL+12i
Z+4e2cqjpsS4MXW2QxXGthL3SnVfow6gwKY3mH+zm6PfURm56Yo2DJKMqkL7eez1tnU7pQpI/qm3
tiDBU0dAOtE4K1LsRTqJfITBsByP4Zaq4XTYOPgxLUuoVOWJfM4Dw6dCQNJIe6mJN+u856GtpiPR
Kn7BrQetINWVLF5nRt3H0LNWBFJ+acwTeGmWzPH5oDVymbxljzE9XlRVuge30n+IQczx+tI8o6h9
+6z5In4l8/NTzQgggDPld/ooiRLL4p7VHQM0NqZ4O/vRt2jqq/2yDV2z1eAS0qYuCm4pZPDU1DNL
BpB6mwyBiQFxWr9ZP202DOlIk71SseT9+Zgx7uzfd4vKnkXYPutZCiAhIKOELypgKN8QZlxBuRCz
mTmLL9vgXamaY3tMhGH3zVN9xf71ADXc3RNGURL19OhTd5OcmnAyMZ48rjmIdFjIr+Twojr6FGXk
hSq6RS66YJLZuufIgaczMTeXHr45G+JpQ+R0oUwIy4J90DRDt9bvOipTnvGBv2SZSU5d/WHutiiW
3a/0CjkS4x0YqxLMpvpCI3vZFKl22IzZEkq4cAnuDnfRGIwIGGFA1pxXTiz/jbecDa8ZS+FLBjJX
iFur/SI0P3qU4ABom8B+rJOzLGE/qxsuhiesgDmvetNhTQ3s9nH0cXgySFybiYcDDHGAuv1hEa5j
/5ibLyxtghhBXe6R9AnBI8tiWwCIM09P6KtfTu6UyrgdckSyoBjDQMkNmRn7LldTpIS3Dz6FHXBl
t+aREk6gHuSHaqJDyzGlLZ+fkELCn9Zl19qOD2AQRp1Wg8cGTzxIuPleZ7cku9RlWfrPL6mKC1Hm
MJtrlSgrWYZsrJ/iVlJT6m5AxmokkiIhEXnu9qHTcOY4i0KEQDYyirMNjdmNISVCb6CClLkyG4un
jC0vk4SlOH9ywmmPN5x2gWo62n8PllFwSQ3sTbD71yF0yGo2Y3L5DiWSOnq52WiCTT79G1qq3ZfZ
AGj4Ddf/wp536827d85Hj2NTdgkSWc7CjW4BdI2wWVMSCgLlNE7nBEVfDIuZFMe3bW6LRHg1KJW9
skn66K+K+/vlNJCrsmPy/zkHCjoVy7174SsRwiBFxSbkw3Ka9U8SwpSGB9KR9IX8nN7fiVmohI7H
e5teu7pwhr+KhCyBjedzacZsxLawRo9hnoRb72GCfR+k9MJkf5CbV+ehRpQq4QB2GzU2hmd23wfK
XSKIcuslSXwfH3jnTzTOWaxGU7uKtOyxDqRMKbSM2V5L/Syao8u7SHtK2c4aOX18OM/w4eyRnT3e
Qi6umhRtQx1tLuvaqOtg4WnYhdgcL5LwymM6727lyBw6L0Nprk+VXFhLH40hiZt83kxINtB8eCHy
+g6DqSfQaKeh2CroDaGZ4vEKFXhg6t6659suK8z4J9e5lFxRQpyTw9Dh0DyF1gno40xdjgy9mmll
pFkTO4GLtm8Fo3e8uj/r1VzntysySZ8OAXOREsgYsEJsX+gSG3ZXsaYYKGl2MuV2MFZm504NKoaK
ZiBgPaeycJuwIiKkbm5DYwsez9ihopgKLZElosJfIYxtuBLfB51gepFNTaL4ApM7G1tME6XdPSP4
oOpHwT4GTJJ19DFZkoDzFoRMdn2wWHkpJ1XZhsSAk+YQZTe6QkAfZ8wrZfcIDsf8jpSah+2mEwdh
yVpH4WV3CnNu5Je+Z+OQINGAQ4rERQRpHoRH/ISPO/DDsJzSyOVeuUovV6eA1T81VlmSZZ0FIBLF
KD9UIb6cY+lNH9QLVhrdRbMf/XOmbdMCLZCshWEm9EiPQ5xB7GvSzkxbSOSiWgXcRq7v15NwtIC0
6uez9zGB7BryYX7RFuYSFih9Lrvrh1HFBXHGVkSDazjBmvxUz7fn+54yG8BvkGFmQP930pTUQmaA
yD8euofz3NxMCb7icJNIcRgRsKnHoqhVHgElnelCsj5IohL3mvBhSa2o7l7+xpIalAzQw3zXbRLy
qkSt/NuqkRYXBxCEu0eHVE4uaOPVhayxhwjr40ACkCov8cZvZoPpbUr26DFYBNibkdpRVy67BFkh
WGMAqwhQPRiT1/VSJSL3ja07L/KHTsN9fV2kyuKI+G758tsinH+08nadkhsfLBbZTtfEFZC+Le28
FmoyFRUcYvAo0X1/axuxr0RJA4abI0oQC/XcR/CGZ+miZ4gGxRsRSajsSlTWq2q0A7rRo+7kl2b/
RVzGin/6Tf1C3yZGpzWo7dM2s9BHZDM0gfO39hgnw6IXPTqztD9zE3PoVNX35BPBxmdddMctQcTZ
PLhogKhaxG7hQHS7IKpIkbnshkVz0dczCW0RUsMdOivd3YuvhZ3zN5QFUEAGivr+NY2/npTkhfMX
otSqF5Qd+Dde2luQ+o6lHdBbBBG/3FgAPV6AXJC7Zm2XQE8M9cEakLGkbZ8+ryAq/CzM1GTDKalO
DDF0xKb6uAUbIbTQSS7Lox4rEF3NHOZa5Zh/JIzkYSeY6zGJHhSHXpKrojCLXgSAV6Qsj1cItokz
hqQnsEDUIcsaSyLQ8DU4QKuMLz5/cvwuEGACAzmX/C7QjIYtSpMEI6PXCw+gFx4jMwLEFxiXfEdS
e4UurOoGPgE5Np8jqLwgDCeQpyZXQNpU3TnqZKoTuEgLit25TKlhGBQ5El/N62lGntSGZy2QPXtp
0qRDDldvQdwPBFIlvbqHhVIy38jJ9jhIqE0g8DamxVvv99B9lmmMd/XBEI5wibKSFXenHx59zgMU
md7m7hRpj7dU6Ybbhw9F/+3FmsLxV6RR1t98N/avqEGiYvnfFzw0oXjBtGQ5FTTkS6+afMGQ96zm
0kHTktUNkVL4nVGE0ff47Fel490atMcyq+YYEMvkBA9/bgxM63Yhf4I0QbvV+clfK2i2yVjHBZLT
UMODAjGZ8S7y0lCQE4j5NKR6LbVOfMSDn76gRNLrvUp1FDQOYHrdIZndmqo9FE52joZbRR+MUjkN
zgVZBfcgz9137Zw3cgcExhO64TdGH6DJ16DDByMu+AjUJW6uDH6mbJzB3ScS0/doaKjRDDzh7Gze
4gawyrTB8tdFWi4ITeDJ/wc7kf3G4/0Ecd3LM56EsSJUFFAw559twbVd0IuuPEJTPqJ6LGOKeO/W
P+CEcMBGsGi5jci1qsdmcviS63FOTJpKPPeP14hQrWLNHUYedih4kWPVZA1kEMhYvH4bmirVK34b
yHoGxmUJPLZEvpuKvNIf2ZQFSoDr84GL3/YAubkoY/gvETB4q9pbN3XFAjtqO9cJIU9Njor5X1Ff
BG5jRa4Pxv9JgmAFjt3wPTH8o2TlYLLPvdQRuEhIuB69WSSHxUOotXI8l2fqdQD1FGxO2V2BCIrP
vwNEIy8Wuz94FKZtlkyNOGoeCT6DqX66j5BO5FcdEb8Q12UyQo8pTnIOX4oueQnrveWx21VV8OQn
t+bfPWJO4a6c/ux11StWbVKvlj8lbe/STmAZVWLf/I1L5H7wuDi6G4koxJvBdVXLBmY99br4JAlD
9zJV0Fo93tilWFv5Nc6Dh6uUkgEps2H6hPjH/eqAhAhlGiywy8Jzn/tSRu3oaWGQcvsMeWDp7jDe
8WNV3MKrvMdEigIYYXeKZMUq8XPOD/tpudnlT+sRsYP39iGFr70LBGEzcDMYbLy1JWfei1Zky1YQ
miYOlc9e1e3RDNShCOxwVKFwIqiBQmOCy/JmzNOxYni35xb7ZktLWQOz81p65LUFjiZRbMmjFTKJ
K31U33HWkmOfEyZ+d+3OtEq6Q0DEc3DI7SDUkaWHZVVeqJU0DecjxB5cUwqtwrPhtwrjZZCiSfGF
e37wjm9+gM0nzd1fnvIY3ILziu3vvr9PYQBix127PCMDQZRHgEAkwqg4eZsPpe3dDukQUzU0ZvU3
gsU/jEJWK92olREMRuiHkpOmkb8uOoXzDeSfkVGQoPAkT3U7lRh4q+45ck2lPIpljEf4HFmEywtB
+3dxfIj0EresjNiOT+wi/3z+3bePcPDmqj5TJCcgETU4bBeq9NkWR4wKP7vAPqjPEW05ih50oG00
BujhgAZ4SuZ79OQ+PsxwoYmtflZopXZ8abkGnFzl4oCr/h5MQ18r56WxvY2UKyqoA4vHa6zZRCsd
g3H2et4W6UWlmeuXaPW5Vc4M8tjB35RvKSIWoqqfqXyF8sX6knPC5VJu/Q1fjZoK2iVsPlUMc3fg
IGX7r2zpBe8ujYdJXqWZxZmeMnMBgCtPpXa4++Pmnn/bWlNsBiuO9ATfp4qh/LnaxlZtrPqxzd8S
5AI67/7p7we7lgCrdyNIk47P9jj8g+LWOL2rmSMcJPN+6c2UVomoNe7TXdCkKVvSfyw9U8l6LTeL
iWtRSHVqgUt51lFqmZRnm8P11+0kQrjjoBDK0GEASjRSBhvs5Ry2JtbFkiTJzEs1WRl7w4T5cnVV
ptxN74TLqvX5xhl2M5wVc84sjReJqgWDmVGat1GgAb6TdPPsfpH1U098EO6Vw55w6SQbo4A8lpNq
vbUc9dLOlv/F1W1fpsGXLLnC9eryYOaDxjUrvwOoeTNCQEBq21SgO0G/QaIRTJqNBT8fjgJHH2pZ
A5eKI+SUws8ARoX/zk/IaVXuvRHxtpUaeocBRP7THRQW9oV0HMS1FuREuLuIbu/JcPi+iubhqeNX
FpXES1GStyBB/xfuukKMUjBY1obLIpOiRAYjxgWeoCCjMosq168EHsa9s0Qcm+42/oMYG6kGf7l9
jpeHMriyvBa0xDhAvGzW1ZO+25moS8oELHCkBvf+iWzSsk+bHrRGDHRKUVux4m/F+QbzWRVPYL1n
xh8ILEuj/bnvqGCFlveVrWociXi4ECkIDtAWmKxWRipEzDPRvxxKoPui63Whb0603uwMkyexj7C7
QScsioHsLDHZ+dg1sf3zqeanAjwEVNB5NL3WXEZanXHyq/r+sKOaxDAQLQDo8iVAhT0VNrQzMcXp
H+i6dT2t4L5grjWVimgykUwX+Ya6tYd/BY84iUQdwb7CTvAoNzpdpFkhHoGz94zkK+mgOv+Tbu5h
HZ5pN4am9H8F9h5ThOZ5zQr7PEV1/+tc5a/rcSjEkpDJuSmzNsF3Jsg3N3UVDfswq8DfINyXQECh
JqFSQq4g3klTM8LF/1teUvg8iEKGflteBghrWbcvTfUWGjungJtLQhlH3Ipi/5YW6WwnYRQnRtzr
srxr/ReafPesZ+9sVvfToCotQpt4shzhFZvLJ6KNrcdX37NMEIoNuOLgnS/iPFwuduRUcaSimE7W
f3sAWizNHsMXY2DfEJjhgoV/gVPrOkZknOI9eTytbq1bD0A6kx6uQQ2JIhTz0TV5hF6/GUv5G/rU
bSgS3YG+m9P6ZJv7L0HGGG+JymNXfOLTSqcfWnL5OxU/7XCndQkVTyNXabVW7wm2mHdRsWfWQAlb
aE+CIO9FBi4LUrQ9/c+pGhskyAzQGEJKzH+C5F4CYCV6WcWSyjM9ZMRG6LTrBZiPMqB80XeZzD0B
FiEVuGbjtyIse8gEJXNiIGKCsQmtf5P+WlnwYHOG8mOyL3RNIGoJ5rPTVDmz8gInDClxSA5ZbamK
uXdC8TqIyMGjo5D2f+OSCMZHsbcgh+15QF3g2f2WVqgIgnZ86+5kR3Z7mXF+CORNGOT8oD2AdURj
Q8wiiyalKm4ua/xgKm7QpS2wmQXyEO7meBj7d1G1H0jn6al+PpsLZLBUwMpbGBy2WOBahZI2cyxn
1DZZqraEANkTZKRXjPMXUJ58cwwny7uuWos1xnLRRlU2Z9XgJJDjh3dUOU8HadxsSMgayeHQfq0O
mVSBp/+cZoMeI2Y+S0u2lwtanssh77hKp1oxuv3hCUI4+wAiMLdmcjP/UcXgB3/kZJf2Mx8QA9Qn
qjAUqp93m+Ua9/U6h4E+eXs5QOs3RwGJ+V6QTcfNIfZPjwXZT97w2Kskr8QD2Muq4wEYMSSi8qS3
WINL23U+nIcKE+xkFo43Jz7Ahr7vcrMzrIJtbpvdp2gHAaICeuLs+98vUtBgf+ubhq4psdMGJ5mb
vjL1cihu8LHkVVro1ukeETW6pfHgjVAQrgPOKBT+PghokZ6ekF/8lzWm9j7TJHwC8wIVdP9DbysZ
3n/x47m3o+l46tvPynRwu8Wo82EcLHRqpMCD0Iqdhkp1he8RGHCuNNdHu2HgJ7uxytVptaoxRpeS
rJDxWJXwdEBxujJIm04fGVrGxOs1qltdVcHAyvpXi95J48ivpqNAhEpkW6N6blKBAXKzn8QPc4iq
QC5+UJJbd3TKqdAqc9Nd52+Aw0+/qQrPOpy7p/MpMeVeBIRldO78ARibj6IjTtLqX3y4mi4FHPaM
ZAv8HtDiIU9/DEeqvoekcKXkV3p/W+HiKn3WVpguVErXmNnP2o5sqIVHZ/lz9NAYkssQCUn4Mlr2
nInoFBAJxqJUfveQXrCyH4kIZ9wZlLZkc1WWjZDPfRClQoofU5PfKNH+6rNh4Y69JBc4x3v/z4vI
fi2x/hRBPNmO8yNrrgt3iGgWalLfxrSmdedhi37K1rcBFJaui7xsTArTaiObKIh8jC/WbpeUnzgj
UfLSWbKq+NEWGhKoItq5J/uPjdSG0OoAXkQ+c5Q3FlZfkrTCck8RfHCwbRN2AsF3I7RXnYGNF0rb
i+gtBoyD6ryzpdnzTYyNiHl2CGQneSuoyox7wg9jT+6K2YSPHKODm6i6/t8F9oqpjnO2mV8hadwZ
bX3UL83woyHOzIhk4+jmQR0VaG6yl+9ZmicYtqL81+n5aYcXgYmFEbW8cPZELl3EHrya545N4XUe
BRHtxpybHbhvt11NnO4OvA6SGYjp5ZINV5K4JXgknMOcX/DrZzsa/TTUw9SDZXY8et0p1TZB9R1a
s4whnKS58R5do3QbXF0R/C2/h01kteI9GfLzcUCJNLHVrTCSde7S2wH+5Uv7YGDmu+d81NlnGLi1
IHNs5dEnS/+Myzo0C6gW5btPd7v8l60YwEX3RyLHD1AtSRTmSQHgrTfDUGfSvvADroQ+CxkHOxCK
or+MtAGL7ipIRULEDl4MsT/g6w+7+UQwmKWnTdUDg3YQUL9KO23SIO5VX4EgX01Z+MNjSId/fT+O
p8xqvdDoKCD49JX+ZjY9UmcWBGl3ixmlFY53ylQPKNghHR6yam+xSmGqmpig0OruvUdSwPIkGKDf
cCJ53IKKmOUAbUd+I2GShJDZkq/Auieb6azZvhcf/+o+C0OCyAANGW4r5TWOwNIam5guUCJ6V8UE
YR4TshaCiaXqnH7V1FCMUp+M1qG739kHrukkwdYgtn4UE43QhCGn92D8Lb8jPD7tZqMsnoTyaGxJ
UTyVBOPhSNstreweh8fN3MTX10L3f04e8RXH/P/JjjMI2JhCX/ciAPYi1Wy/4WDFzhnZ3FJUl7py
/rmTKhczdLBye6paPQDCXcbLB/OaDC+cNGaz7+/nU9TGWD2ZXfwvV3iltxYXYe3NMrwzC0CerusA
p8u1aW2G/1JYCf0PALM5SKjPPT1NGKqcRiIwlY6mq7r+guCwRPS/PjTNBINGWul8CmokgWXzt/jT
OxLpBXJQybK5YVrsexN51DoafyA3blsgYLNQ+KUUueoI30B4BIoCuH2fo5SxdoHMRHzVO2TQHEYe
4iZJJYw3PVwFXBgLApvIvysrrr3QXSQyOjLkRh5OO6vEOXbFU5mW/+r7CJHv40mx6ZC/Mq06wQWX
T9tHl3GrpfpJ+Ptu2vyeJ4M3Kwwtf4TSgP5OAxLubEU6ssh+xY2kbMqYtmixnHsA2fgOf8ef5U2q
wspoIdVCFmSeJIcC5u27mWylLrgrcl5XtQ11nuzEegmEl35qGngYUV3RPz9oRiVzu227/yxoqjNo
47P0aqP83mrmAUznLENhYBJUTCkBuBzcfoF6Zndtm185KoA/sxfhh70yQ1E1C2xJ+lCradpRhjPZ
PSD67Un/kjZkLxGsnasMPM9Cin9m5WtEtAL9a/IncO9l1W2btysqaLOOiDdEhIOJCcmV/mpJn20K
LIcvaFdiTeQdNRhEUPavRL0HOjGplVV6eog46YoO4W9ZJsYKklP8hEB55OPKCc02raC74wEeaSUX
sBPNsIY+wni0pKQqIQB+dBKJKp8ROsxsdX3M+zTpnyF628If2nuNfpzC0gSEFlFNaukfA1Gl2XGY
GmqD3Q0hIyiBGrVld9Q5DJjog+P0dnOGGs/Te8Z4klTjcK0hrFjTpfPODrDqwAHBgY9815csBnXx
gdiIUAs02YrvtlFsNHrMXIhxWeU+ln0cKYlurEYr4YzWp+Nh4ui9G17SMe4XJKEW8z5V1fB52PZc
ZbFC2Gd1dI7hzwLpneQhLRS58v9ApWz3cLDarSGdrt8kNsG/nOB+f/1QmWDkXBbkY2FoS4SF5Ggc
PGF+mciCgdrDw+VpzxvG0GwzjrRi8arfCzeYx715JxtC0gkgEr/5Y0P07AK7+w36lX+tARBZvx9Z
fAKU7ifgUK6HrU1SaO+J6PpHHoRBQ4Cy2OdKl4Yas/+ugsOpT6bOXRcMPheXvnMxQsAwqbErMjel
VJ7t0+DtyQYhcBxDvyXkmOjDRDLzxjGfXbNoxtanDRYMAaIAaFnCVwFUYmLWHO5tpAiGeUZ8qyAs
PWD2sVqLOuC7m2RxkoyXzpa65jvOmz0QjBG5dJOhwQDj8Ta+TkSgJ0UD26k9FA9p4CmOkjnAzKLF
l4BJo9U92hrYLcjZakuOXOheMkWWWnTQXwWMlf/juGGu2xdF7uv9BPCCYkNUcxZWFE5BgORJ8fIG
OuoH5kTL2QLIFFt1xNAJCRjjkl7iEOY4bVt0oEiqQuGhhoY0fNl2uXVOAqGginZv9jDDrGlrGNdv
xGxzMMdTqShHy+PQXXvbsS62f+2F+aqUUqVLDlqw3MQRe9bNgnY3om+ziBjBTigeE7yJ5pZ8MvXC
O8GvJ+R73GBwzE/JimeQRUIZTW8AsMN9PYhdp/qJk9K7IFr/SWMSWJj07sEJNlXDoOxgQUsdq/zu
JDpXdfCK0aMX9bQoefjtNF4l+lOSaIIWzm2Q97NDfg7VoqRnD2X7+KsSFWu9ymI1Pt9HI6qY4rdB
syTD3AbzlOn5TlBxAksOhefqYzDqrz9PTMImq75Iw8A9qIsx44SJk6n0/nre1ZJxAvdPCGpWkgGx
lEZ8sl8i3wshevho8gY6eP2KfB2aif9ke9/l4/ESF0sEJMup6gkOKDEDElBMl46oTXftqKjD369P
9bB9EXFxZoimCiq7sygyL6YK5/CkkcQ0uneObhHKX1r2vAWLLWVh7PSQRKuu7gJmLzdrwLqaZR5Y
tAu3EELKVqf857x8nhMdTBFeDJZQcGf8pwTBmuWK4HetOqYEYTL2DN+TQzFOyfURQvquezCwhYiJ
cxF+yOSwkCwnrfK5vS7qGKqEoEWGxfrJQ4q+3+ua1eCVIb/VJviJbjSzvS6aQNnF92pLdwc+cjH3
ypgyNQD2+j6aiVeDAlhrUV3n/MbaNwvjdmm+mHDgHIdE2yX7gsLcle0tcI+odbl+ZVr3NnC/oKqr
4EFzObrOcPwZDDz8u994as8sCNe+PlGpv1kMcZNsUTW1EwH2tmlUdZT2fLlzT5kGEURmSnlzRAo4
NqfdP4EaQ6zk9dYRiEK+q1bylFcbpfOhEsAxYnek3UCk06qcze3avwGwqPfosSH0ZOFEuc5XAggk
IYw2aq6EOHAWxLLhtSzD9m2IJcjFVwDVsmYr/GNrFXcvgwI+o/76xzUhzyFqABG8XyDQexsGUvfS
nGXJc+fDLrDyn9sW05jo2O2AsZq+Ypw0ZFfldU0oCxZDuR7teORL8li4E7XTfDI5EUMIKHLArj0l
Rc1PK0CRVV9FyaFaCsWMMpKuwNX4cNk32B+RD8LWOWVQUI3yf20aeM1JEMiNOmmSnx4ye8H/dfHa
o+rmCNezWZ0mxQHQQDvvygrj9N9JmxWQHEMoEiyYW4jH3/Tyvn/TZBXdZ5ofgJbnOgfd+sixffTN
sf5ZJ5pozwGEY2VtHI6lKDBpgdQtiutKmB8z1Q7+Ugj6nq2lo60P2Qlmby1IU1PiQbVjGPK986qh
+x9JY/gZQRzPpp1BtSnudxkuh6Pk2X/BCWA5OZ5yFi55tACAWkbiBVwd+oTHYZhPJ1vRsloyxKTL
UFvbaZIfDr5D5SfV+YxKvKvNd+mB1xRAP+FgAKP1is+ZggaaVCtP/sbD8iR6Y85tfImmrXPT4sR7
hjSO4A8Nz/H+gZvs+T7IozZdzL2ZJdqKGoiuNerRhCbJ0jyBurVapt1/GnvzxU7tLlIv5dm+Q37h
qRc7IrZ9mgzljpliFOntvCFGDVbuo35PeWF05zmO4yMf0IjFlU/5QkXSaYigfpCE7yMy/TmXqgmo
SVEtSWohMtVpmdng6xrrv6XFEj6Esn1w81v6BSoGIW2/AacH0vOiZM3C87eGQyyHEt1Wd8+Sf63R
i1vMDqnPb4bdv/v9ggiGIp38S9xQesmta/J/pS3HFJUMDrtmOVuIvaHSrsNmzWnAwc7wU+qMkNY7
VeZ79YH/Fm4JQN9Xofk0wMzmfDQC/YkDREztN1jjA9TvSxAA3UBQ6TOXe/mK8SweHM9o6fBtFjwj
+s1D0oegttI5Qw4USqogzydapDZA65BRxC7e3jWuM37qKvvWmrc51ZVZ9lGWHF83z1QVRxVWh1jX
WudE/nwGrW7K/wJApAL7mobArt/XwdWRyvzCp9uqyJk9Ix0Kuf0zXqBVR4YliPD8I8aFS1yGM9bb
FNoepUYsntydk2Djaw40J96rYHU+kHzpBZeSbD9q5e89SKoJzDXHJlSqbzjI8YlBJfd34ewjotiP
CWpRqEDspyL/+PvueVvVW1dh+Z4oof5te2GywZPMhpKmPZM9lUfbe5RnIg/QvGIBaKE6+qExVBWH
IvFkvmBMyuYkkI4JYxmkNSlWChkWrsVgWKCRzkVafnSdzXDZwkAK6vj3EV5te6GZ54jaz2kz8rIR
JzuGBHgIcB0/4VaknzTvO0nQ9YpDVaMJHG/7bV4SaqoGUcba71/7KEJHEFdS0Ed8JKNlQ3iOPpsT
YSve2Nc8gRKfjOesu/vfZDOVwnccBSZaeyzn++9dTqG1R0OwhFJ8gAnW4mhhc51oS9GbT2x+TQc0
BZJNELWPGhrbqiIZtbxjGVH8UzwgWjBITeeLPy195liuxKvyj+QD/ECqOv0FD9Di+Z8/qNVt/8S5
m9oyfh9ikMt8aMJXApwOoIatgblnfdkOSOrIY18IKNzbCffAV4VWs1SNSykoJzpXAUHdP9kYT5f6
1EEn2kxxWOF2ENVnJpLt4y3Q7GE1TGFX//m7jhpL96HQiFUlios8hfE8JlvFHctTvT9yQMIWMer5
78bEr9op7hgMD3YClXs13G8vAJd4TdyydBksQhVWsP0uwHNnSQqCAoayQlCCEeblfrqeMbIsaWJ+
ppaDA9DS3GJBMBd4TU8TV8YhgrRXMo6mCLX2nZy42as6HcOUWZPBZWeXCxDFgVwB/IWrijwhcNge
OeX4HM6l35f37ACDCjs1R6WKfDqdjrkt2Dv9GVqbzeX0ZXVfEyyAvUF/t6ciZqSASoiov5FTLvO8
L9GzoYYBZ3W3lgQZRMsjaC7yLTmurV/9FScFvPfELZP9COlDgvbf2linYNdtoQTm51dK4H1a7quN
Lvw2u0FG7pkJ5nA09QRB+Cfur8rNUOTfgQuepwr1EJ3vu/DpBEq4XTw521XUlvP50KKFsATZScwC
fFokICCcS+mtDYC2BtjOlN6xkEfHF2aVlx6L4vGmtErfjCH7I/hOCfEZKLhCt2DQ5TyRx/OTHNJ5
cipsVtzl79mXlpS0NuDSDESUE3KGsQsk/hDmh6xRSTJGmJ0D0aLrK0Qzw9Jxpiqg0aWfa+4H/WCk
6gL/LKSP70yZ8QgBjpjp24u5ISuLjPrx38nmcy2kni3anONIvMUFvvG+KIIQrgadZ4rN9goeMDU3
dW4QJr+GWL8lX5tNUeMYCTmWL4hU0ehOb0BF1oZx7YQ0mACmmg91pesa20IqHEcd9Who+G2MfA39
bsSfuCvxM0ENknuECCR7EVXVCIHNEja5vB2CtX9h0fgCcJRPMmu8+k6w6Ijg3nXZZRREkT4LyNH5
IdYJ4pbh+rKIfHLofk8W8EzlvVSAzXZLrO6egTKq98qXZjtF3LAY/To7TzBc7Pfd4bqZaBxOrZwl
dbar1U6TdkDe672UzyE22gk39fCSBCQeTIAWySYGQ2vUykaYNKU14BAovOFNAiq/AK33grZ4xro7
ohSzYStHzsF/fX387DqEmPE22vWtg9CO6HHIBWpUy0QGDdSiZOMoHxJk7Tt9DRhUwM8ss7B7GeMS
e4O/cdU2N70QBHlSLHiHUVdg46O6954ryKr8JDTNMjAQuEP+uBdmqxG0VtmhDTduR5WD2WuqLhBR
B5yt2JVg+wv4wN3bCWSKj5gvTWde00NbmwEpRjXfy5uanB3lTcgsRPwgGMNN518L+t0M04azv+2Y
sKu2xiFCn3xGRZb7MfKMmXZLN0PiWTePTqt0uX9q19tYmtdZor/fnErnsJTJiK1KTKTv/RgJt/T9
RLGT3Y1hFo1oGD7mTNDmsOcTi0QKuBkr6x8sX/KhjJhz7xrgjr0hhgQzPgdNFKvawTLTzd/3xw7w
BBqXcYoEDWgETRXldPPKvijoHIwER+D5q2WPuhDnvsD5DTq+Sp5NaiCkC/UuW7XcAawbkiCKq++G
CwrcNys8Shu8ur8v7MUe61I+aXSkek1V79UBRmaGeLqp8KMy5BpORegnzzOriHd0JXSVH65HlMTJ
7eoxSxt0RRxaCoKj63G9pZJ9tDYCGgJInMqCPass0B+heg7iOOGB8Wl06MU15Zlg8YvxCm1X31Yf
hG0OhH1XvU+b/++1g/rXi/pdqTMuSIgChj3RX4gqH0Mccb209KTt4mlrdIHqmP0sJLbNYXwxKqT4
5M1TmkAO/jG0ciNTN/lnNqRWk4IvIpCi3L4ghGBm2MuE7dpxZjms2QamLaG9pKU7XapgN3Lo6W6R
ZtEBG1iXxXXEDUC3brpB0F3aEK+DUw6If96sjs4OfAe31Gznwr+2zO8vBhxiQw3IB2aNz2ic/RDG
f0HYgkTAJcLag8GbYSlmGQmkIekRLXgt11Z/SGgrSIoEftZOnSdwn/N+SRBZHOi7fAKXRteSe/Nh
Mf5fMK9pQ8LymH8aTAYbe4gLJJEHq8y6ce4m0tQnc45KRv63oVoFG6Q49D4Lvhz8aYBHZDiybsCN
yhIBMg0r+Wr7J4ESar8Cd3I+woJBKk8eQXnRqbYjvtNjw7vEx3hO65cOHblXkB5csAMtzJWswkNa
BObKdF/2+KRM0h1X3Ph8vYQhL4rUhijHrlGpZZePCk/RQ4nbWXzG3Nn9DYV8MFtcGJOgCmDAXXJd
D6ARjmsckWxnQA0KiRPPwueIJaHB3s1vDTI1tXPiJLgVYypnTPQDCYQDsCnuHXWuGeMV0RUgA4MW
7i0x1i94JJ0O1OztOP1QnUhR8vSE1p9zo+3bDIsCGDQL8Hg8/Go9YA3R+IybX7fHSH+7pOLI5Wg1
cd2CxBjp7Q2CW3aoWZ93QzKQIlb5Zod0NuGvl/0i7r6tDStudIA/cY6ZKoGcpIAOVJhmTAZRXrqs
O+5M4HPa9jdTxcaBexAOHrB88toMw9h3gBqp9My8XfrLfIbuckLPZcyRu94iRz1C64Kc4V5Neymj
aS+JL4qkZKDoJyw52v/d+feeU3EqL/KRMdZn7PXJk9RDeK6LP5Bmu7F7phpYn7RBQnQZi2n9S81S
HkYFWBJwxXhduPwKxn5mIqmPsydYAUR/zm0Fc4J/Mff8Uywy3aSLQ6bs2uDrMOAjTdpFpgObUSRC
+nH6nsLBYI5r5KFLOUBXPmvwwHFWgnqIYDuznVNzQkRma2NQPmnoFlCRz/OZZVo1plue4ks7K6Ri
bh6sA5gzWuqEL5hMlfK2zD1ph4zKUV63NpMf8jtUlS4aLf+5Y4SJq5fbDTlU3QGNyTG4Q0/9so7l
QFuSiuZbrvj7P7dPQt2UuXaj5pdhy+gsAZtL8xlfDQq2B2AjcpUKDpUhMR/mIzRGG7eGo5b/6SJr
EEdij7o+AA1iK4YwBWfHAbFElZoWbI+InLB1MYNaxnTQpE+X1IosoygHSishEvilNcrtDdRtF7kT
abzoyD2jlYAispyj+UoL3sxS0kYaSY9FdLgylwIL/NTAFcP4WPFr/vkz6eB3GB3LM5DruupdX4C4
+pgJ8Jd+QUG9k7Drn+JyNJvDq36q1pTOQzD/RbEKRGbvjwMRhbtcojJNHV3hHnWrtK2li517z+pL
daGZWo8Bm2HtXyFAByGrEAI1M+TMkZHe8hKiQ31rW8Ba7YtmREY70nW6lafWkJkdZik2kOE0Yzjl
3+J85Faqp6ljyoXHzNEFJUWZ4jcQqswxaNNu8yVTFqQLJkr4Eb435AlhjBXUycwizaug0JvmZIX9
EnHgSS9p41nq6qXP0myXFdKv7/T6JdgsbybrrtOKQANuFyBlk0Of9VoCj38JauxOKZ2TTP6h7zvR
kAaF5LN+4xnUw1mt2ymT+5RK6tocv7TO/ANE0isMMmZDtTrPh7EG5a6e9ErBPpI4iH6cQcESu9BO
qZkatBU4yJcGcYSF7ROUmrGt+WG0zu/2kMYQyVIfc3IBa2WJEcpKxFrFOyAAjBssTTn9pxvRg9LD
bnWdgWc8xad34T6sx7p98TS2XZ4vhUv6yzvZnQdx4wDt1DT6AhsJUW7OKlA+mNncOUA8ED/jOTfp
zmqvhErMGSz+FEZUxl5iCF+30OPXPGgiJkF36WGWl9AagY3blaxNcQzg3a0HLFpK3QJhRmOVA+UZ
MaOOySuFPp94jyJAsD1e7hvbrLUSqtacEJRKInwYotguJxBykqGxDugVq36ZrrrqalowwfDyKEFk
1hLcy08ZVx+N6QDB7GAks2N2HBQtJ8wYsOc5+IOE6KNbM8yzjmugUq06+UOMtcUft7lNMDCTB6Ha
xUgsdtc+uIUkuOmvdbf39C/K90k3u8gEVR+oVsaEOBRCb9t4dwPTn5lNzCy72VpvlA/kip9maDLl
xv+smWO9oOW0oe0tW1oHEaNQg263QLctrhiVtUeNhDXl9+MITBNovQPGeyqPDGE3gv7qfEc1RpOq
qkKSqJ5xkJqCTEQ1iXUK/2lCf+6Sjz1DFrdp2EtxSPXJ6H/kPVW+RQo6BmBbNdouaioNzpp76le8
e8xXMaKVogFJt7a6apEsGHKqHGd9NRafg6iN4I4TwV5IPfIsCU6EWmzVmAdwu93nEu0aRt4iebll
jYfG9OjBNQZRLks5JUTsOyPhR8MEHnJnZWXAzaPODgKQIuIDoorObZAODxTdYkcmYe0LTs62XK12
ZEWgJ8eWc+Y6vsEFRFXbh2Tb1AuIZA4RQR1auk4WaW58Ji3EV89jPO1bePNCS/ruVqXqHCbyjkdp
B4E98Qnoy9lgAmogk2A9mM+jp3FEc43q2EIW2nMbA1DelmzNjEggaVvYz4HhzhP38nY6QGuLuL6w
WqR4+YWqr9JVHuEY2beTvpV44f0JSi8pYQdanMGDrrjIIyxr8fyYEQXC96rPNsPNhU9mE2ET2AMv
csYL/vg/ojQTD4sG4a0rsgcQouF+nhd5Z2TBQmpYNbXNtpMP55HlMF+9Y9dCF0kAWiQ8chVSxRTU
t7q1p2p6/TlptvZfORo2uSuTdhzcJSxDVEoazI7MRiDtTC965TcdRVZnV5/sMLqKAsigktblWpan
bOr9z5qWE5o+aWUoZsIBj2n2TPvgMRNgBuQJW9zvVs6hc8BsX71PP5hoWBb+CF6Se6uhIBTCL9ja
b+Du9a7+/3WoGxcZuc8clF33aXmCUF/if8/URewbLLHyZtaKxeZeC3aSinJTb3hDSIQ8rIgL8d/n
+UKHx+ZnbxGfIDmH0fgkCv2vLNp63f8ORNsglm1+DhelRMPQAyS7EesvybLUhSc3/FABuSEiPdvV
sdrX/ff5HdLAeDLW3fOxbtzvt7I34BDY/vb9Nf9Mx7JuDDjdk7S16al940yRioIcMG3yVe2TcZRJ
XWYxW/iNQPxrvIoCuZfCyRASiOKF/Mlh+FUrXzmpjkIKFo8I7JQGsDjHxApicirPYssTmYy9K1GF
8ysPTBCOUTsB0OQzsEsQKwyrLniqkLkbDyMWxmM/1P+rtlohQOMZFjytmsnEOv0DPptD92RSkWgJ
XFooxc09bPXBWxpy7Dfu8e7/dkNRUXeLznM1BiuWgCxkuhXgFAy3b63Anh3qLl1miwV7CEV0eFMn
7JmOy5Al9bxF+U911S5BaeUiKZl95lHSRNaaUkIPFIFsrC/8kvAz8iE6jB3RjxsQomuylwC9h1A+
VdZ9Qh7DqIFGh2H4j9vlDjdDb4slbthQkbGRA4OJIV6MXAJPlgUg+8/Cp53ABC9zbr2EzV2DbNYy
lTeuCkBoHZhXRaTsNTlYgNlE+wnvmO7Tz6Na0sgFoKT/W6+pdaIDpn8s8D/aFabdVndi0Zo9o3HN
kVlUXDa9ybb9uthqSc1l3eBtdzQ5hqXRe2Hqp13ZNKyXtMqBqDgzPYtT+572qHKQw2skfrMHx+Hl
iFHGEfj/IwBw7tFzP+HOxI59ZjShqQKGDWMDJsMGeTtVBEXN1kCc0TcVyj9YtOa951ALsTc1fX1s
18AIn9qRfwE0cGQ/Mi8zHbp7maRtARmtKuBQC61Dm/ATtL0Frv8v3/4S7MQLxckgNn7rJf4Isid9
2GqqGFIqwGMTierOJLo+SV4aCZy3tflZGX09SMwOX6tZ+FfC0yKTeEqYrKE43kJFR+G2UjsapKLe
H30arW3UTQVFDNsyRxRQ3N0giIIeimBpKeuz9nySoJUif9tBV1j9rWltm7m/nx3xJT2HKX8mCIm9
muHrIZTPPQXjtj26e3+EEPwI3eKA7NcuLAPvAaFxfdt37RDLjQOpsic/FxsmACg52eiXkRhv3kSj
ke94+aFk3s13cWCUvncvs1B1M/zKdrWeuvqo/KXVrqOiPMF+SSYOT5W26bITfg7iqmw35o5fuNPr
TYTwtzhWXAxEabQkU+//j9b1jUc3U6yJK31ntJNUQOg+1f3aQwCg8jlfmgOl2vJ2uzgCLwOG/LHD
6RWA/becP8hVY/Ty6ktOrHy9j5PXfDPBPyUgaRFsbaY36FbmamVgXXWjMf7tbiuOy6Jd4q1pqaGo
mhLw7lHRVe9X6gmrC1pJd2DrEhavBvvoCm4OuVIMkZDww1FVptZRV8HkEOxBqMVDY4le81Pkd/Jr
eJI5J0HBxkDAYnJzLg4o5ShyYDTHR0lC27exmkwLFz0sBRofCQAnlg+WJiVFbkAwC/F7byXUilZf
DcUCgyf3qu2bgTvfeJdUvA8YbEICBTef+Wk9yueckg1htsCsUK//VTK7w844XVMY5KxLQotIGlIy
vJFekE3HwH/7aQhTPmSb9Ejna9Dvr2xyOapR/KibJBAg9W+/8H/2g0vybRqc9vUV2sn9caJCToMA
0OaNmh6J8IXxSTi+vmuJ8N+KhDJVphmRoIM38e+5+BdIOGk6THBZpvWc9wm2lUC7qnVwzk0pMhtz
7CdSXdg2LwqEY5HMdD1qrgJjnM98j+qaq3VcZdOIGcnjYWxkidgbiZkasAfgds62R/wpPxfmGMUm
otAiK/Eeij6vdK1lOP17LC85Du9Ziy+AS8M+wX+t65o+O6oP0TYNQ08iJOlEBke08Ij39jlZoXli
UMlmbJeONIFkxUPQ0tS8NObnujxPO09ER/vuFXZ1bNv9uZsiYDEg/yydaR4YT9buXJ75e/+8kNmM
FKKVxDX2FrtdlLP0h80DrhGGiuN/vxeZxk8mc5jcxkxhP0Gcy/Q+N9JaqzmEliVvXl66v5jnhJnE
QCM5zD2V+iAldYKwS0q+FZErB4oSZ1TolWMkx9DhguNHLDmM/YmufNVmgSftjtj4x31+CGI4yGp9
ZaOqj81EfcDri/6GP42KHuwOPBgYP2PQy6Y3FYu6RTq6UvvuwMSJajASWr8W91HGvjJtqg9edoc7
aEq4V+HL3ftIFuvtxNMIHk3Iyx4khDj8X3X8+KNKLC0iHxAcVY7c4zSdu8lg4FTEFrmrqM9Js9tq
kVu3P3lF0UjaJ0L6ncxfGBOY08dTn+JvTrRnUnI+NyVctxhWESZEzuXx1RSIhfPHk7gJ9LORxCp1
WmYM0IWxXA27gj8EZvT3DQjLt00i7e9RtX6gZgxr393+A5XHbK4QqtDrb7BRqzegZHC1nWKFp3tu
fxX/YVLJw6GptaAqj0uD+KTQmrEpBZkEbZMLpkdMv8m1BYs+e3sqQm30YQgnGjzw3U+msVDgBkdr
BsJS4nuxn2okwnSvdDGg9+xQPP0+aLM6Lcfd032ulqP9/fDQ9v3zZt1ESGk3KfMSHL51prX9KL4G
itZN4EAm102xoIEYd5cvP9ZoxBJtBIHd3NdGq6wIa07JjnCv1luEWgsBzObfiqayy2j/GfgXVFDf
QEfY3UcWMl3ER7x52jWgOVrbD+s5qWTCKAUBwhZzh5/WB7sVbxZHgomhMDHC1jyWNqgBFhQ0RHLx
p2CD77AeYzWS9UcGc/1BoASoGJCpRQqtQP3JmsHbHs8a8TILrVWES89PYN3yEA85hDh45H+j/t1R
5R7/t43JVMIULQCviVpmLd2MI6i75Je6gMDpK3OqdgjV9pOCd/4m4qAwXVErOtZwr4HEm+XBwOOE
djJMOvejHtuBwyLCT8JjNdMSl/dg7epG5mrgGgeDatZvyUC0BpnbGiWLzj6PlPwSBWkv9iAUpJaa
YluwBjagec1ULSc8Yr0tvrQUoLc0JT/4F30G7vixNSGyrjwk+0cmlToU3lRRFnenvkpc5r3kQDR9
yaDvysiWumW3JbObC4giyqcyV4i/0ua2xm1bTTsOAgEfmHkzJYVk6IugLOGYCb6soUFXejNKXfHM
VVjeviQ2SHth1n+cdvLK8ZlZXuPLs3PIK6Hs/t3XFAkGYCUG5D55HIFmqcDTfu4sFMyDQS4gkQfh
SZXl/zFJJLS0Eqc0PHgaFsMKHVWfLTkRznepi8C6Dojql4mCbW3vE+tBbgUvNGFcPwWWzJ4eZpNg
UHaxS6rpIZYjuL0hKLz22kV8hdFOZluwv7Z4Th7f80UC/NiclAgLA86HD2JLyHY3is2RZcovSncH
gHJZisr8qvkSFAb4NQ4xkHSBqyQPhxlFLEkQKvBqqfsE4M0hCovZDqopYTDxhOTHonKQZpB5b0yJ
LcAMbmRYcUeB5jI0jNW62Sl7ufBWZh8xjBfBo+2AUhWUGMyr34nPXFXk7/CdQnQGNfboIfuWfxG+
aSetKxScfq1elcrd2z0+O7jUT4b4wwDfvNv2OIl2dgQYhgU69StP+bGj+a+09+1esltIRVJoKSzc
f/wisprBiKeheTV3aiP7WCa3deDcqYAicVHWUzp/5BKEMVqxbkIbKVGMXOcUWn0Ai6swFl+qskQo
zwI=
`protect end_protected

