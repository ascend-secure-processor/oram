    parameter   NumValidBlock = 512,
                Recursion = 3,
                MaxLogRecursion = 4   
