 
	parameter				NumValidBlock = 		1024,
							Recursion = 			3;
