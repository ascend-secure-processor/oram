 
	parameter				NumValidBlock = 		8192,
							Recursion = 			3;
