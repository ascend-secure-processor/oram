
	parameter					IVEntropyWidth =	64,
	parameter					AESWidth      =	128,
	parameter                   AESDelay      = 12
