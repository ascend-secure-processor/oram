

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ADd5uFeDYZ+DEq8KIyJW66keeFkHhbBXk3eHLjgw4OIiOeao5J92cOHTBELAhMW9UQgwdTwG68At
++qkwhMZgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F5LMTctMl3znCKydB3X9VK4FC7OTej2McP88vUFBVwFibsxkoksojcccgBu4MtNddfDJhJ6HpOdm
3E5+Nu6QnW8soH8GGAzW7Oc/ag1UdipZvl83pGJSYCVeIAwl/WgVkelDnqZ2Xo/rcp6o7adrGezk
9bJ0htKBKptY6PpWYFs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jLdLbLUlhx+YPuqxwtpA5XyT/uAxfQ/uzU1TVQHghx76BE1CXcX7AxCDWZfOYU8hP0Et6SeTRK7A
8cfy2IltnXTXh4h7hR5tEe75+HZK44zyS794aVQvNbfz4wX97uxrMEGVlmWGyimDlPg8gHw6qisI
7cTZKEcCNmYGECMVQ3AN7v43a7EAVII8IkPvmbzyBShWE2YbCi/zzEVkgYVl3b43PNKAKgvAgjQJ
FjbHyfqsrY0CcqM6RtlAooCGoW8Nk4WdNpkJ2zUAJ7PuNIGWSX0Hp51ADhlRaUkm0S6ONZ5060DU
t+UWaUNOyScPlEU0NadI+tZ+YN/W4A3rd+l66w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QuShWHqXcGyP5GJX4iKQ7yTlLGknHgNgU3wI1Or9TGQFsZw+kaI0Azye+yC+kzyG/+3037Fd//bQ
oAO9Od6RqtLYgQ2aPwQc36LYNzyCOpGqaq8W4qYSyDouvCBFUPOe/QwyY1XTNxojR7RzAcsmtV9k
NWUiuSuOz4BJwSREtvg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VNYbf6u83WiYl5iiQnBQTWDVZioUNw44S9KQQQZ2JxoCAWGX2eiozGYYCv2P7AciLgFRmKbBSB88
9fPElXK+F+8xPoJB/HmsxSb2nQe1D0ntad5USt/ilsepkBnFXdv6qeQmd20u0FoDbDpIhYb7Mdqv
dLsiJm8OkLcaItvPsYfiROPNBfacloRYI/+GQl7qiqo+8DGL1nl/5srJzSW/W6vr6xPtZy7gW/aL
jG4W7nuLZaBpaDkQ4/0tEcXtQZDc6Cn5vHARNBsnfTArlLQKfq+5TbugrkdSK/zoPJoCvCqocjjN
2IrjuR/OoKkiFSVu/8GQ6HsLxRLUb9Y8eNOlaQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62128)
`protect data_block
Xh62JTdNcYWOOCLTvDckJV/rK4VnDhBsKdd04PVC2aADL7yR/nVVTUsA5ZM4zrw3yJ+UOUGc+x4H
cPCqSBGHsJtRT79HQ1T9d/MIggrLtVZ6tCxRyE4PBJaMwMegn4IDSqXz6cI/WDwprY+sLXH6LB/8
lJPypN/uqBx3W9hrrMtIu9wgo6oRdo7qNNXxZxHrebeIEVT4j2bd5oBMQxvvlQN1yqXc6+K+tNf9
nL2KQYQf3PFYvM5mIbSLtn5a4P1Q4c3p1bPl/rhSp1xg58wTerJoyUmQNNf9YudQna8tSXJ5YSHa
bTI++BsPjLyBbXyVhTPYCTQWLGFQ16SHxD1dp/o2s03tNCv79ISGZ9kCNgbTziXPYptpzdfEON04
ZasueWPM+78V9cYMBsHBFQivmMlIgsFEApdHcx6RDOcUuq/K1NeaYe6HPrqcE2efUy7DjRFoQ+zO
/lrWXJsbQnOnPq3RikEWSnqoKFPC7oWbDouFTBXvK1oT/0wId20iQl+ucKwZf/wqnPK99a1KX4bp
6iy86xENvQCDGmSsC6CVygVpxGn5eycV/CPBd9fWV0BJju5wnV/WMYpbFiLN4qNx/1cTP7Ug5G7g
Vi81w6ZY2XvMp0HAJ5oAqC2DVcbzPZh9xSGipSv1qA3bkhJ+k+rPBYbS3zWtG+QCaISo/NroB8Yd
Tk/Qqd0Li7R1jSnlloxy3JfIL454/Fpz+ojRWE920sUstVcg6SdIcL+NvyxAphQsiet4xlFj4h0x
jJv7o0LJktAh7kwemwTnPzrfUUarU8iYt2mw6/c3Rk5TjGDlcwffXQ/4zgpSyDkzmRwdO3U1fMNn
v1bZ7BQukWucfwLNkB9AnZmbzC9lXt3QdQRZkkMwwLJyxMEj01NUTJCx6edDjYCbYyI/DLtDdsLH
e7ToL6Bx3j6LMoEnncXHFa1UCPqNf12A9ZA5i58hfLyrL+h6/GBJAMA4uEzTOIVsyrAF+YquYKvd
P8m+EuVDLlk++6fidTheAbmrIlsdW6f6iMKrlqRbc1zSw8txHdp4OyjTHAc75pWbsS1Rvvfc75Gk
Id7ZfILJEDgmAH4eT4l1mc13q8SdnTu/J3rvN8wGvG9k4k3knn1VzLhpBZWcaALugexwhWmAl/mR
+s3hjmy68iY7yzOEsaPis6xZNpCx9RE1Bl2vG12f+a/o38mxmRkQwPndwH3wrCRJ5+EQ9gDITV8c
WYkU5j8+PoGRbKGM+FELJ8HLSHrGb7iY00Gk3QuziorbdQm85LdRhQei/gXsXY/8crIetEzTUHAL
i3mOVMKbsRxeT1iyHEo98F3gPDb25BVVvn8k0wnfm89Q0We7Yaoonf2HM6Sz4kJxZkxeSYG5hfzQ
UeC8OM6W7qTOnIhL3Um28C8yTsJfYaiiu66F1fCDMLKK2nn5TtYeDGqvkJU3J5jP7AuXw0nT+GLK
VB61dbzfNq4hEjwpQ8FRnckqNAvIrx90g3Ppd4N65gIgTkG5m7gHU15Vw2peL2JhRasC5PReba2l
jPlhwSlLyN7czFepPPNK1C5Rk9nfxIuRey+eBXUTBHicBMwH5QvGhTdMfl2DT/0aL7vbYKrpB24T
Aj2C4e9hYpp61rs1+Km/sYO4aoLbuEUu/jxTPn68QZdp60GGd6X3LVRuqXbnPQ6+v5PmpUR5XhDy
nl9Uc744R+b85iUZaN8RaYT3VHHxZ1ezTBoBoe214rELjtxcULW616uo5xJd15jFaH4POVfhK4zi
PSbs4ZYcwrTdV89B/hpo243xPJAHKXqQf3QkEA+dOfqz+g8WwSWgEylIBug/kG8O/LUxKNlw1bX+
5JVvzn0nIrqrfVFyG+fO0GxXjOq2tidyrGtBOZ+TcageICJulYyMwqhov+OAcdSCuQZmhU74xvI4
FnuArlX3SFEDFnEo6/YRtXGD3oRjb/1LV28fdUCMRzXcpKn0Uky8tkVSCzTBJRu8vatugQhFJUoF
OxFO8XIrIXU4cCap7Gpwe6u2kz1DRx8cbmon73mxY2bHZ3Ja+IHs2v2RDUk8Zc1RkRSdJfWhbga9
3BfdjOsxUv3oHHKg6zWYLhP03UpMW1PnErbKMTCN3dpNVoAzRBDWBI/bZkgRSSynb8HXTmoUNFtE
yg4FSzqVaZpjVd00ENL8czfJi9BokoLmzikw0NXVfvAfBSV5MFI7zVxXDz8mHcjdKrzHQiGeVybH
MEXOIxz29039JdZ9FE2zvwH/C26K1oNXYIE9PcL3Hz8VIYKDrykxtBApigw8NRg7pri9N9FFZE95
J7K7tA/xnHQzzyf28SOnh7Ukiiomf+iitPy9gGuFfySMi/D4OAvqu1pwnAERxWbHiIlR2xYpGrdG
91R7bPBvfEGTK0Nwon+P1oyg0mbCrsAvkAR8iBDWiV4XKLTKuBwdkrV7wQlCZTb/6/X02Px7Qw/4
tiqTrCeXo5QmYFXJ3TWec4gFdKB01QJnBJAbTfEuv8AWUenGb2fSkCOTyjG4+zxlB9vZ3/KSx9bS
0raDkNZVKsrdTtrh7Pj07eTo+T0mJIWbFTUa/8f/ez28XIJeZ71QR2o3STWf5xSjCw7jZ7Phh7Wf
ujvT+KHBr20l6SRV69QbQaaYzEqtOlpZMVkPm/0l80vmsXNzKIcIf8xgBTsTVYrce/JlnVA/qTZr
pERxh3cXQCVDnKVGn2oU04lpYlHYzR0VVbMh0lY4uIjtPBtrn3CWDCek32uIWHreoKZykoT2JTNl
u16Mrza15VVTIAfXJUdtZKeE668+a2PVJcM7OWVJuUXMxMXj/gZA5anPrMR0bh6q4OQsmHLBPh3t
OqbISBCD5CFzL4HazjKiKN7g+rdmiOWSioMVBrPsr/7RbNuiw9uWQoBZ5ca91FzXPvg7UCHcuqDT
zNzyJ0Gy+YQ6dVUXgQ4ZmP2TQlHeB4b8DRoclFiZG/PrH+VBPaQoycaL8vKeY+9w2x4S0c7Oj7oe
XuFVzwMTgzp20hIkRXQR2sxgB636/MXWQYqYXuj7ZJMh9PXi6TH6DVoB3qPTbn1gmEW45POry31R
pJtZ0xFuOHII3a/I1yrLuADl7dhmjMTCgV1m20eHB+Lprl8+M35s5NA2YnIC8t21znJdTsuTlGor
6wKlGvp/oqEMaKLtAnCo9i1T9XGNEkVP3zdjVwfmeq9gm0khWTP8OCK7FojSwTkLSWNErQ276gME
GE/rBYg6sX50bhW4IusNPpv6tzAjDAZoJb623PyiID9umeCk/dmbLBUfaibTevCs6Jk/Lg4gASWj
hOd0XaU8jcJoYzGu8FmAuMXY/PDWBXUj7Uj2T7GiPccRdskA6blk4y+RvKzT7qusWRZEiXnEkujo
iTP+250L44bkZD8/QsOoIcRa0Dc+xKz+MXhNVi3O1665waK/kJLQJF05kltWmfH0CIAiGRxiHPpf
MVdBZn1KQK5Kz4cGtzxqXls93nZS3dW2CUSqQ1uIRF+YasO30HIVXKkna1Xx7gSk2G2qBF9oVWbe
/+vgMGMwUUlEbB9CGWagbMh+EK2UhaXOkfHHWgaVue5VAmvnTPJ2Ns2Cx4MIc2sQ+jzqac8Ldrw1
asQN5BsGjdJHBXQwyCe6HEmLeifQ3yV94HZ5HrhDIpSxNvPhbVhw+DTAdUMU6Z2KJF2noF91D+PU
pw5TOWu6nDZK8XVpjfe54kZ0oAKuTa73B3qnmaT9vGS0mXyuR9F1Z/ewEQLWzXTRjFS9SgNLRtey
qhlY0m52kkU74Dg6eDBRtN8eHdcdwi3BOspBU4a/Lz0+HSkfPPew7l/x2yij3oL89/FBp8tXkye9
GMzPC/6HNBzdg0pLY18kub8yhrkTdebPP/0neKaYXNIx0sSblqYG/WcT5uUxucnF4zQ4yEFoD8oX
VPSHCSJ5AGeT76yDBWPFSTkKB/cNt9xha6+FFk6nicOT3XUmxYJj1Y82rW6MLL3reZod8iByXlqu
gZ+lPo/gIEhgkrJG3F0EIflHnScj+mvLsEc87JIEP5tmp8fgi/LnIJiYstEGGhvD3qfuDhty0XTq
vSDG2tBRSmUaNnl/jgFGn5hK/rk53sMVSjlVcJiMj1u4OlGuxoxbByhk4yk4YLCBQXN5FF2bMfOP
qQQc4bt4U2QtfSX6M7yJ/F0yYrq59aOdF73mtA/sZUW5Zn2UTA5hEKJ9jhJlXWSPAtfAk8DFfjZ8
hCmT99/h9lhxg02Zl26ItzckLioNynEE+4mYpYVY0hsCasLLTjC6zT//nPVxnmBSYstuoZ5l9PBw
vr4cHx3xeyCo8fdSYxQ2GzsNrGIpprLzXEY8BPDWvushIl2BsLtcy4OFaeVgkk8aw3ZDg8pNmHQg
C6hlrzc99jwPwKkKINHJkdnuL/gw19HbZH7s7QYaqqSvfV4Zc8GkqJDLN4c5fLeMxUAVsMIdMHQ0
ZdD08sSBUEPSdCqasb5UKs2KiPe4xcdUQg4jMUUAYPyreGsU9x8XbB9xlwKjhM6OJf/JM0Eg+LyN
Hv0gPhurqJPiZt8KK7HVKy5umLOFLAmsT/vP+7amb+GqDHM5Bk7AK8NSc8G64t+mDtI++zpzVKrK
dliad1jpOtJ9bfdWaLOHFIamoHMphgowHqxHdPoA8zKehGXbxPSN1Tc00QYKglnTLvJZef6XO57u
3JcuAwgtsSsbs184/EoQ7vGe48Qpx9hBngzJxziGjYxoDNUM1TKrdQEi3GtB1yoTVnNX0LcTL1op
gCiny0k8faPJlsDpdRfhkfZJSNJACfGC1wpPeKGIVPxDZdo1dzm8VAwrcRqmDCvD0whTLXLDBMV3
NUcTqkqG3CS6XAYedyPTMzCqSjR+S1p/BZR/oVPHKLlqzg+XufPL9TankcZsSTM5EZVciG/39o6H
iUZ5VP+eeJ4aodFq0o2+7PJAyX6ZjkFhA+Nzomuy+ZORxW3xSaQlbRTf6e1HJCX6vL3p3n4Pl7ok
DItSxPXiWpy6F7tzuhAG5DWqNl140VM9Ub36ltBnOWddLEWxzar6YFcv/SY1g84ZMv4MWlxSgaDU
9uMoiz/QcmnBcBMCQoe6ePdlMlUEBSjXhKWmJeIdmVV6vBuDdI+8VqyQTLX5KzOs3FK1WnNR7Hbc
qx7w98vXdECeQ9QtIGNF3Ww4ckw8t+CqVFakLpuJhoj8ErpslcUmzULlyBVO1IsXepV03X2ONjKi
Q7ne5hhi311kLcO9+rJrK0HmeNbSejZlYj3g9SL/yDGS7eOjnJmQHxUoKfCB8eyfy9nDfeG5iHYy
NnXJh8r+SWVKhDyRaqiidDL0W+7eS1V/7lIujj4F7isvaGXK5MLkbBGwbUW1tK5U8EWec0UFAI3T
kNat49G0wTUTFBHJ09LcUGEvXAJ5ueq6jiViVEQSgqnE5/xQvCoa8tqr60Ih55mBHewnOIEHIhjB
wPWr5RJlZGdvirWBuuT7xN0OtQQ3P7DvTCNDfXd/WFgGfoV7KukNp/U4K3w53lSdvN3JKcMCCI5N
HaGsGTH8cnHubNGyIiL8HTZNHVDAGawgVbQzVigSv4fWaq3TyjeeDIfeEAEnbAS3AXRic6gYuBKI
pjUYuH6InNmvKAIQYza/jsr4zT22OpPNE37Ys89Wjf8W41lla+lgtQueUCdQAtiSOXcCYAZMIEUO
njgNPNTqLG24k+k8dPhSduy7FrSrpoxG8UFVEVFc09/M/VyykAjDT0lyXX42UKdJa0f5Cn5SsxUS
e2KuhArdcIBt1/4EljfAA16yfHj1ILPJYsKj/XM+e4hc6+Sg9lojmZKoHREERFbq+/5DL3dUYozw
bekxa+f4c7tUl4dqMmEWaAqIQ14veDAiKTIOjBnR4kBp8tDcQ8j2v9L7SCbg1vJHGSVJ9H8KoZ6A
IcGQGGH0/B6yW3pSw+p1/D809cei0g8XP/Pco7iT2CmTZsug8SojgT3PUSW+NdWRvWlXBqUKo0o6
zzFhulMupkMMIEy66mSpqgR1bhAOFpE5FnZeKAVy8SWTDjmU/d1AJ+RaD7kkNQH9rMXZ5xkhQeRk
dOiZj1NhYOKscEuBpuKg0edzdVh7VlpXnjRjLZYWi/wxpT/hN9Px+fieqoU3t6pYA1U3/3P5oNLt
fTIIe1hd3F3S0el1cCKtJWN8o4LYfkrh/H8albPZMQn00km1gJ+60xcFOdxof+JByYLL5essxofl
0gGJn6pyiXIH8dnPC+X2rpyU5E+4nCQvp8eRVnjd7nhog0zKFyYjMMbm7hDueH+6gzTGwzwXC04d
FmPoZs981Ednf5m/r8MTecN70ZuzsEuO/MiIa9vL8vswDnpDbU1hklDHHld2h+sYmFRm7+sjQs90
lEyxBFw/SUqzGYxVXlOSyFcc2BxOkhBRoZC6T0H6LqPTlOq6llORQhGb5Y5i1f1PO4y7RwfevTsh
sKhwgzzr+DXlEDOE/5aRdGLaxTCJS0YPVvTbXvaWv43pH9atkd/AHmLjOcW6+xz7ZJGzEMTHwVcT
VSjhx5QmQKPsbbrkjzF4bh9290MpUhiIRj7e2AEDykYAKWDOWo+kj5ecVsDir3Ry2WmmM3zmbGKe
t17buV3tPE6SEx/+K2eLNjw8+4w/EzIEsod5EgoxUWKuqllMc2nknfjS/svM6WV3D+QgnE2o8A3L
SESICvZ8/G/m4a6YBrCnGhIIDcBIRr2400HfF/5SZ/Zikiv6rW6kXEiLk6bKPJ7OpiL4hh1oCvc6
3UPt0zrbi2uih6b3lWh561U8g5e5ck8A8aMU4k06j2wGbr9htGEEJrXJdQPIZKyv5HTr4qoYHfyi
jneIitoCqQX2YjTugvRgVhYQIUc8j4a1dhkXzofKMv1CRk+/oLh2vgaMxucu/mRCJ+taSocK3Ebj
79CbfQTrstpbVa6saAOiPfTpCETynHWKWvAKpziz2QCCkRr+UWDuPCnnHeBxTE2G0mQX+fTkSkS0
M/G39dicrMqhHFox61hMBXDfMIJgAB2wC8X9NSD9hAsXI3D7Vq4FN4YulSVv0MJExm2k3JJdAWxc
3NkYmLES4hEa4IAJ+wTO4pPg3bVmkXim9dDb/fNqmZNEUeECZLrx2IqACWwZIMY2uE57RU4ZJjLr
iAT0nNAjejyklMtKCzEL8zSRLkexpe0i/dgh0e/Q8Dx8mFTkpid3lxk8aLToqNvoq5jixNGHF0Nj
VQc7FEP7Y+ZCnnDk1tkTdYArkvYeRqROjlnVczTxdq+GBcqB1ro+XeXaJpiC0sdRWXi1RJG8Rk+r
Lz975Z0fx+jvbqvaHTrOg8gtop46ZTMhE6sSdXmyGbL951eXf6UQM8vtrFTPzuabPf8T1/Wp5+85
nWcMSiLyht/rXHfHJQ9V0hpd1N7Au6if9Z0WC8FnN7ER4yefmXneHCtxqrXreW1nLG9Dg8S/Yead
xZ00VV7/BcJCRXn/6ivp8U8KT64mKLztfqiPlKOIMIS8gCZjW41jQUKBmmi+yWgFytYRndOlb1nt
9RSiezj6do7rBIezivT701IXFqGm/i9XlWSPSqlwaJNiys6fdCZyWKpbdESS9NxOFEQ8jivZsWIR
fxClPitUKOLkFUAKR0QM9kgs9H7XnApI3QBelpeKS5xPCqSfvBOD64KKSpLr/1oY2BqlGHBE9MRC
gFyBj9ilEVOyZ8WFUr0uxyECIOvqHYBpJCyAh8tp+SMlvpwWN4xiOMvSNWPEDiSBZoQIhUZzS/Wk
KBkIvYcDIuA4szpkZ87j64ivhtAftPisR6DB2/mi/R+hseIls91/CDqu56e1McO1v6zrd7rqf8/H
znvKRrRtExhMrwbj0RYKtLYeYkjUUSSeDYYTJXtdDV5jIALOiK7JswAfFQCHjmjjYEjenJGB3t2O
KD+npLuCH04BBbcL8lWIVLW4fdbfXTfFJINybTyh06WvP1+44WLoTG3Ga9aZHvwd+pypizT3yKFE
r6/JacQIe+TnXTis3CPmieB1pqUnPyETrp+0rePUamNqv4k/A4+Ob7CHH65TeEnKXigm6YsLNm6M
lU6WsNH5oPqhn9Q3Ssa88VChMQcvWh8kiCqyFpZOfS8/ZqoCBFaoOT0LPWI/QVbpE3pp/iMuk8zr
/dln2+54CQf4BByIbG1oO4fSG5VQcQzmruGvGH6Aym582bgdZ0Uo5whKjZ7YVWOWkdTLTmt9/Gc3
9oykCc9OfkfxysrU85Kg3ZWDU5Q9Pt0I2ZzPAdhWcnxcOZsJ+SSGzkLv9XFs6hcnEu4JB3ixcMKA
ILgTeFgWNagmhD8nkPmhgXlJ2TQpyO2lhZnoSpsMj+qWGb6LJNjlBoD5z5/n5qm+KG58FbASXgpQ
ClDEh4KM0MXWJfS2p9rXNdb7r1SFqFNvop+SVGVvlfINLeO1UFg9C3OjSh7HvFmvwnuQwWDCRpgQ
BtYsx4vLFGimWVGafdXRR1b6PcozoHaC3qBxMXiZ+o5YPp8e7V8RoSyfJRDpKoQSFuxoP+HwWfTz
TPaEpkMThdwVDDDVhSYma+LePziw8KlmYrPTaRP4+VmpcEuGisj+uy2qfsM0iaJmj6PHcKY8yhND
d6joFtxhbQ4GtnBlmncdbDSshsN4sDjJZGRMc6KmijhRF140R1rE+MA4dLQS6stDLDDKJ2RGcFLK
1Y2kxCuPP6Z5YWuCRWP8KiEH+hnEJyTAHYx6egtfXKW/MjCWK0JDwK100rDtGpyIebAC3PRb1cc8
oOh0LaW8MxUwOcTAcPCEiv92urcS0CiVEnYl9KtXMyMpZdVrg2DWmoRhdyVF0I2NP0ZTrSy+1sxl
vPCTSm+ZsnORunmYxihfqBkUQZ+tOh6vcW5mMZ7VXpPz7M2liXEruythIb09azmlo/bVutiD3tQ2
+Q8zubpc3i8vg8vOHedPu+mKUxkJG6K2S48w5wFJ7M0ZF13dB2pNsCRoijuYEhVlD54l+PlSX0g0
00oY806j4j7tlce/LWbdGwNYLda3L+Wz+No4Wi5fu92h4GYMyJXL8BrdDAY3zMivm36QE8TAshTU
vifd7Y6dM/dlIbj9djMKRizb2sP1c0/iWFOZWqLS08lPoShCtqYE5g3/IK5vvWV+D5PlxPGK8dHN
XKw3raORfeV3q+qnIpbYhZwEdzWlRpykTpsgg9K7sxeV6SzQrHtPwS0K+wRiTb8uiRuZj4h71fMh
AY2gAGOChSXO/yz6eFoQMX+7esq6/3S4NvjLY0lEkxVRJCH4JGIsMDDY7uabwrcuyRgd3m1tD0yz
svmRgg459gRK9Hs/WWWy+duiRAR3rYL3GWH+/vCKz2hCAwXBXLgq496hTLH6RKqceSgOvwtaggeP
NkdAKcKYhjsFrbb8xaC+o4xvZg/QxwP7klj6Og3mw2X6HVGysSvfMMxwzKaPw+zwWXbPcKXceCtD
7M5YtagWok8FrYJS6ZxorS45G2Qxbf5JQ9zyfIire665tL3le2qkhPPJJ2pqH4er5CY6Fy017IVb
D4HabJVcST2fhKv+MGUZ2zwd0xOhwguikUaEUB0/uOFEaN3gsHuQGlwjrRYGyZYcKfq/DqwF4ZRr
CPjoGWGwA4dc50PCSQCbfXklDP5Rxvc29eFI0kJKmLruYSalxyIDWfppNfQeIgx+YtzTz5g3g60m
hKY3FJRWp0w1sM2h6tZG6vnOInbjPaIrops3JuixcAFXgrwUGzYbv/7W557GCC3N3V7QyeaWka7M
4l7jpNdLmhY1tE8ogriwpfwSuJYVlJ+dVdWbuQxTxtTipuEfY0EWKHQAFNV6/NPAcEnY9fmSy5v7
hcupIiQK6RwMbephYnviYoF/2a7rceT78dtioG+f7PXDAS73Af6Of1goyWMoP2YktQVqmr5eOzLK
A4QP+gNA2LZStyg/lTRL6P4Dwc5IrKI+1/deQsZt0xblckAqFJMx4o3P+axmiccrdyQS2HcVPj87
smnQ9ZmpNmL/jjUXnrkWVSmpLrYeJ+fb9gjP+sEhsHR9y5xxTAuBnmwNNysUbtjen82G6UMj3+Ek
b3jMU2xqX2ijUiEpnnNyBPd4/jw5TrGYiOCftT163jrw9Eo4+/QUb4rsn4f5FMkX6udsdtkkg5Pc
G+ttxtV8UdxcLtfLV2MNvv6IRyfEMYhPGgzdDWCx7HJCNzijtndd2cPqgvZL+ho5bDywzXXUM+zO
cLT491buZI3sSlrslZG2UEZlC4sSRD8zdeCKLjNm09DELkgYmuRTQ/XTo9IVirIR/Ev3ThM4Kbfe
iTso8EZEgsGPrgCEFN8OsJ/cjgi/4Cd73mwVHFZAAtOyOoKx0FHu0kPXJcbdnIs2ESMfxKsph/FX
E6pip3Oj0RsUKs1WoK9S+UdkPzQlNZ1tlJ0tf4pTjs+IqrknTK3SLPJLs+rUddfjMEpiNEXyueLG
8BI/c+3hq3SqT7rAqJ7Rst1a6FqUA4pqNPFI2VwRtqJ/OzcK0GeadreA1rZtQmPcgXgYRwcayS/K
JZVgkTN32x3yHwr7BA2BQ0A6V7rhzixSM/5rAJhjKF7L/qB8kB0ry5fBU3RHb11nVVvurrpe8Odz
Y1HAcM4/LNPsL5W0Cq7/eC1O7IXaXeNSvRIm5GLGj4H7jysntedJTzFXNmZnT5Np+Yb7QmcSUOTR
up6MvwCKRwEIlSas0s4XbXfG26V4ab3ccIgn+HSmSastg3MTkKMk07QmzTyPc1ikD/ICQvCzGdZe
iZjJU8VwZ9QHB+P4ZdgabYtvDdlz80r9JsRj9PN79xXquWl5FrVkZb5esHYFP2WHP5AuLZCULhpm
HXy1EodN+HderoNXCJemel+cpmiqdoI73LAWWLp3Bsa8baASydOvFYC2UImx4CXDS+mnST3bestn
MV4ojiH7Lqlo5WpdXFauKucuqLPNb+SBYisOdfaT6n9gaoUQUZUxDgL0RlXkwe+zKTOugnkAfjSc
9x6JKR/6h0HqGs9cFUrM4b1Kir6u/d9/ptJqkyOLS65p5FTRJNJq7AbMW8YQ/TmIqfmqAeU2yB4b
i+7+9sXtaT9dAUv5beBr4bh5d1J4PBJer0BXvxm59rEEcoGg+7+nmc23WcXDRgJcFemKZ2FDy5AA
VtEu5AOeojCrs1vV6j2sUW0qm7jQKlw/jWeIsCJNo8cMcxp+fdXi7FRQyWaXxEKO1qUi4gqEzI7F
zGSr1xzpklhC4ykueULL1Zke1nn5m8mvuNHGyXNTok8oR+UHyaoc4umwidsz5ukDXfA6TFqcw1Ye
y53fcy6iybQizBJpn8NIvi2WtATm3606IehnEkwg1Ja4MJ5SrKUdII5XBDgIIMoNovVxUfvoaIBw
dYw6iDUozZYOTb0rL74uZ9PJ3lW2N2HuPKjt3oVer27an/kOHcsGeQk32N/ehm0IhGz+Ku0MAfsr
FaR8fap4+V4jXIFlbtjLoQKQ2+tJCzrhQzbp1kpbsayLWj27Nltkz1xOC6Ez6HiFbHpDForn3RWK
nVv5d70ajA48WtHynVeWYARxuUMfR9Hoxo5iDgvngmwiZhBYZMRJjMyHf1fn6fi4E/Ug0uqquyE7
1NSnLAcxVCgVXn55hK4AdPzu9XlmIAVwd33vhLsTMvlE+vTZk9/sWgSWwMf10k5ECaa0y/sf1Jq3
hzsjyZxyHQRYZ2ssC/kWB/syqdsY0lGo69uCStwMZ1ZEt2eG+ohFprIP52298Z5Lfb1Nhpbjm+rQ
2T+nOjEUKvN+G9NxM1Ts9q6OSNQ/JfvuwSZBngHV8ekMayD1uWVKjswg5niDnOgBX0u+VptMriru
EJRSW4pJJ5MJqsAJmm2UyZjU3m66/jBZw301H6c+ey716grn/Y1bkURJndXksuayjEIO1+4j6LyP
zM9/XvYDujuRu+QHTZA5ER/SN5TabrEX77tOSn0F9WRUFyzzQkpsOKIOPI/G4eVZdKiVUajPHQh1
PxKndostPGe1s85GmkJf8Gjxz5I2Wx0kbWXDIOR/a51wbtKDLLXnO2eQBuxDQ/o0G+0a8QLpL/Ef
eBh6UrC2bXuncDYfdFUKvguO4ZSqC6AsvP/bbis5Z12Vr1WhmfPk7lnntbkrtkJSOX0p2wdc3U/v
/PxCTmMfSWpyVtj0IF+CIhwII/tOKDhn7P0KyRUUjcEYjl3PMk7+iKmUqNLTiHWGijinYFPpSQNI
FpHHUviwnte3I3Oh1Qat0ohMJ1kGqnzDExs3GCG0Oa/RyjslpRXbYUBzhX5RpII12MuvC0fMuwNl
f8GGc8PL7yuDpwaF+k5j+9zcSUbuhsGgTSNuhXlEfKyK5pGDJGfHqGC60wgxEcArXnDnNq+FRXLE
3lgzZht2GkiMqcl3fKBK989WpPdr4Hr2+YOLSS65nUUdjroNatQEg/NTLRL7bvSpIN477A8NeaPy
G4bi5HbBlvvPaZzMrLht47chhZeZycDVBwBE7kid+U58BBX+R8ElJSHpx3Gptt6VKIXq6Wf5hdEr
eYcE43+PcO53W7sq8Lic3SWqA1RXRC/lXzSnL0pDC0Nb3x2z+ayWrkT9PgVx2iV5wZxt/5WbmGV8
sHiqQw9EUDXIEDponGH3JyC/HSFQCHRqGxVJcJ3IXIrsF5n4ooN5ZBS0q5XXGukixfYKFdxWE3Ym
fyQCOJD4bKULsyHy4PCNhexJs7FO/SqB1tiOJuaZR92IzTUyIHV7jENi8tz9PiXRSj5zHOT1mwTl
VyyMkI0QHa7p7jjBncGAPB7Wv1fEZ+6WA71wKZb79DxH73q5A11xriiWtfflODez+jllzLItxOn+
+3PKQqVkKFfeEkMRMZ4TPY5wWiGX1U1qj9Cgc/MKdtkFJrkq4ws2lG6NBKsEmxy0oBXnall9hxaU
rBepz8/bd9UxVD8Ve9R42RETiIUTQLqHiZkMbNoIoUktzh9RjuTW26FPIWLH9Zw+2vTjHnd0ac6/
LXCWs/cW+2iT8lEnuIDeaoUjGBTu7/OaodeKjM1ey6ylu7MLZNvfec4zH7he9C43lpaTeyYjSOmT
i5RKowadJRnFtZso51aHNfuoSPoNjKzjSELNw2C5e85Di3GqJvE/j5O0fIhBRBsisQA37qtQc+pw
V+BM9Xs0k/JdQgfau88IF2pVyQWEj1rLsHHjE1idC87I6G2vJSY+GBA3EF3WKNOfz6YYOxr7OBbM
expiPUsjbuFcD2QavWEliRuvYpTU5SekWz1e9X/ioMjG2kt13SmyK1Zd6GXFTT9HkPmjQz2tSqxG
gL+6xWslNGt9QsA/kF23Ojl5tylchbVKbkec8C/biSnkReH6SLbUflS9MPXxrArvlWMMfTQxFTpr
V3ddr9T4BjDMKWWCK7L06qh1T47dmTJlbdPzD1W+6Qp6sJ1JGB7ki9inPJmKz4bcSvkO96RRlAR3
2V56WJyNPAz1FCFfEch9kN5oXXc/NDD2ojVMDkkN1eiqOAUrXCKsKJTXvvb1DPRGWhwWlpxIfH7h
e20Q6rl+2JSgttoQcnlhP8UhhsiPsFm6NQNWUCzSBtwKymcvvrASun2MbJhHAbQCDjp1rRqN3sov
KU+T2ixDhrZtfA3FBv+fJfAeMZDDNj1EhwJ/vRQkOv7K1rHfBfV4Tu4GQCxMmHp7CD1wBCZcl0aW
JSoJrojBd7U6M/VBmHhDlIzecEZxlk30VYdq6qTAhl9f5jgab/uN9b4pcLo4qbsCldn8GLDq77wm
4+xvr+8MAfZVq1nQiRitev5bcWbrGzQHX9qDPOe12I8Hguq7XJicNDRPTFDx3yVydLkh68uY/YS5
M5MfNrIJvxvI4xJvSyqHTSharD4n+RdUufZwmbuK5NeS6f3KrJ6wBEk2nBr92uQTUafPVbJx8yZj
5psmi6lVZIyDMfx7hCHgIxHEGqdislhL/Tq0mVGyFOcLRDJ+FjuvaLs3QI+T3aTROtdwQcbn+Yp9
QCeKHsL5lyNYvbM+TxSFuCEbbcaGtskoeZV+2zgVjoY8gWIhCOaSbFQnzNY1W+4TeugQpboXhAY5
rnniRuhnWPA286X89MoNcW4Lr3x57k6USEqqWNz8+/RnZ2LzLsJ54FvlFUhY2/6mkQTo1dpidwQY
lYYGKEs+RiOQSOLyFPXJXOOuDRbDRfXcrqVXPyukJ7oONG5/vSRxHxa9e1JsH2JxvXoeqSyqttsP
4619zGaHzSnlb05iRvBe09gzWcWFHqHDUGBk3zn3TGssPdQZx0hePNKoUo81OYFch1xAD6Hz07VV
vHhCrXY8mTUC1LpdGhyMHI6UNS+cx11o9zbC8dUyM8ehEb3Jna2wxhsoGIY/Ud+N7huALLSFt/3G
zvXuG8L045mWXrfAusMM4ctTBaDPEaZgDhkdbkAYa0ItBlkEXuhD6QfAgXBZhP7gQEZkw/nS32Wu
ywsH1C5ck7De5k2ERH/90G8KClKqn7J044u4nwZGN2RZWeGkAg6w7Hl6kRS2wdaptZtbatSHdz7A
O9KjzuK13eNgMz8j2mfHxROfQhgFc6qbypmY2djKvdQN6icOSPo4jDyxtD+L5XAVCKVwGPRcCmZj
yR7L4TXqjKmdHpwL4lPt4kwDzX/jOaKCPAuz5w46LlQ7UgQsz4vY1MdFr81rVQZYzQPauzJufh9n
XOXpysDnauKtV1X7IaaQpR3wVCE8tU1D6yYccw67viw7pjwpJCd48nJ/g940HmPUQ+CYjkUqqIFR
hOF7nkR+gAGr/oYmU+rlLWEGVPVTnVMCmCJZEtPfliv7ZOhQnHgUT/x03Ym/IKJ/no76RdK095Eb
6k0mY2wL+MEE8lXHOweL9txTaar9/t5KT7cuUIj0sh7BrVVgPxJMXXopytLU6kFZTSfbFKVNJjmm
zDzR/iFkIHpTmNC+h8p9YRUOnVKx/BwDBR7sIN5yuh7r7dT1kWp/lVFwEnP6Zmf0bLgASSurM+4Z
eGdaeKhDh1ftwqnlBRjzJyOBHbItwWBGZkxYT6scyJb/wPxhXYZu7Qs/W0/dhmSXnYl+BO7C+JwD
qlnMH2jXnDxdJt8WHVEE7nJQRAP8KoWUR3ycYhYk20/hLzA2zlfptdswwo1TaUmCObiaaqy+voDu
ZZGuR4OyVa1vluLfaCaf3XQhVm2KPMv+OfPRSNG3vucNj54WWNe/xMGj1qlbvhBK93LWUeKgY3j9
HiB4KuHl9MUZeCAz5Ocgkt1aKUq4yiMV9Qv9U3xWBuj3V0n41/RGUvsH4DL8gVW2xlk48W9kNvdc
flFFcej2uNALaJkMnwntFmPhBdu8yP0rQ7T7L4/tCEZp7TnFlaFh0pENtgn9eU4KYH2yj7+kjgtH
36/f3p/KLI+4sGkroWuTuYe31hNvWD3JxR+cmYdfn5W2s29qD+7W4EwyeMGVqKYEw2ysqTcUYrW4
2jHpm9XzLNhcGqVvgFG4U3v479hQfxoedFToQteUfL8/nrzQz/4lXB5visOjB0F+Zbq5KhS0DkhD
SWwCn4jtEzdJcTQPZ10ptGfk6KSNSltOqQijQcusgMTBy6NHQgDNiu5Z5DzqXepxudm050BXWY/u
nwW6tNj4iA5ZwHTqEQqHMtFAAos7QQYkLgfVpKvrtCsFwAlyWR6ESnfstrqTXjSSQCktQhtAdZab
n0sOvzuKPtjowzk87uZdy4UUJ3bjMigDIFhMwz33n2XfIjMDa6cF5o6feXm2lys1G4AjMHr19Aoc
Juq1ridTEbKMuTZ4BJs4l2l4H9SW2o0nirLS2wgKvfoNuX3fe+MV+MAj/GFMB+yYqkUOkFQbDuB+
ihym77QaUDqPfxuC8N9SL0+cfRgM/Se6ZugjwkMo+XnWUUI96C5G8UY6fJ12zgdRYcXV1ARPt5WO
BrW92I5F9YMyQ9VAylxMg1mgngVfIPp51NChDvDQp8MNNwSHIt5fC+2iag9J4SQRJb0QtloeL4F2
r0NC3baM5Huy35zSQx/WfCdmKbu7XL6GDjLaMTTCfdni6YA+3u35AjMRuj85Q3o1/lPQRU8NSXjq
ljzepXYX/m/KidpXX9CLR33q8rBzqEpY+p92D2yKutLBY2sldYSJYPos1VuqG4uj12PxpL37oW6T
9/RxBfwE/DWNIewZJdMwRg6GQHrvhDDIMdN/gG4Bbu0p0ZDPi4NdThxIEztaeeI+hkAUnM1+TMoW
FUI/ViE3mPZ+OCmiG6Z2xc5ZULz/6h96iwRIskibMFxb4OGEzmh/IDm7W8ESVXajNhzkV7rCmMDK
mUYhtRODmZaANtl2CfVzzixNBBp03rgRh6R8pY9khTy/G7mzyAue5CHy1K1qvTROcPnIbfj9HrbU
FIGuNAH3g0aV44QZg13smOCFBG5ci5HVU5Ift/tq2j3VgF5/DR/jShOa9OVigM1UyKY41QiAezub
BuybLh4I6JRNy3s4c0uPzP6Xj9HgUXvJ99Fv6f8YIpvP+kTUsxIMiww/SWtwwPfMXioXJ5WdU68e
NkXyjpfS6mWXEpEAMlftHafkMLTEimHOs9lGgoZcAvhWoYrTgmQLeE8D1BBzNqItr/4K7PkoTSk1
hIQmyLXvmfMV3ZWr9sVQpgoVF8YJ8r+61yaUu1boWcYRxu0JFtJDYrpLDF6PBhYKpW1guraOjOIP
vGgfqDaPDCHvcamXATSLgLJT1/pORPGF4A9ah0Wdb6WZELYQItyQTjr9wGj8iHiv67pYmiRrWx6F
RKfrAvtkBa61A6gH3j3Udug/88OFkES/ZvYMfymCjvll6WP3JG1fT4KcFzhu22z98qud+395XNCX
KRMZpX6vu3+C6vxOH0SMUy7Uj8nH7hstLeucCXZlGL1JBQK7qng2eJtYLbA+C1O0m7zWfaDCAIoT
K1YLnkpvy+NAhpg7mqBOvejtLDVwPHMsGsid6gY/0HH8pdv0sm6YZ9s5gKGfnI4LVtPRg/ChKh13
h/sH0+xQZLPjjjLgAZtg9A65CIpD2G3yTQJyeSUCMbz1PI4PZ7fq9siiY1OV9jmDU7SIi10dbqBx
9UUXQqNHsUArGu+EDkkKVHxa1TkrznAMzDnZEybtKjSVUlDwx6knnsU442WQJNFTH2zIXBcjoc2x
R94+BP5BkD2vLJzRTddnKWUdFE/ewUuq9dzTykvxXkS2cjQNCpWHrsMom0VCAoc7FH6/pFT3Dbow
n5pfy8vRbXvBn7olqHeZ+HWgFbe2NUWnMFSuu/uK64WIpkkv7zVGOMs8GyGPZ73q2RlE3yvVV+aG
qIcKCmakTwXeAgzOxhmpsTAXN3R/dSPGvLewkTI13KS9ZJzW3CwYR5AEdxXqgQ7IUeK+NwdZ/5RT
poRF72QOCrJkRmoD365w8kmrPwTgCVSkOCdeFI5MoDaX8uysMxtep5rK3thlaLkAfeQ5V+qyPukj
AISkYVW7xWhKBbJ7Izq3Oxbydy9il3mjvzsjWPiDVZxVVaUUZDmzspqro/lwehF/QhzkZmmearQI
WT0wKkHMn2AqxnXN+POQO3eoUcXB8OhVp3BepeiNw1kTVm+126xhqyKhwCTQRpeewvOxUikydagg
pkwVPbFIRWOrcZa9EMNWVhAorsVdpmwa2USRPppbcnch2wgcF2UXmosXon+n8pnfz4R5XYYu2F3M
/Oc8EpSi1I169/Q9ab5EYjRRqkKIWl7M6ToL8RAyPCpV52+Us10uS9TTDXI9ZCqqHCFXV+aKJuvd
C31ufwVN131wW2MnvuvzPlV7knKcTC7jJUyJpnCOQeMRYABKfUPjSUqn01AmafZh2GREvVfbi10P
NH6GK1wsBA9o02SrJZ4/LIHWsJ4PtORDPcvZL6x0S9QJKW7qpRBLY5qCTEWI/n/j2I8e+02ocmPB
YmbOFyO0DEWgjr1rEzbQm1GXDk+UBucUuV+TmT//tBamUiMGt4amaBk07h5bZP93qqh5VMyvUtxw
Q0ba8OPyNMkVsIAw4GoIrDkMzVyy4HfsAygYKat4umtniAL8/K0IIX5PywpduF4xKo5Uj+gmGCCH
sePrZaRpUQjXfIwWZKh32Tx3Vq5QKibUcWn0k+rqusRgkSi/FwhG68ZC2R2fpZXmZ3Lu1XZWcMVY
7oDF4y7g1gz3JOL7kFUVQ3cFe3VV5lfEOFru83isVIirAKnolT2H7TQyjefrpJhGicDsnvwHOiRa
Ao4gfu+PjRqT5ZXGHRuVeuWCzdhkW6vP0Y+SsXbYYg2YT1/jlp9Rr4E9tsEb+D6JqJQlIxFZCO/u
+uPy11Q7Sol5iuui0rf3FPdhvsnvEh0kZfkARTGEXvSofu1Ic3xQz0kOohyralENGFuAgyaP0lTn
57K6biKG1MMUT/uQ1mEqBFEqEqgCPSggl1MWuwlividr0AIXiNn4mQ6ZBxm+g/73XJAMLEqebqvK
5exkFs4Lgb/OdoqYFxSyZDKNyjO/Kb8csRPAA9r3y6XWu4HgA18lcFfSBDvra/V0GjlOBmESSNYX
9RUUIyATShZStniYh4pzWOz3OTBBXhESq9feE7hIxGym9Ou+RCGoBz1udYQ0mWIxvlEtdcMjrhpk
84itMMx3wLunF0cC7EkI92l8LhSf8NK9lXeNuGRDuv2UhcTzJygOAmi7E3H25rymydDry+wHaWzH
eKENPaN7p6xgelLZIbJzLJT+llcZq+m6e82Lw1mRgm+KWJ4Zq3UIDRpDgCUsbClPArz92K5osV6i
wjBEH2erEGW2HgtV+8xoy03I4BGRx9bLjddXo/VHH1p4sNdYW3ditKdMRFBNElcA9qzQDZrQh/IT
+Cde5yH1/Ia9KzXu5Xfl5gLMl5eKC5OvngQVg8bzsSwYQY2c+Z7jr/x4KzKnlQUo07xL8QsbRV/V
J2DI63VnIxfn0GxYpsRypcDAXBLt2TkkTUImlqAUgTBJF8fxIOlCD+lE6tcYWG+GzYliHlJg6aaM
MbO+OGe+68iIUDafgEGJyJSPshHw1ytEje1NNUfjj5RoldOcJricTTXKbHrfGpUlQHYjVmvEup2j
hlKRNLeI9YI+5Dk93JohtPltFXLMs37i6T1WODd/XYaGfqb0VWi2+34OkqC8lBKweu5o0fV5OCCO
9sWZkqRylW2cesXJmE5RXYlqMC7Uolkx9u8fQPLhaCMvpHz5LhgnQFx5g9kxXupS+sdL5yi+gnja
qsnIyP/wzf1mTWW+mD1o6q9J0UVR3/hKgkNXQ/XXFGx9e8lXAYIczPvOQniS5o1SkNg+XAwuY9um
mnJycq2hH12qmdVhAxb7hhAppp0fks/957av+WHBx4FAGyJIQQdAH77OkKmnDmfQ6YHztqkcON6K
/4NhFNIzWSCTZAMOBC8kkWNH6gkmJw6sOCjZ3ldz37ZMvrnxm2BYSIP5WslZsw+OO+v79HkrlGzT
mFDQX7Ff8zcLE8IPtAiU/ozL6C2H5gCkHvmtvH/Hl7HofzmezT81grA0H1gPFaGzxGfjjHjHUtP3
YU96I+QMOLTDQ/+Dfsx4F4ur2xY6z0HtOSSFBxglhlib+SCqB5xYNVOo4r9eT9gkxm2n3ByqcBJ5
xJ+T7mhEj22Us55tCYuDwXf9isz5LWcRNbO8w0XyOFjuwaKab2+8s4tiP4XPKutMEKkc8f+yeSf+
A0iRC2ym66AiLhk5LdWbRh8Q4V9gX+oAMN5+PWMijcb9NrRBOgF1VtL6mxqzum+GdHeJ4sdjnH6I
lOkcxyOykpLkmqdzWlTJPoUpTlXGtzLrUUhVN1i1oh51Zsu3/SBx0rabnEpaHKCPLfUUirpDXHsj
MNWr+F2zELqt4nnAENKflgwhxsjOBzOhKKRw5I6QEFCLJldz1UvtkVXj6s9gBRsx+zZTN2f6kl7G
frxs1iwOl6E717j94Uq0+XIrn138yCZXC6cQBHiY+cG+i46Ioqg81+0edAzqkTaYWUsfkV6+47NJ
oxp62bckyB1OJz6TreavhBv4Eib7SDBwQZItpn9U24k76LZhd1GXWMCwLoNMUspyMbPx0H8UPGzi
9pT4TE1efFlvnLyVhGp46tZtJsZBD8rj6Qdk0VddYCY8o5KHbmltyOZFy7T0BYlLjckBi0An3VUX
YTp1GH4kbtpZIyhdsckL12NrUSoTc5zWEtsnmoDKQuiJtLnPDyMKuCu3Q7xCm+7VZZbiVFUHxF/s
F79/uuHwXTVG0MBMzTSHhS0oMOcxgIH7N32geyvRXOaR0Q5Nku2iOhPxjrygpZBEOkiGt9OdTTI/
oGpLwKUc9CLtB4ZZdEOhb5QHn4jhZtdT5Qy8+rh2PB835JWTgsbTGW4HbH9lgiNPOPzk+c9R0PpU
NkA405HmAeqn2cJchV63iusmmtnIeVoXRaET6ovUdbDXKI8a+4Urxm8M/Ff3j8x42u20t31oAG2h
9yScjFAU3gUxx2buupiAzNePdvr+UzEcJTfeA4ewn3xQtB8BFPCns1u0M5nI24rsGjoJKFi9lmXr
ajHbapgHyh5A+qL6Ow2CTIxp8OLNNh28o25HjhT533XxTruzliRpRFlUpclMzHUXg82gnEnDh1H8
K3mtWijAyv8VXpojv6x5sOgDpGRYDSzrmJCQr2L3NjxRM43EJl90BD9cH4ZxFgoCp2FAQ45sbDEO
eeRdfXW5zcxf/M4LQA1nQI96E6RLAucEyQvTdG6hhQfxkWTm81cvXBczvECZj2z6NRUTceGlg3YD
Fklh6/WdL4kHFVxXOsgF/KufCdHQSIk57YFJ2zRGyilpKUvGEILQxlS2KaTJfaT/FLJ3Q1IOxJWI
ytFCDH53xd8WiRw7gkAiDUV6ZfHPNdE7qcsfU6QdphbUkgvQzDyOf91mbymTywmo7fStpkqML6jy
ylUe2zb3v8aaJq2rTeHjVLT3jLVSu4RCSF8FQvvo9hyESGok7+HrDK/sFZxD2LEnYw72kv+4o29F
LGWyygJ9appWUWX5bw1/I7xDf2zUB8pDiWpO16HvT/6zjeXjVeDNzGnboMbHb63ZmA6UPhSfk+CB
7nYokSZoOaBLBsaAFV/FOuUuDBUtPikxJkDG7e9RQqqUqeEpyJIqcdaDu0KiMS0WhycRugzk2SVm
rvdi8L13n0GOhc63UyMH/oJmbpLekHGHh9WlsDA4RsWQPjsGXWrSrqA9kkZGtA3nL91ALkfkvdrS
nUe/ZWqT3MpmqL7p6RNZXUqoBqcpqqElMRU464QPvWz85s9H13alRWyBb56uBiIELdldvw5Zww7A
hN0vtRgnYOCelyHX7OCA3o3vytvTJ2Iys/8G8iJdxO05QaBEYbgXTT9HUY3W/w3yMC/bpVr34Fc6
wubbDUWCP+TmD0PbQQWVjz3NOHgDWABkHR9zRI+GnPe/+tQiVk0QxgXxB9F+JasuapZtLkPenJd3
B0b7yp4RD5nrgv7zi/mqV2To20Qt3g7xBKfwb7qRgt0PklMIPFGB/b4Kfm+f2KdWG3i8iFLoEVa+
r/g3QFGKc2AuaUJgMiJf2X7WEBLtT4QsoXdhEZ1JB0qnq1/roYZ76QZ2P6qhnXaE1O1FT2IPlK32
Jw55GWlcEarjQJSxzGninux9MZOEpJBx7F+hVgbLxq4cZQYYesCSuZRHng4ZVd7KUu71sGl/LW0w
susadllm6MQ0ZJIZZZit//7pYRPNT25h8hDadiDmbzNYAIH0y5GZWHwAMqs2XkWW9O3seoatd9Wu
uioPXjIZ0TB6f4p4M9smk0+L2SZVsYJ2Ae3r+dyj/mC7SPXyWKH3gmrVtq/ZgpIfNdMZakQnaVkl
TxR/DxbP9Y2Knp5Nh62cPWhLWN8FMrIxns96ECjK+9KU7XlDuCpbGVA9ClR0pp5KTQtUnhq9f3Xc
eXH1mJv0d5Lp+HsFZPtoQHHAOWb0TXGYPxxDXfXXfrhxuIlxMpXpDZu5QFs/fG9vXjEIEtV8O0v/
BCamHabHdLtWpYQsIHeV2Gb9Z5de2rMv1l/MXuTgDVfAN/coEkr0GUWsAPQJkq6bwSUINt+BDy1/
OtpOv1XAsrQTRuQLTRqBITI+HQnu5vTBZZW3Dsh+jR4bF7DquXfWqDRTe95VhyBPnyQtJvusjAKw
EdV7Xd1j5qPVFiMCy9Dr2d1L/lLyW6NxJpLX68384DUPTFyYkxQzx3pXQdc+Zz0MU2U2U0cJk7io
0vX94uUXy1ZUqG2yCZvyf6KKhPpfdkJPAj7He0HlGnnIqF/Q1+NMXuWVDz8qBFDpIuf0Bgjl5AFA
Am/2CxU/iLtx6SSNKaVHV+giX622jewELYbm53yOnEFcGSebiDpVLTkEVYSzMJ/xTnl5TNfZRlqc
FTwJmkdqrb+Hzcjl15zSZyGygkZiadkyWhxRjceN3NDI0+3F1eyhdpO44Yiqq4xrUMQd46t6m3pw
tjMfsva7C4fOT0DBqH5YmrWjeJPzSK5Ppfw5HeE4o5Otr0oNKL4ERtouTcLgLGLlByGdJOfOr0Db
ccgX2XpWE7ISQgh+7QcOCLTcA8/VXGtZ6QDWwraE7MQVynWWGS5iH71NAW5sAic8VjuggQL1bWJH
XdRdTdxzXmHAlN+YCLuCajqs++eiG7OTr680BKXrfsIXurLY/LzPZl4HK/a/Ff4muirX2CtHeigR
NTbNzWGvvip1SFzwN9vxIq5bO4Fq8TwGbPp5Rthc7w3bSFQI/hXlUnbcveQOxmWpKVvlQBGpF742
MVUOSjOoBxfZNqkdtyp3yFMtJZSnMBSNKWk0DKUYkJuyWhErSAwUeSR4SyQ7cZJxhpk63VQF6yBq
nwy5V0iBtMgI0HYMxxNv4lPDQAJl9ob8NzQQAKglpbMex2Ddeoi5vqZw0w9VUgKQRpNk/UzuVs7P
5xXRUWoO7PzH+2/knsMtOfRyFWKaa9WnGqc3JjUUf6NY7dsmvZr0Vzu2u/PaT9e8XxUqDp9c+/y8
9mZ7dYrZQDhj0lff0dni02UqcF6/r9YPTaxic3Iv6/gJLKj2deFPOvD+H+KkGiGcVr0qvPiNUURg
PZT+bJ5TbUqvcDPlZ7lzg4/rlumjQqzJoDGo2Z8QPlYpoJnfgBs6w2XAi+9LymK/CFL2tsrYRhRq
OobSy0tDqTPSEdQEfADwejEmY8YOeu1OowSLM+DVX1Ny4oORHH00T2roLL1sN8y48fXItezYg71/
ds9Zm6XnG6i1OZnYEuDseegmtNjmhh7LF7bKBBv4vvCZAfEKNT4Kc4WAfxKE+qcpLeCzNlWoVsek
Kg1B44orK+tu1F+2LmlopnhiWEwGxqNG5FS65dmNYTUGq7MiQHvRsf1eL/GilsiS/2B99lkAlkSr
adJ7ZVR7qTMlLXCT8G+P0Fyfo5+e8jG0qTTpfXPLHnyK1i2Uua3MKQ+vOXUajgZX27brVCAMV9zJ
0BV3QZh6inKu6yVPgn6R3e/fUYGhF4sjak4u8wTSdEJPxFPnLRx71wzC5ciKjoYoNB7EIjJdYMH6
qd7TwgOe/NPLesRtrOoJwxqNK78dZKRzzpycE+8MfDimoo9qYWLp1s9t6x9KrDgBiWDJVLXgGOEU
0nYFyqEI6icx/5bGQ6ussW1Yz41k+r0pk619Nd9x9tvfJdVwdWM/2q8NKuFeTk/02/+WJ6CCde36
ZOOHEVqEp7J0CWPSvHt97oYvOMge7Moy2XwzpxLjgd5Lea+NwLKZ40iP7pzwmyBa7VDdQKYfGmYj
Zb37nf3VyDpIF8Mkw5nsOFl0IVVFQLeW9joa72aDgYNQBSa69TrxXhaQbJaPqdqmT1pp4JxnKAq4
U8JFTPoqhE92MyorLFiPdp55L3XUV7F9t7emrjKo1Xninj003t5tUd8TGIc8t78ubqvhNEjJkp42
L1xFu73+04/Z8lIs3Pkk9BWFjvq4xuDmH3cc78AlrmUt6Bb+9UopoptM/jbdD64ifKETLYFwWG3a
UCIfbsCyBdJEXxVXyC5Df09Cr09Ow+PYCSQP8hX0MtlEzDEDgOwXsi4kjAuJh6T0hahzKiiRuLcB
5JorM5iKiBl5PoNoOtz9YhbkSi+cfJY2OsFeyugI72I+rlBhpvzGRgJeeMscU8OdeMoSYpyvkerR
Wnko90nS1nDPJFaylAFt22i/qhrUN4hr5/FiRfKt9RT8Q9wYBxQJ0vs+ZfnW2OLvspoNKNhrvHpn
R7/lP6x0+96b7EYN5FnPKJUX4kwBYuO2jY5pzGah4ljqhtvRxhrFsuBRgBD7Gh/OQ8u4J0RGIJdj
ajCk6bFE2kLxGY+TkYOvi2qpzyRfJUxD5BJ0/tYtqX5ovEMCSoRZBdWGHFUb4UPB929bY1oU7xmZ
pcBxotLkOwpJF8QGaMQzESPGTVaxC1J2lg3jBodqr8eV+FVrQ76ahUePkq58XHLVjtGkWHZ2/EIZ
dxx+JGoJ7ijqs6bn55NEo+5mrSystm5nR3DARqcVciTTSZBu06fkCV5o+tg0XCeEmWIlTkh1VFon
XB1XmSc1+XgWTZgiR/Q+kCtOXsPGg3UPe15RJ18ELdmKDAN8D2MeAZhD5fvgIaNjtPgrNXKYAunD
e1OO0qrZ77k+4FnmhO3iQ890buanVC9naRxt+I5cGaEmMkY8Hvheo4bbe5wqQTU/5kImCW/ISJ2s
F/poiAcAR9OMYeltD5YxxZENYXR/ocSgNTEADBwWHU7RpmkSjl062D0xqDLmKt9yhRhfB8S9c85B
jQIfITZp77uvhSEeBbRLWrtpwNO4m2qe99nYlcPm246x/GCLnwEGT/Rp6TRasq97OmRSCKhZ44q8
12XYJfJIUQwJCqQNvXYJ0aDEWSYwM1akyzWpl058ErgLj0IZM3olQoFK3j+jvjB58fbAfNDfzMUW
EBR+rz2eJsMBDS2VahF36KZYafXcREK3CgZqUHBywpU371xlgRlmpemFeMiOK6Xbj+rcMM3D/Ny4
U968PEBMKiRjCOBpeRnWTw7OGFYvDU1VC4w6FWUBF+UDX/9Ud393G0+bYVWYZsBFoVVpHCq0iMl7
tNSoQqwYQgyboF4DP4/a7SBOdM+hygUQs8ppsYSz/RAdvu8Fl6dvQmfcUnbYKspsOOvlMoEV0zpf
r9iHWrCykYtFoMmYz+a2I1vCKaQA6UawUhA1ZaQFDzgFctK/g+7Klzamyf6znmS06CnbpruHil3l
HbF1+ifG6GkrFuyZdShJIYhEXeFjrojCoDcaQkov2DEGb3vwOnNOuEL8bRZQvSNCKyihIqSYOvLd
gahxu/dydRi3KgbLYiVg5XNHdfQd7O1ySuEjER/85XCt6jeSHuqghRtzzqt5HgQ0HOhaDe3kFZ4Q
1iGBZeBVUTnAD1ueeMjzKSms24NlszmhyRM30P1OKrlFc1IEGJ33N3pox4V/EOz54b6pqmaD3F3r
8Y7TO7HTNZM4bzy9NlHtlS0pj8CvHGrDUAP9xUpKFreUqFN/HzWabDttEeyjNRuEIAyvIUqSg7A0
KHoMpC9GwUKvgVuJ5w9xcUi/oBGTDi8lZ8Bx75Kzk2cSghsxyG6DUZ0oT7CzSZ/Kl7jQRGO7rw0q
ggoy4ADSw5ZRuC5IPw2NSNegya6sTRZ0XTU6H8pEL6+5oYNxtKKgO05nPXIj7WQIXqCAE/feeTXj
ky/q5gFEMj/K+Q8fcwwRjymVxk2wcwZ8eW/6Z5L7I9hq465hbHMM4HBhUVJ1+lECUC9v4tvrXpRL
wXHfZEKGuNkpV/2201bTFb78QZMwyMnu4kr+3g4qyRcQnwLhFo/7e/mdKwYSMHvfcMsRttrOlvGa
Rc+jIOkeVI7z4lDtT6Y5nHuBgic7/bGrvS5kF1jmehS8rF8Q0mUhyztEgIbX9oDTXdjJxdO/6iSO
ahSGoPNqiWrLjMmp8VNwz+84IPqheDqNYY2JRjxj7rXIN69zhTxO/wJfZx6ADUQukJk3VLdeROg7
DaMzP1CCbDebSi3qfGs1fP7pdvVWikqYEsibEUdxygnca0D/C5tPcpohAHovnDn5qM/Z3JYKn9sJ
kTcN5fDK8WDXYu+2yIAvQWplEolfyFDObpfitCGOTJZsEaxeRZPzhxHuzZOy0Pn/A+4gl32MrFhl
POyv/d9e0TmmFei5YkFH9kb58Cis4lVSibYtKZXucnRfrg00vx0x4WvGurzCrxaPawdkdj8SfSCn
rbC5jP9mt5VAos/Ps+yHjYJQtVCAgwfH4hJuo1OqYxvSnPR/H2H6DK1fBrowD60G+kiMaoHidHU1
ygQE1pIe50SwdwoP39/NJ+tXGc3VcKEbUHtQJMxWxFiiO7l7TVBzNKcHZqkNvcVPUTxOS7PocTHH
Ao6lLnj1QwSgPyeg1E/ENDNflyqEdfJDvo+1YS1YcxNIPxVETQmY4/30/Wonyuj3ThXTNrp7qDL0
7pmRJ7TcFI033urDtRaP6UrDB/TVQj12UKjT8uuosw05a/WC2Qg2Qz2IwRSxdYsg2YH7GqKIuVko
X3Y+pEX12hgMkMGK/n4I72RKr/de9EkbEPl8wYHvbQ+e7bMoWlreIWD7CLtFiXgg59p6jsALi4MX
8hY0UCzAsUBdatTbDlYviHwYVd8+z/9YHv5JpbKH56PiDOAl0DaKbcwvsfa0KeQ1cKGpEcbX9i+d
YnLL28jps+mk9H1ss4pi3WKcIn1zd/c+3unkjdQtx9R/wsMUD+N3hKnhN5VbLN7kUTnM0KwHxaWH
xt1b2sMEdly1DJlju7IAHb8vGngSQf3jQVoZFPNpZq3OjdfTeJmpcYtAMd1ZExDQvSkpWhHd1gG3
qbiXcRJSrbeQpjx1AXHXjZyxpH4t3tgrlvTYk34ABMOsnzhsKRBPwycLQ1yfKetJRSrTD1xteg4d
NfV13cj2O9DSzdJWn9u1bIeo+Y38+c9a16q2ksvKoMOOWc3U1FuZc3yYnksnPQedkIIqa2pal3/R
kHyRInIJYCsCGsVx6u/agOHtNMagfNVPE/mokv+jqCDAwFOkrhtlWoV8+KhXXD9WliIm89CThm0d
SW1wC5BNIQ+CCmK3joiewkyU9/+VbMBmUE+ePHuuc/1rXlwXh7zPgX0lJyjX1AvlAlTiPxMAJx2a
qn9U9wOs/JzsQX2EWCHbhUAOE6coKe/Ooqc9CQvXas9siLP8pALzaznvS4KbRKQ6ZziOj+S2Eiy9
r8vZ1oavDvLkOYeMVfVFy8rMe5Ai67RpJHGnEOO30y9d+7xDo6g2QUimrtDxd067eIbe37jdI1BI
Ju3toslVIlbE5fIEFY2N//hh8OjREjgTw8BGFNVNpmnxTaA3Bnp61bWrxTSx92v3Qr1Qg2CVoAhN
xB7L+u0vjjNGoPWIk6E5H6IVbXduu6w8KdUwo9lC80fFKXAgj+/lQ8NPxvOL66MIEpe02w7v59wi
dOGAt0h3JCJDyH5lYbi2aPrg/hEnjeuM3HwvFSTJEkQZ+0xjCIhs0dx6cuO3B89exvQdO5iP3fp+
MpquxFAtlBw5QPh6MWGDmveAhpLSn7W8RFOSvMIOJLUYRtAsSxFXjvzGr8S1plyvELWH3rtwgcYl
ULHunPKohnotubtxzxqpMQvBrJKtJxGA/FJGzuiNVVLuRJBUmpYPbCbdbab0QYw8AJj7X3MrXb3a
b1ziFpg3tPoJNa//oH7X/2oJsrYDie/jFAfceRHrsf+NqvFiyGwmvkmOPzVnVtZBGYTcpzhDJvJf
aboiJYcri5WuaHBlknvxTlDGG2tfRbyzSMGlGrU3HbKhOHoqsMYXYhZfzm2h2ByTvvRo62raVDXw
VKGAvfUGxXh/YkV8XdeIFjFvggI2ZvVAdjHhKkQ7EJKvfw2EmnMf0XJovZKryDBFgpFfg8//lMoc
ENzDbO5/CXICdPqnrxYcHkyGNR0LseAY/dDKDMRbz+c59WcXZx2tZWMJ0BO43xIbYlUxYY5xl6TR
8YRHSkEDLnu8uqtpTIi1S82IQPSroZWP/HpiTrCaaWc0iIEvpMlgFW5+jGJuDwjViETeM7QPwm8R
Uj4lLezt1f8FbVacf4W8IlF1A6CUXBOww4kC7XkjDKYD0ERs4J1VrvfSzaCtHUcMPipqaBB+Pqup
sduAAd690a0HNTIuvRzk9ibaRYtvZYbEiMUr8ZCBH7hS+m0XQdEakzuqr0PjvugGuA/IVtQc4QqJ
KBe1g7E+qvm7+v80aVdSK9526arly2+rrtXJQT2lrh5rCH9669d/pPmf/DJ7pMkXtAxIcED4Ih/S
1qNs6nsNJ6kDT6jGYCicIPyNyseEBEDCYlVtNYgxBx2bpkHI1K6VVJRuYlK693NSCgQl5j6dTO4z
Zbj5NSlPO6iZTmJaiPjLSxs+Y6No4jJugQGfkUJN/L7eyhPUKiiCsoEATY6tNvo1w3dd8XDDiNOy
o+X/pzkVPKc/FSUYwxIDxjcWQ2xx6NHH40QsGqAF+gqbJZ2UchftvrYQrwrXY7SAaDpV6iGc214z
F4lk/4nE2olIx32Z/KcqIFIu0Q/lDdRcZv2KO6uy5zYGrzntZsEaoUuOcWXIWYefDXyogidmfRSo
9+/n0OyOMtu1g/B7bYBC9G9bjbTf5L0au4l6bMilkndrZBLeI9YobkYy9+VZpMg/jU2PIe0oTJSZ
+CXGAo9bbTJNViOR43rUKZFUmx7z0zpW37Q2dbqZ/UcMJUnHJc6fZAHhz66xRpCyt9aM0ZHf354p
9+EC9MBX6dsKpdK3I904eQEvowRIbjJooQ+8uOW5U9i3QU2WOgKb6DZWfl1RGsyGb+tGgXzpqd9M
4M3cCdi9yEuCZTDMnhAX3jIwgE89XryLm+IG3jfoAUlIn74AEeiiIro9PJnniEprochXUEAtny3K
lco0pj//Ye/pPizjdNU6RJRQvS/2ajvBxfCeBHcPAuIGl2PvYlwjRvX6uNoLcdR0NRzR4wGRNuNT
6ev299X0L5lbtS/mneifbOMA6fcnA4aqZ4nVp9ggUMmlesya8SH9N858c3prSljrBv6VomYqkinT
gmn/k4gBVbz+tz+glpciO4DbWmIgDM15fGZLEE+zYin0sLunqNaNHMdCIJgrIKPahTusWsZq4s2x
1CLufk5Jl2vHqBVO5DJV3hOXM4l25n1MOYZyhWKDKluXxpfn0GDZGKfVwl2eLUrInRA7TuOTb+ZP
8L1Qpq+OYo+NpNn0eQbWAm9OcJQp6+ZypBafHTB/mKa8G51k31fR1IZULwt3CXSkQYSZVyzffmTG
FakXgay/73WreMYmGCfuFjrfRoHY6jr3PcFEtfozmzwMcLKilJyAPC5D/j6Ig/7IKR0NRXq4gddE
L8CfTDQxKTNj5Fy8boozj2wVaRTBM0kOSE/TSksHKZCTFFqAM1D6xwnA1O7s5ltxOTrfe0IOApPN
6z3Ji04oyB/iNhSyGroaGJ2r+VNnC2jkLsY26UenCwnkJtXpc+2rGT6yOmhgaoSIyRK6aff1KaeB
BNsOhq+6Q21azFvNuGnU1azV4iVQcUQvJhOY05c1EgDcBF1cSdgK3qnxdMpp94KENqfTuFoeqjAs
q/bxN4cXT84Q0G7FJY6D4vNBNF+zfyy1wpOmbohuWXA6i64d458ig16ApzeZT/23YJu9csmOlsXq
zTm4BAw5tjInh1DxVd0It7MJJ44ej4j65iRL87WYrAiwdEqyBfhUu29HrMm1BXAk9ym2YPsuYlIX
ArXD9OAV0QaNUHD5rP5cdcZuQoOYFD8fYpSlvcCAY1yPhN2IUCXmCgzIIf+xKC7YNUd3gsyw4ZSR
hu6HizqJP/Fz2yNZiR/gKouOxi7kmk28/M+dB2rnr5ztBjMdPlFZI1/fomymde6gx6Dg7cdcNnnj
JigWZZ/GAYJAc6KnQ2A6luHB1Rf0pfg3ZbBxvR9mxPoZzeUgZaJYBsE37Vy2npZC1txMf9xNF8sR
t5wCm1DjHKWxFQDjaqS+FlAoQ5VC5hgIA+OwkufXyrAvCy5CDTdt5/RpyiN6EsCDY6GMkRKnJfhf
PO2kYdDwi6jdhMJPt3PTgmwlJXFDnhpS5SEzhAZ3YRfTcAiblzPwDomLzTQK9i2MoVrNHwdLsZRh
t1dcRzNYhMZDKaIpIeLUtOCMgHaJNhIgJLVlGT3n9iGlH04H39pTH4933x8uUd6tG9uSmwL3PHwn
MP0fmAZnpH3oxhh5db9EJIGvEEYgbNCo3YzHJPOzfSHNUQI913RnO1P53A9WNxK4G7yR2IYAt/wr
qR2+YmifQp4B0mOuUSMGxBh99+zAChd0CuhEBBGj01HQJvjcByelw2zlBAIfdELzBeA3LB42Wm94
B/V1w0oq7W+ccg60l8gdRindb9+8lBlr5niVsnD2oZWEhanWW8go6h3s4yd/5hsLgaiGdG4n0i/U
Jca4p2m4ZKOhB4+4R6AiYd88o99h2i76v/3pi5XwX6loqRFgnxHSXrKkum3PWEVN8I5WRXYipkVM
cFZuRsnNk/t0gQFhysPn7djeW7NSMpfC9ihMtjNYCiSP0Us6VLCRFYW1cz9G7AfcOW3kwSHHNwxA
4nUwZjB4J772en31felKRIOKHbETOYYiUzNZEtZ6IhgrtaFDlTPLhtY8hAxJ5+rdkW+bJoLPhjLp
ZgNW1Tz/kqU+xUY1zEiQlKKbsCDRnsUxJW9LzHAq0bqdH3P8HzB0ur/1tRMrHDCRTG6ntTQsevE9
CHLDAr+UKJqaDYkOw9TE0gmvvbkuz58ov/zPhxm+jtgSNh+y8WXrQMVeDhc2H84nixHNsgpwWW5c
EHxysmRTingp62j4n+iDN7sCCrSH6ZlZmbJOtV8+zOv5EVdyUxeIYVAWUCGJbZStD4R1nP33YKzq
QKY6yWElTP9P7YrZ+0JiBafF7jZbEzpC2Z0/LwdDaCgPokQwK/L/dB8dMTtRsM3lXHC33/bxqes0
nDU+saodFR79FJU4FqAg6h6iszIuG0bvFd64M7n0eWOGhdc3zOxIQERCln+K5aqzsgGydS45me5t
yKsyGinHI56NVH612PSpVCf4i4FtCX0Ffvz4VkKC3uDgNKNzTptcACTcLLLlsU93e4ge79cd25xl
gH7YXo4m0aJnNp79wbx5CVh9Fyoi0GP7SuTlHuT6mkWZA/Opdl324UNPrfDxbLPGmX/O4HTjSFMS
VucDvyjU5+aRmKm90I0ao19GevScX+6OX1PA6Nu4ek2RJhZxXZFxBNsJPQiFYfBDS/ajzflx2JOt
sfEY+Lm/qE1NZ5YoSyrjVf6dO4H5xH09ZTSzQ5wvSuzXJzIGBKtyD36RKTMa9+ySKeIOdsm2cj1m
ZUg0Xee5O0u84vanc64ZhDWAh3GvBBSGC6pmaytPjTiPgq7Ypco9gkBoSJShfjKVMtglQb5rlyrZ
RXp3pne9ch3m/mzHf/tJywbJOvK0AX1wrzlcIesdHPTjqXq0PV/XC+TTpTJiGYBpft4vuODUntz3
qhfCRFnEsmNzZIZdEl44POlQyoIiR4hSSXKidxjk2xau+D4SyrO7AvRe6pAP5hnGd7Vw7CfDGwtk
4uphbrx3PrN493DM+woNPSPE49jUTbLwYWWU7TxvawfDjonxI1dHcd6EuBZ+tbYlNkUTZ89cT6qt
DIKZAOu0LMic+YySVDVStjGQHsDkPgQSX3LJLSxjpl/hKPlUXtn1WE+GXIT/Y2Nvhe1qDNFoT9iZ
8fdLqVWnBakQZ181SryCW4BeuG5RIP7ewWgTER7JqDMYYJ3c4cdolqnqGuIGnT520NRsd5RrQoIM
U1cG1HgH+RWfIzvmAzlhwBEz9cICfA6Jxh6jXeQurELlJ2++m6GrxjyWOYE/ZuvpnB/AMlbubjB4
/ivJpcb6yXAuUDGpGdAarVSV7o76miEhw3381SgOUyvFuRYusAKV27HezJ/C9Ej0ENPqRparqaHD
6lnkjkjPwfsBELcxINS6W2efLp7xwzx3ZHQZF8Y9+lIxlGj7zbOqmXwZrqUmjwkJAP9mhaQqBeK/
iULE9EaKnWNwu6r/LOOCqlvVCTQC5mfNslJaxAZCyhJYqmwEhQn4zB4rT3ZvU/YBKJhIkNaQqjMa
e3nfUxxL0fJZx/X8I9htTjPzHtMicchuABt4NvL7tLtUe8HQk0ItjLDvUaT/I6+jn78NHVnRxMoW
wZLSFrhGeJ/r4BmlfWF2/zo+MLUyNYkbmrnW4fHYF0ldNf0aiyaXDUhlCLcCeb+4Rf9WfKa7c+UY
EzJY2BajWkH5yIVwgQwAUXyaZHjNJW6UmcrZlY838/qV+nOGz1huN8AVBJMEmrYHMvFttWQzWpKI
Jbb2XPF0TpmEYNl/Ra4xaTqPo72vFQd4D9obC/mokvW45kqR5JrT4Efi1Q6hDsP3zvhXZDHu9u/C
P0ie045EUGuy8s5uBSu1qLkyDUowLY2jUFCJeznu73W4Pe1nU7kSPv6LqFdrnRAMzuBemuU9D2la
uQ63IqwDTSBTEIPAjkCgt5748i9wlxY3Hll1jhHvZzDjM1Y4nB+xIXBp70MvyrSrrRQ/tudwZ7w2
CP95d1Wgvh+nE8i3i/XqDj7PK1aTJKJMYoSygK1cs+GqZCg5rH8ZcWJPrUNLokEDDMc1mu1/FcRG
JalVzL5ZDkQgMyNhx66bNaxSjWHS8RguAZR5FQjl91GOf5h/+KdpeJTAZiDl+fw7qKO+h9Athu10
SLOIdH20ZFCE9pUnkB4dXQw/L7jwh58OYuX2FWy12U93+mnhn/X0La4FUpcZgiDuDodw+cMWByXy
iyNQCDZ+GMCIVff6jyYvaKA7km8/YhF6e6mWqrLBar615hrJFftMkZcbIIM/uo3omwHdXkXBw3jG
mawkbifjzat26en7ywgtTk0YveYuXfMHwfgR2UNx6wWeN2PT6UR4e9oq1SPwFe23c0VgJ8oZw+ke
fuCKZnSr/jKMdnf1xCQJTj1joybOwtJLa1QD1BbfxpQS+36ggX5T1idyiOmwjMev8PRUiOvYAr+b
H67wBpjWN9YZ3TFOonbDYKFQS13UuHEkrgffAqEGrZHW4ww8b+xT/XIAVGZS9nAfJXUd/Hqvbf/k
4hZBb8JycJi/BdF/eKj9+BCGlbtEL+3Z/b74CM58/IpK0WhVE6c3gKwB+aHZXP6HhSRHde63orgP
feNucjg4XzXeiCrUwp4nhWkQ+WVZv1dJcAZbz8sCsgL7gBUaBQmmMktnry7a6e2i6Y/oFKHQ5Efv
yIzUzF2Z08oZcX/2orfw5oAnueqhdHj1JAgoH/+e3iVCYthi1t2aKQHEVyfZrOmj6Ic4Ekdv9vVZ
By9kUb2bdAYH7/sySzv9Fthc6EdKZxKFov8cFddAbOT1PER3jpwqEuIy//dRPEGYIshBztKTJCf7
qt4db0VtAuwytBlnFNGeKdD4Ojxeq9lLQzCK9cCc9At6LVH1wseSpMksEnEYoBSwsKG0C+PVHrHq
FmuIYYeQW1VWzeYLpEGbmQI7Ftk8zwY+zwQikKYYw++QdUB4/LeeEjQGU/+U5LCUjcK/3qY7Q77z
fUl1nya4Musw0jE3QelfKMxWAX/YaXqoFNpTYjwT+wn2MbULpvDGYT0wF147Hik53Bm3OKd0L9k3
mKQU08nMNxyhu8uKBztEEDKgDYFfk8PimncFnKgAhWQJcSD0Pd22VrpxvoVxHAALdUOBhAD7EqKB
TbelR/qn2GBpHAvX7xbZVZmS+7/WTfs9RMC/oN2X71umoAbdUud18J3b2qQlPe0tKrHWwahp+2an
NTvFzRlu3qwofBCTwxOA5NqxeSB4Z+P1kZwmchtJUETgzq85c1dBocExz27efsWRuK9kyDO/zlvC
HU948j7iDGKgassWbb0ht6hdAJ/vkwBGVWWBv7a7fxvlY9vPAmiIqQKcbg5I2SAT1nP5ZwWd3J7o
uCx24JatKaw/F5v7jRbkvnJcn4HS7UD+2+IPKhunQFonmn6yH/mSLfDqqIM/r4yiBTsPU3sDwVoZ
JRo3xCa3qjoH/otv403w9UBYUS0iuIqbaDiAj5duhdYIEQi6ji14uTrv5o4x3PMjk66aHJ2R3Q8K
Mf2LB+5qgXfh70huqOQ2J7bt/oX5tsRbTnlSA6r+O/uqmAlbHKuenzi4DgNh2htapHQcJHPhSh0y
gTUlIOxUNGNIarkKL6WP7yKr9wOmgR35B15myrFWzDlKN9FowMrlZk7DV7jVbrxcTQt9QNxwO+y2
RgDSrjdn8+plxjiDyFp+ljfzZ4YRdftzNCr2hkwMJlmhRmkhDjU11bglNhJQOY/nawzE8s97v+Mb
Xqfu58CLQyzU9TSJQbRIb4rFoWMOveF2wjhnJBBNqW1MQl2Lh26sJKBnIBARUsEwagtcP1L5hcWW
RRn0KqJNujkB5FvozCs5d/C3YWbA6D16ai+JQvKd/kFVxSnj0H37nulm7lOI1gcBWlFNqWC/opmw
Ts2Wlzm4vbkGWV6QrHJKPFLUSRnRO66EMDX2vcLiRqesPxtp5Z7+nX/Cu/EfnPJrEEgExYvxFugs
AhUKYBBaw659nYMta5KvLQMTxnJsjb3PG/R6H3buoF1xm8eSKJboi6A8jHnw/+CwfctdCXyr838G
jWtM9m+C577GJXbHA9ZS08mIOyipcTN1T/6zw12bSSTwNO8wVKmgxzpBnJUyArA677CwQZE08pgp
4f6Oz3BJCzAIFhGrMqGOklqDdPW8G7gvD5MikKD2kFHQFwUNkdNml7uFHZlj9b82TMZSKyFgywID
gUHEcvWPrm/UheO8e6heI7vSp63wXDKeRwHXkBZK9UgoQwMAOmEMSqkJrgYZ4I9sSqq0N/krK11+
fLkctzvoM2Yd73Q2StBfSPoaA7kcwDD+il3WkL/0v7vu00NtJjCTrIEVU8Ybbcsy4AGS34I4waqR
T1FuAqIJkv49kLgHtwvrIDsEqVpL7attN3rDpwMaY/fDXmPd4u1/mAHMXOzOQ/3JYdDN/sHfr4YH
9M+gMnX09H7kqhex036TaC2ZwvEvbc90i1MeYbUPRZ3kG8YPNH4QZs2enddJ6eJtnwf0Hs3PXb6M
78AOO0BoLvX8kkTtB5mvySwZNBCM/+v/JKVy4y82wEy7X29UDhBYPVEQ2VpJMA78I1EabIxURO94
VxYZWLNLbKyPtOQ2+cX4V3qgeCnP+1c8a/ZCKY/4lwdOWA7RKTNga1TLkZMd479GIa9qOoW//dcM
7gqYrdiPZFCg3yYgxRCKP11ypoFIdmUX0nrvBcX4Wi4QORKxzf9YzCdrlSAplVKt3w5PNbP9uh22
ZNfX1otoTC4EYDrd2AGEJf3Ud8EHP3Ixhq7QJJQfDN8Hb+htIgCM9TarIdFbRa+kImrxinUD61Eo
kmZ1ZyWmsMJZBSSweN0QcjzRcA+lcyX5xYKZZ20iWE9DUOkKLrKdKdPfFfBwmDAu4AtcDdDqTmkI
q9luJDbTeKhhB21sspqiqOPOgYwSAUvL9D485Z6e1eDKVwPfEnr+vDeHTLBoIBEdX07YJpNXhLbN
VYUZv2DV/jZ43tSTQB74Btv9vxlBE/ATGlj1WOJfXOqh6br/XaVbEGl360u23G9XIbF83zgVcZlB
E/8C+GaC5dL33HZP0ss6leVQLpaqYk/ASt+LHDdAjEFNgKBg08fGR7sH9OhFQuKxuIdF/fHzKh5E
anbad4em4rpiPjkmR5t8p1UFiohPmqAnMmsPwwTwEBfeBIt0sKwADKAmi0bZv29Vx5gDGCIfySWq
XksylLrOjP2H3obMjISMzvjqtOuad5cTAgYFd9T2/7iRBJaZAGD2BuuQPFu2ILz1MNAFRcRGdY1X
SnHIy7Wgj1hy5ZByjmOwAmQVeKXKylROrIdTgz0De8UpkeAdyBnS7WJH3stkbkaUJfFYmRhKMi5X
byEy5btw5pICCZluvS8QqvekkrfmVzfrl1NGeDHd9vuw5wwfShyjwN7rxZ1E9pU0w/mdtuEO36A+
giX8ZSplFxhmKTfVjXx6dv4UXJ8Yow/Ciy/24tlA+IGLmtap8VLuHTDCkRzgKgVwd1exi3LGwTMv
L3gwgGNLk1gwnoXknAPBqJX3WolVVTdoiV4EpxjAMpsbuS7gDPUeWC2wTHqGc0+HsE1E6QXoAAn4
l0f9YnAFgQBggtIwKZbgPAAM4MPz7NWOuSZtW4m5XZJ29fslruwDH7tVX71R1V3d1zU8y3U1t+Ft
4s4A6EEcy1nkMybAkzPNk59z8zC1b5ntIuTvRGcjEDen+vnSIhlcCJwnKMp29T/QaJbXGW2Cx/qd
zFp+dOsOBHPBzCEoKQEqQYCLOgDmapH79uUSCH84XlqQuYmjW/sOBPbm7rsOJPFTfh62NADuEFAQ
PdHGLE96Ork1imim8w7oEmvt8TRBmDNHZ8tNn4mRNC/zJf/aUJfIcK/3R5jjTrs3yDBFcYKcXFkh
mWMNEwjXL9YLnEAZVa21OcHiYWYcuy+z+6veoT/fcHPN+ZoyAd8KRlDnth7Hl5SGl5kmik3pulmZ
cdNyX3WOwCU61Pa2vmkObHygnz8J68Q0CQxcBzE6L2WbhogeLPKFD1egkaHOiIo+ADONR/XbZ3ga
oKI4PLKKl6XdMcnKpBFW6rVoD/CE1BznFIBvFCxfuzAIOxxZukXgiSMXExW/CXyBdj5EKpS2ncZR
j6+u4KodZtuXE6D++xBtq6TZV1TRr97Qay2Xk39/YPo1eInYeWY3Ii+ajTgcUgd9EtrGB5orzgny
W7UUh3+9exlzVtgg+9nZpYnHJp87H2wmY9YguJ+n4okJUC4o/iPyJDizNiGhmPvzpwuPxfwiYQxW
MX98HP6h+o2DeDJDJo0RnuW+pyjL5eR+Ul/lhbU2fuYomlZsIyxr2FTDAKyKnRI7HuxR5tl//as/
8WOhqFpYci0eDbiny3c08NNmDE3F3vpinCZPJ2vFmokZKT6ggblf8cMtnQF/QbV1K4hMylGb2dey
qhRvjJtl/h1IKjkHHzDBmO/WhwmVbVU+XNrurXZDUmR1jD2db6LmDUAxJgk7tJuCG3hx1ftAm9Ee
8gJn4GSIIFIxFr9VXDKVno7BKwlV3JZMh/GucaG20HMSi92Q4zBhbjWI8sCk3GXd9qJi2ioC6eCM
LTDMSMZRgdMcXaiA4BwsNY9guqctEQ3jYmKvon/KrEonrmmNgPVtUuDpRvhcRPcFZoGqvNSHicpx
viuFbu+FE/YLJWKL3phVZpRXVsBGu1iQWpSkdxxqbH90TNAai7ivp8gT8myh4QQYnoLgzzd6H6et
R0uwDOFwsrRq2eFX9TiUiVWTKR/MZ3a7mIiZhtMjX0/9JAsXa1RQlJNY4tbiKhyKgya0vGg4mC19
VqkJF6H0xnwvYZcxuTjA+P4BBoBEqNJMJw+JJt3LmgKR5VdgZy++BvNNO0aZbpNjI1V/e1tpnBAs
G1uAx66zF65F+wZBqG0iq/USOZ1ONo0lhLG4zadcCk93KLCFpFUDzERtguCF3AdsLxbvmk15Vbj/
WwdIa8PwVC9iLX5aVVuIRRkyyGma3dK/LSv/wjbOf4BggB8EhkFFGLR992O/KQPTAYrZ2By7qTcO
nX3YIh1HAJGP7uARXDMsTx6+tGk6uKomBwZKBePAPgCUDPbTy1JOjalrzO5hHpErNJ1KLlDzNBfv
SsIrwBv2n63uGOx7yhMHs6aaKNLx8HzmjtspTvO6WJd+UIjdbHPll+ChIzNIBeTvDErQlnBIRklM
vD0uzAJhBG26yb2QuUDWdW9bPOs8y9x+WQJ2wW0xGBHEt3M/RL7gMecRhgiTPba3RR1igeYWmPUF
DtNyl2ppxeVb2MeKZ9Y0nhbAQCWvn1qdzw2BP8XR2vCqBD9kcZuj0Po9xOS5Xt9VXatkiSt6hGpV
sDPamAaKXkeDIozkZPMoqIjris0lkv9sP/0J7P2FpYkJnAG46P4f9m7uYYTgmF31p4GWPx8hp5+3
z0vY0vMxY4crI8QB3/gDvF6KhJDQ8/K27DswSt0xWkWXwxbasn4GV4FC7yPz+S3o0IQHyittc7YV
ow28cJexewsmluDmHc/tXv1gkm3kosJl8Kdv3Mi5MtSa9qDeG/sW0iFFicy7ph4p4M4UxxzQB9p5
tRZvU0MnDj5/+8vExFBTNnEPZFCViX/HqD3jZ+v1MOcBWJz2IZ7VM1kmSWgqHG+epUUtTxJYZTdS
f0bGlZ1Zor5zuJpgFB12VSBkUuJRApIwbRPtA0zNhJOgKurXNWG5mh47rNAXjtjQFskYcAg4Sb4t
/Tg6c0Sm5LSC+hCAeOVYRj2LSva3COF9oxfFZN3wOF6oKaddjmj8BaSP5vy0qoGsU0RdOMlPyM35
u9AR2hZpxLfJYG5j3IPuhTQhepEiYk6G/k/NXR69lIaiQay7ub+JV6K5S2NYZE+nWDWYaP4xuSX5
H3+EUPKERkndpW0jtP6EqHzKUdab8m76l5oTI4OqwUWUP77BqD3hpspg0RlmjwwA2qxqdu4PMpUH
TxdP6ZQxLOGV273sAdv1ij8Z3xC5ySqXt0zoLPC8hKTF8tzwLrP+qy9JBXIFtwD7xboBmD9Mccco
nfc9lLYEteBJ0X4klGrQBo2k+KX2GYLoXFkYfvHN2RW8EZJy763MNzboomJe/KiT9stKqYYSaJaM
tjoZncVvedB2u+EsDbZ1VFPncwK0tdLtTOxQpRCeKbmzP8YZ146yW/PDilxVvSB5qKHoxG8ef/HD
RIaLi61z8WOBYr8PeeDmHc48h2/5qo2RsWIVdEIfs7PqlNppDWqs1ayZ7EP6Yxct6Hi4WhKyNIvj
Rg7PinAInGvcG8cnw72xogMxr7wTJTAQXNTTbzklOdGmoegJYeiHW3/VOTUiyPxAj8fUcAym5yn+
4bzhLvO72aKcANZh01Yn33A3wWO/e/i1CILOKx1BQWkN6eW/nSmcqneeRSpup+2Gw0u8T7llorxb
yJyexvjfvtwQ6x40+zuVsH4xM/cMpHgIYGFlSv2gPUpnjMwynIGay9vGTKuwN/bt0+paKtHlBkbJ
M2WyKUGorlSkPjMlxrppSksRAJc9cphAMP+X9govh2RS9mkDwW9QVvQ1HbohzZqZlKgRGJrmtWBg
DDvJcA+PC18X0Z86YE8LzqjRRbUWl7Nb1S4um9zPC7EwqGCjstixSBqjkvyIM5cXQBbFNkA1Skyj
yLA30oZp3yhsKHwG4U4OKywC+5QW9cP1v34l9l78UqAFWaDjDhxdXEuFCCzXu//0BipGw8JBGHSm
fBcpVWv+Q1OEtLqQ4Tu0a91G2xceQ3rVROO3HPHjJ/Xj/1x2aSQoq4lY9nOUCv10qKDUKHVdKib/
5mIbyye63fOiKrpKMpb8OvD8V7K/fx5H5tJJbjMP+wF23s0/xJyKq3ChsNiI39otiQyxp+PZuqsy
n7Xi2NkO1M4pfY/0U48ZK/xlZbii8sKVTidCCw0RlayQ/8+3h1a6wm3sAeVE8bN8cLsMcurGydzu
IVVekk924y/F7G18bf194LFgBlJMQsE039WO1cRA01LDiov156m5lzbaamAM/+AN1mJdtUVZOvUh
0RGMsOlsBrJZaj2oqf5cTqJb+tUGqMtoyLRKALTZZG0D4x3l4jwBBDMrlllu9LVK+tDazpntpwGE
XQ6K6V2EW07niR7j0gF9Uj+2TixnpSh2cxzGveVFyWrkoPXAcapFuqwlJCuUJugHlataEIJ208Y9
hsGIVw0WqHQPuqKIVKPpsWFDDHte/WS7O3ncTqxEVuytVk8/RIiqik2F66vhtyPHriCPlcqBtsk1
Jy/0NCvqmeQCORgyHLcE26HjIxWvrD9gfkKheJFM4Bd0OEg0ASV3hinEJr7ZVYPQmjInT23GZA7A
8IIMuUsbcf/Ny9QFz3bG6siiblZV7a7sI7essvNSdLnTRXmIzqVRHg9iEGzN2BUhDUKEortCMlbz
ZdhZy+4d/wrdQcJEfvo0OnbGg2Z6hR6DFbxgNVvuEdyTM73M/xkiM3A3t25jo1/x1htjMF3KGnbg
kzcqtP8z7CqwxjD7Gy7+cKbmav9O90mJ9oZKflfP9hengiyUZ8W27FJf7deeQKYb1XRHtZE8RQeE
uaA1scF5Ff/z3ax2tKxP6uLev1ak5yre3+UAUBLA8ngPlMjNA7g84vEbjOGdleHYT7deKWo/sYIx
NPc9xNgegHq+LueBBfOmVcS6lj8+evrHBonTa/fJ46jOGYpoECt+H9CkQmlVYbzKznTf+d7QGtpb
g4YTjlBrR6mcKupLeJe4ZpXLlAAzaIRovPhhy8ju8DTtTmzegPSywrq3SfFHZWiicQzziC0LXjYV
vuEx6mdmNd7tnW/bg66+9c8hXk/uvDFqh6o9buwIMgrLUox+EsBvhMaNoe4+29wNWTGCklZWSOjq
cf03p9dvq90bbdNdGO/G4qR3TvrZ9Tioi7ea8VBJLZuXaD5ElM9xFeKQiTeTA/5YxIcXI/zRdXba
HXgMyFWwer4oJPkCtGyCyzCcLoe4rSAHI/OaKbspTSVIofMNCGdM5gqYcdtEMBAFXBjSi+8HqiIt
1P3EUnDXw3ePeL4FjZINTXF7+fVTl2au58HT0FN1DQlldhgDKLgShmPb0ydMrNBH4Zm/88NiIPi6
ooOQ7vmeYoosXnKXsghu/rhnj+NELJh4S4WdEbIyTM3cZ9iLikabd4z8AwKkawvFHmMUwKZaVjY+
zsaRuAsvRCnOOMfiZlRzhM81zjAEQTKyiU+5ynX+IY33/8M58pBRqq4G7UwCtOB6ilfknLiw4ECJ
9UDTZt2hB4t22kOuM9knDhNTx2CXQkTviNDzulUNNSCDql/YmEBZeVe1LgB9DQprtRIv3lD4PNqe
jcJn4mtDgGymlY9D5vT9voXUZMuwQEa+ugvTEGdaV/MK7i7OZqqMhCC69XBgyG9RrJ++VbuBckmO
d/oniXcuH4iZqWhU7xyCyxE5nRbqIaio3/LuL1r9mQ0xCIlC6fceGiWeKCk4xS2irxlLULt/4wsG
NJUEFz4oNI0kTPTincWSYwvSrehFtd9zg65SsjUjxPjMfqJWcSki8Dx4GN79a/Rf8kTA8avnnuae
zn3cuALMcvRsDNPX1HEInnAxJPWsLtf8bKZSQiPrXYcn/923B4ddW8OcrH9S2Wg8IIxRIxJ0vDC/
ORQydRv/IT0ACbWKLJWkugLT0n18cr6howWBP6nnwQmEYqRQPPw+tahGG0oQkinmeO3pb2htbhSp
lhf0f25sxg/pqdSZtQS5pCpHFYQyRnD+PW9FcBmBF7VvbugiyEUOnkQT+X2Y2HvMG7/IvrjpDa/G
p4jWUekELjzG2BPKs+RfX/+FhZJxRsMzfTPlINbHbzNvHoKncffHeZ/qzhZGi7bKpeXRz5KwOW9T
GIoerkyFuPa92dV4r8mdI2XRe/f4Dq5EIXx+8RLH53rXc592MoUPUdgBzlH4uodNb9fvTHLT7uGR
Y7RJ+DcBv9kyAuuIf+jxHXkrMRW9tiNjSDov6RQeZZJd3At+iYiyeOdFu3s9YO2AWWRrvBO8bs/Y
ByJV4SNDTX/M2JxLaG7llGta/aFWk9h4k97E2zaj4qUk94PVeDoWDI9oIym0+q+vemKucsCesoGD
quhK5YBSWPR6h0LX3fiO/XX/xnFFhAGYXmwp/ZUx5ifDeRK3uoAtLaeYHtwvCBrPebXcSZHCVYkq
KKfyxhCf2vdM0BuGLNfuffhhV6H2Wdnxw1Kv1Se7Y+UoJYbvEz7C5naldQlbKeoVw/z5OfUIykI1
OMvh4Qlz8BO6sFZZP8ppiZFBb1lfs5vpBR4PmOc8WZDeke0v2XGe7SW+j5PLSCcxMBvjr5VP0Zeq
quacJyQw/BrXXgPEvBySYIbfDNDvOrvoSTkTypedTfeWGv488IgLzqnS+p6sQj9WcfYRJDqDmhP/
LstAL2jhNJUM0O26lQ6a/ZrFBAjJT/EVEif5m3nDt08ms2KBxh5q3wVuzTHSnEna4xZKDJxmCpTJ
rRfU1p5O3f+uUDE9lnPgujMRn40R6gQWw0+itN2mHJ3Roy+gUGZQu+qC8LjipsZaBPy+nRHfRp2P
4IysZfb32NhaISPxJou1dQ3VN88hH0MHWqs2ixUqAXVQfnPCOJY6vm3AtxAhkIzL4QIqeuZZ6X55
4i1l3O3cKVXz0ubRCUNfFtBYuI/OKsKL3ZIeht9BBKbP3okronWTtwLbxZd9Qu8m2S05GiHVf599
7kp2ZbMBa0LgsiFR6CEEU2o44jeujjHq5hVcuy3bnY6Fv/+bBhOaU3zoef4dlYQ618UjTVJtpyYg
EntHjpUiUPTSYOkhY3E/7vEoX4aX6N70kLRR24rB7elVAvqaz4ipF+NVdo/8cfEMIcMzcoL7mP9E
omA3oDNzS/o2SvyHqE/dtdA/fStAH1mjWlO1qBQBbK4SJ/L9jncdJnBFYGxkS3dff2yti/dzqRFF
P+mnyHdnnA+LEAPuYb+CtlFb+VVxR30YlkTTWjValfupiAu/dqUt4MpOB6B1KiCNpQdiCz1CUL/8
zIFJqylLxVYu2cHReoc7DhpqgGORMMbxXXjEdbMo/mbwOREh2WSO+IfNzDtsabaGvAEDYbrw5Vcr
VFhVPrT3CG63aXdXkdnWZk+g3Pauql0/0y2msVOBAD+S1+zZAs+npX6oHXC0zZgTfXIzUK58Mk+L
KiPb6JDL7lemgeuG9qC424wdPtY/sQU0PFB1AiCkNKKQ/csVRaRnREfUqZEdyDTUAd3x2GJXEdvU
LF/+ijFPjNZ+NiEGhwl/7vCX8rfla24pGiygXCRHcd/ioAioRk0cwv5x0rw/Q9IeSbdo8Q9lcqVR
3TNmf2cKNFCEaoroCYfTtMfDYxE23kv6v2MMjVGMXXpSseJb4/QPI+i+4MGoFzAwDPhYoeeH5igq
G7uUMfHXnlnFxg4DU58dzHfXnBd5sO/Z3oJBU9IOwEecAo4PqmEzd4zu/aMszoezVJdo/TVEs5sH
0gTgwaL3FJJ8Wf05naUDrXyydgDaQwXSTHFwujRtoAvTjsuslLcAaW2KLnqGQ/2o0cC8U7q4Pa4z
VOoFATNygptPcrBRwKoCig8B/cbP1b8DnmU3amyzh6R6s55WSMG5rqQN3H9gSzXHCQu+etTjD6/A
dn1FQAehZ77DUnhxql3/aMY+WCT4FyT99ABPtIXmrMMIghxITQ6ZQgw3wxcbtmgDn2Y1I2k7sofV
hpF7KOgOnF1usVcGuRz0k4bKmz9rmPc8mfyfTUonldzHQzhODa5HAo8kWHO7wnkALr917K/uHeBx
lE7FSiACCgiHqgIa+wmm6PHXIPnnxuKUleFEf8heQZl6/wrPIXqvag7owYyGcnKmITp9aM+Fr4KI
Hj3O4TGh890SOGGkJG36yDmC4BehxKcG6a9WtpvQdWOl7+MIY+tmmJkd41y7W2F7dAcrztIsM+vh
dfsZNfqSBT7XsdudbLwNdjEq41YjePkE5mrtqtgkn19i3yYAplBNFZ0v3srA8mH8WlfqqEPk1Yot
bY2LEms72UbF91rOWV9HmrI36lsv+3p+ZPROtbBLHlc9QUWF1GEehkufbXZoY6NLBt+4hr/ixlGp
hs8KwXd7kQyjpXo2fFZiBADuNw6nqIj0Exyr0JtfMkLhc+ELOnkAIF3aLrmBHWTveKBa9UpM1KAd
M+oI/5qL8EPyWD71T82ZiUi/NAazYtAqA+9VFWdWve1ra1fiKeurK4Us2nO4K6tLwF3fvHUWUYn9
z6SYH2jnMIkxv072v/ohPTqKOrMKCeeHeZygYbrQmmbKtAUO/gPc5fsNNtmYbylKKpIvrLWH3NX7
D5onJZvBNUpwO4KsEc/+PaoztDVHHhQLCmcmr1+AlQBw8oxlAOq/rk9aZzz212xMrYhN3SoRbpnK
KZqhU9PjpgJwAaY8E6LrPcIJHK9jP/AkDzzsdCarrMncECaylCl+x1Dg4+PNNPWCoF+mAh6wO655
hoWjXAYU8ZnZnJHeb4u8TzoAjv71WwuMFOprGwLfHpqv5bJAmuvhcJhc/jX7Ujd6AlGhmKtuTiVI
vBrACFTYo5L3IJpwEpFb/QhAYfApnO5Ql323mYSs4POnEe8vGgiw4UADIlUYPEeKYNO3JxGwhJku
zk6sVFhBgJTFLlfo+Qin4BCqkSE3LURK0zF208Wu3prG+ycwGEQZXIe24noJKHiCE7NK5rwYYgsD
o8sBdsTNNvtGCLTihBFYhGbUDNxFBv4jQDnMU3IolVbrrqTlxNFPAN83BjENuXND8PlCcDDj8R2C
TgyTA/7aA2JolCQa+fO4/odF31M2sADK19WDTcHdQM0enk4CNJYfNK1bK+ovgCBfjHW6TAspoNjz
zsoXkGRfwwHXvAptoheHyJsp1fu6WeqCL36xRvqG1kqIP7Eyq2rIupCNgbQCMKW+tVYfGgRMuRtm
zuCNwVz8+KVIMgiBxzTwFzq3faHFWVWodMhM+NjON8uMLQxbQytqPhc60TDhi4NUvXFeBR43NMBg
QwH5/d3aZ8yHhIT5bobK6/WjSInuyufV5h4uAiB5o6dyb8gseN5RDLn6HX/3nWPdjO4GMhjJRj6Y
+wgaJpcc9C1g9CaCrW+iyJUXtkGsH383PCNBkLsx9BGvyqVf225vuFfi548wF7ovQQvDsG5pJ/4E
HK/pNAIu3/Fe58C/Ka+/mU4Xne+yrWjKjJv4hpPxd9EyMAhZcQlHvZGC/3ByAH5KrkxeCbQhps8x
WFuzErAorQ4c4fJygkdpIWtnoBnNnjoEV0wFNqOZzw78tpgxVUXHxpI5pL5z/HhQSnt/tWdst4AT
JMkzEz4vevRW2Avfh7SFkBOtk72aiIbTcWZ7d0QcTN422AEM8Et/cYDIOmlYQLY2VRHfYYruz9SD
vggWweEmZzyuKRrM/fDjHv15hyr10FqbpcJsKivgO6OudGDJDNMUj20A7KvGB/sid1t/J0lPXCqE
FHUAnhPq8phg+wOr4bWYWGn0eKRfYUUyOkYyAEFQWp6SH2tFTDG6+Gb6+SVEqFr8qwFiXpdcvFP4
UPBKURlj0uL/l3KZz48mdFPVHvA1IVZApVIwOSwtclT+IdGQbkVxh+WsjlcX+H8fC2gF688k8d4j
Tvrgt8nuoY7FcJxQ/F6dauRD6vlS69cmVFIMI6TumadA0BXsGJBptvVdMytd5Kh/UIzHBiYGQHpa
8+u2968PIJX2fhlrI+kevIN9FVseWYvBtMdT0BnJukRgi1OT5Srh2Z1h7kJhhVGNtdtMSYGaY6Hu
4XxySz/W5LrkoXggfz5Th0dnLZ8NQ83zpT4gc8WuoiEN1gyB0mouFt+JrysdBZSeR6kCILW6y03E
/WocvFsujtA+7jnreAfd7UWa/1+bhoipDxQSwK0pPbPgPr2LFIKKOnw7bRLAdspfsoZcNVR3Og7W
GjoO5DutO2INeRo2BjwlxHhzk765Yn9mNTk/QfE6RQw8vt+IiUZtKzblfKRts4+wnKu6orxHrxdF
mM78oNZcmTM8/8yzJS5PSrvynFmPZTs7TU3ySV2FCB03I8IxbjGIXkmNQ2l3BRwdGT/86Jy8tn7/
o1RZkSgs6Uuq4oi7O4acCuMmniY/vbajxJggVBuPjgaSHRsmY112cVbrMVMZTWZyzAm8ZHErwB7M
RohqH2/ANcF+lVz6W1u9QqJmYz9Mah9p2KNqrdKarTFnMK5gHAEbscICnwecVP6Nb36J0bduw21p
JbFalm5yXoCNaO+iO6CKsjwziHJm7AwuwQxIcz0d9TAKxflAmvbMlpTUDIahqiVM1p2pTZ4YGY2+
Gm5R+n4vAhTOjp+6Y5uPJbWv4iw62UANsCmSUxdhtr+uv76HW5qA9i5xdTy9RO0rJtOFfak5H2Od
ePTJb1eucUtFxBdWtuiuaV9FstL/1VUhFCGz1E42ksJIQH3x2xwlbi9z/zXqq4hhaDbczkSB/aIG
lp1c66/3rCXhWSadGd4ooP6EKc5iaMU99m3SzKDdREhwK46IUWX5JvWGBqIMEl4dE4XDRdvg9Cx2
yaP26fzgYsGb6MZimJ4XkCLqjeDlMKqPAoUkrL9oqVvqUlXA/K4mqk2LoReAFmi79/L87ZCNpAdy
3lJihw0NCtXFCGT2q7PEkws2DZY7RF2BdlYz37GRR5r5GYcNcKeEH64VoaLNvm+e2szIaTRvhC+n
4hzPDHxUMEbjTn+RzEfUClIWI3VCTCLDPRxP4UNVEvohomEir2USGGIuLY7Ln4eMpx+nlMcXd+Km
mxgVfeXdO3v18tjE/190IJEMpIHF4A3XIe8zHZ/Uw28VaucfdGUpc/ItzZc3SZmQPHAuqUnvWCPZ
IMPFJUYIUDnzXImjedrB25RIE0SWuX7pASzqIEgInRK64KzC1Av21j4cNZFUfCRmKTD4lTMPrG3F
0lY4Vpy3nxe7e75o3Qh99hV5kawmnMnse34RnYB+e5NmJ2mQEHmq9doLsYyKPnuC55puS8ooOhLd
iYP+u5K/9LkSIMegORgMBzYUQceQG6JZsrG+NkVpbrgSWFoNcedPS09LujnRq8uIQXP4hGwiC1IL
11KoF3+t06G6fWJzldfvXPE/zw1WAoJ7k7w1+14K4CYzxznWnpyh7PJSbUhRJnOwpRfYGe7nfFEa
fnpmLdb6JN3DneuB3fasSrArXT2Hrd3NbNF47LyQqba47HvEfCkbpKvZ5X7zd6676wnktwf1PUr1
YVQ1d1NUvuonii1QDjpi1NgwdvPmC7KzY0JuqtGS9wubqgyspggBDuV8y2ElOfD1BjxfFHq3H62D
6oepZcary5LUxx9flGAunyXRX10hfsLLoLndvaIyFEkld0/wn5j3nurqunWrG2SzzXz04GDT251C
sTs3NYlWVYyZEnr4aN7jgcWUb9FXum9x0jrq+2sFfRrRCq/OTktx4S3GnEfmcXbaY5a4w3gRm9a4
FMMLiWM/UgpO5gvdegky8Pp7Lw0P2VMH2gePZT3Y1BPBIH+35mlaos6xXizzZrWH/AxKhlprja++
9JvA55IF5LRw16c5GNJkFeiboXshlPNfIUiLUkt899Qpf5KFSlyl7Q36ep0SUJuisBFqllp4yDmK
GMq9HhoaIduLnLQuqHNbMsbRasHowsUwhCYcjknTXmLzf+Qipwk/dEwY/Khx0vEp9rh/qwQGTgI4
iHfZfovYrXtaqLfHk3y8BzVwuodKyU3bmpVwhyz2Md4zxTafRZ8T2qLV8XlU7yilmYc38nFaxx4n
NF80X+7T4pI+9wT897NpWRmdWKfSGdEjeirxRE8N2nInOxv24FXbVOczc4irInZIupGUldQs85jw
u8k8CJYZTXqGBUosqA/sXW9ODlvwhH9pG8jyqjnkvsSthPtrqDJ1MR/nWS2obNfvHmiqsDONMl1a
M6zS+CW5S7jE/2MR3kW7JyN2N26OJKy8PxhOnIr8vxrxxbGl58+ySc1xqeombys6IQOjTvqXDc27
6bHs7s/w1z3HroFBy9ewVR7SMrlhKLEd92nFcVHpvBYl5L3N0g/Est2qMXrUVO08eGaVugclyz0T
xNffBQoZVkeZeA0cIGII6hagFCgnpzc84TVwX7vAbl/4Ez7oSq0QrocM3dJpqJsXvkzV7qWAnQVf
PQvPxulyjCf7E6A7eYx4tHnIsdrHRIP/FYnfnG+JGweTELJJnJGLZzAVlL8nZ1xa5X7AXBGDpAjv
1d1HwC9BaqbuK0cqGwosl84awhDa5sSpF+s7KyXqT6BiIZhWYWTPPsOcAEPIlaC8ZyC+96/Rt6aT
Jv6nmiXsF8YvDnAghkVSFc9UgAoH1mnEFcomJ41YpiPAdnqrlGDdBK01URK1l47bgNsa/RkYNmMm
A0SMwZF9OsMKqtFSsEYthHp78pXr0++OY9+hHQClRrpkW9S8+8hVe4cW8qe2ckqdHBulZVIrMYAj
0GVKcB7KN94ugxLXB9+NRwXXQWobHlYNIKpWjk5lKjZOszmBZyth3490Xy4prBTnD+djONi5/yCi
D6zvef4gwbLM0gQWbb45eUzrDPcsfSTRTgc/CW1sdw70aVcMrrh7kYJyAClXKWyHsyZO1PWfdhot
Tyn6U1h8g07solbQ9f55H4RZKeq9EQWE271NrVbRmhCZK4oZyy41j7rENHWe3asBmmrTD8mCLgVU
nnCtIvgDywPP4djeJGntFDkcl0qAA7ZS9MaXHIsUwJrWrx+ByYuI+lLAQpNxbJu4zTA6VPQ0cMhM
kIJUYnmB8gQWKmMZZqcvFU3hv4pyKBdwyM6iXr/ENex9PRBKPS3USFeobAR/6uQg2X0SZt2Umt+K
kEgRRWF1FaLn/Kwq+vF+f8HqwcLvXBsBckC3ADVzt93jlKeAEKlZ9ceMzIjZuDlqBlFHr075PtrW
c+nX7jPM6B5BBRQdSWRYkl6+C6ILjLiJKC0zFDfCi1MKu/rRD8lxfm5hXzOG7dKloDtkNNs3oFD0
tVMW0esp46WhY+kRQPJXU9mdxlURmwyqP+o7TTA1q3UDCiZG8+aR/a5PDi0SzOr/UHqz0Bs4ZA/6
k41AegbZSFTnSQSkmqGgqwDkF5v0XTaN0i6a5sJ17uIRGxrEv9Hv9qEj7+hzm+DagY/FTJULwx3K
9o5yWqcVRbprL6GcyECpUeBxoNnoHPt+yZ+hkdhOJWr/4PLkeD0FaNWKXM+SrohpDqQcaEM/QLgX
liY/QJvVXs+P/0Gd+e7j4ZVHUmGuUnYsaQvKoT3QboPP7XlJjj9nbKX08xElDa/yy3BjISNdFjos
+81L8QNpwBlQNEIg4KHNRMlCr/2iN0n5sFGnwNVw6EnckE2h/3W/ops6HvYcJb5PRzjMFxKoM7k3
8NY3O7DGRIZBV8qafCtVBVtVOyn4M3IGUmMlxXg1mCBCnzPBM9fFqSkNwnDZ6kObGL7fOLiObYZ1
Ix7g9wblEts7kwCYPniCFNp94Hq3ySxJ40F6lt5YJCSXsvrHxHi062rSbC/1dYjWntPFHy/7RW+U
Jo5IIt8ci9S4Sah5erhRY4vcd9jcLbbnxw5rt87+5Tm/ciXZKJctAvBo3RUnbn2ZnFnT3kUoe1FG
rrgsUL8VvLFyrCy+BGXGrj7xuJdTsKz0VgB3p3Hh6YFL7TqZIZQzbE+SdVVD2W3nDfgFKqWLfP5k
NPIacbqwc6aJTusu3FzWRTSlcX/2eYtZOuqnNdyOeySu6sP2fBsldtdCriL/dmuySaBTuwKFVcvN
Ij0Bi1e4kifIR9q5codDPmOW9oglhrO9H9qU9nFNMP1cvkRGrORF1S2sP5c3QUjkkDdCRgcugUqe
jvnjH8W6av9c3QsZXAGB9YB5n4jQ9ieKssq0T9A7YoqpOGGM9L0luo576UF5vWYaX0ofJj/nfXry
7ePAVzrYEMta3CM6bRPeKOb+OoOu5ehdl5+UOvy/6Jmddr5Ou4YVWRLFzplAL2YRcYcmx4+sVrU+
/+BPFhjC6gyFaFV8LGGhU7IMs8ypsiMf095x8GU5hoiq9Bu8YQp7XD1/MZ+c9cZ/kJO3ohMiWBvp
UFpm2HBVCKpINY0bOUxq+GdbGgx2we/6loHbOx3WN8vxr834a5H9Oa2P8I/1c3Uvc3hxVYwBYI02
XZsPD0OrcwxPi0tH6sQgkjHPlXVtjbjCjKBBNu8Az5Ync3bsi2E0OZ8edEd7tQTfKWCQbm32RLf0
mEeSWPuHtkGoLJJFPHSIPde3TqseimLtAhNnzcmST/0V2v8nPYyZ8xEI2QjXCW06LF1IJmyt2fWV
uxTblGiqhhUcVffy5pFP1twO6s7HfxPMgnKFh50slGvHf+dhdKqmdTZizrXormc28OXU/2muoqDO
TQqly6pgP9Ucqd16s1HdleFBPCw6whuwiekRZI9ZxSNw/Hbjk3sDzgiVoJlHUF0vJZcqxpM/80HP
qLltVIilGXddCbJS1HPa9fBdbrSYMXNHqXw3AdvKxdm1gtcqHPI1zvFw7FszCo1lGFHmULlli02h
X/j7YN60kjUocweOL5fTtcPcDHlc5nUv1V/FqBlPhkcae+p89BLdmpA6WF+vdSY50ITQ5lKgYBiA
QjEmukriX2yvmmqdsVdjby/TM7Eng0DkxfehX3qrL0lwnjgRr6sQQ5hHg3Epe+cU9V2yoTT9+Y9Q
fNZvhYR32F7PF5LAiIaoySbnrsdFQMG2VuqfYc03fmnptQuZwMFQlFH+HqlRMGGYtyK5d9Sv9Doe
AAjaVQSCtVp6mR0KacXbj/6WEMOJwnPvv9XEyhY6PV9PhWMZ7o4ceYuOf0EG92IccspjAS/yrwxP
Vqo+zZgVXOwbwwesbShTK5ir5WoiOHcn4WQ5+7Q8aAnfOf1CK2SshnRTsxVDHB3Hg1mlZcH9hNL1
Tkht1CHl4q2F5uU8Tf/K8hNGXE+ad2I38Vh+v6b048R/hH+CsVa0IzFYBVpx3kREQPbjGUcBAOUH
RERNHpIWPdDmRJapz5pH9kxFNgPwbpvGzHli6kqcptVp9p726kxJNl56raond08FYlitpbzC3NoJ
bCZQmMEZVTft10a49soa81Z9IpZQge07mPT0b6i/+JKiSqTLDPrX4LWpl5+j+g9wGqS7R1ownWEi
gHnjW1so5nJh2BFhVi6DGQxXi3I0PkSGDazZcHPAgWtvojxRl1VsfwcpFjcBehoXOmXR4WKRxdJ2
SJ1a3BQGxuKLioAkt1yOgBdNaSaBQTH5WUF0d+mNPv+JT0TPhY+Cd+IE2j2Ypb7zoitzpFiB4BER
uA00GBg4c1xg+fb1xZiq0E2ufaVebPxtMQwIxbN3DKREKmK6PtQFBU8R8/hA/MItiNwU3GMyiArc
0eNUcWi4AjUNOk1kn7fiDUuH6/VHGaNLvDTvWympVI/fDZCn3zsNO7NPLqqXbpVJ/zeNIt7mzAhm
U+sqcu8NzGsgTOyoB29o5kqY11lkbHTvkBGTsaUIa2pIxqRUCc1EbnwZV03Zvnarlp2u+xWWquso
38DAiaq36IYzGEPCnF7SKz1C18qwbeeP3kWavjOv0d6CkObTFtplq4k1SYRrcqBxjnOIOJ7d3CVg
Wo1EgcHd9hR3sWHLvK3NbpQz2MEdWcAyDwFJ/6MuxeeOtsAkXqLCcVu8ywlITwL06QFulLQCj/pW
WO/yqY1xTngje1sV8ac/XKbGS2pZONn8eCzpkGQ57WdOXR0Cnq44IchNir9PpViN28g8MpuxH23a
SO4DnNKyZFl6y2XP8bUkWfMzwTcW0qSdoGzKCTGpb2qg+HOr4Wt1VNAee/KslQX3sWatIjqtsgDI
5nq/FmnkV0b32t0J+Qj1znUC2KTuf7VvwLysIgiAIVNoim0ll/9YfUKnmUgzwfEuFKXshItAgiTd
RnUFxCdo8bNzzDOpRpdWXWV4FTJRWY8GzkR3bm42hXslWkMq7XNMnPi4JMcBsjGtwBV4kvyz+RC7
4lzuWFi4bVO9c/rI5wupnCJbAk2gotI7ucj+D1COyEWE4lyNGOfXKeR1U+voILZ9kFqCbTgB8HUm
KneoqqkD5/0ioEWSPfP5ufp0BH6WIc6/IH/hG6S6OUKSaj9bRxDUFMK8jK+XFATdPtCaF4zOXWVd
jNoRahMHpKPflo+zOnFM9fAguSP8V3nsSyoqJQjOxY8ZTqZHFmsFqN5sS20a8NgxY+pTdmhlLwK/
ZvHrySPrNhiTdiBMm8WlHgY9Re8pzR3oqAUFSHLtoT8YTpjrpzWyYywANHL+TqV0T4kpeYuT5wg+
YE8CDJZAVbLmGOJ5ysR1z2aLv2dEFGjT4KLEIYV4O0XmfJMnFiVzUXEzMb2ZkFBH6basZ4laMFcX
Ac6G8fJDY2WppLxB7Bj79oOkCsI9bgh7pTr+OLh1kubyVy9IWSuqAcJd9aW28r8q5LLg46dse9hS
yRk1RmR4XNSWp/tqB1aqYfTT8PK/KG1Yr23Fuz8LEgGKJwtA9vROxxpuVpg+9U48fIgIcKW2J9vg
f+Jg9Zlux3E+EjQYtWgWrtyTXGWksQdVvrjsSlSvoNPeUEntrl15VgQHZb7zN1IKSq63Ij1uRDMm
2D4kGuCvdzI65LQctOPAgFnjuUhB6W7CFGPG6PbYUeON6Syd17PL+ZPFjcZcdQ3yzZQFXSbRj5p0
BeCz6MBRWveipOHnOJ9X2iO14iGJFIUmvbEh4Ofq9La8CtInVOo6j6WBKwNSOXFfstXpAeOQ0H7U
Lm1XZBz0NRGrmL4HGMrpZdDnNv5xm+jbWa8pVssQnYn3KXrZF9Jm8ll5BHaYu7TcWAeVX09gW9PS
35Lknai418I71oVhd9kIBLqbkvPEW5v1XJvClsejaepPnQAJRPN98JBK/iX2F9982tBr/7FbZ0ty
RZaJPgmWRgYdCZ4wcywQqmIBpk+pRTo2Pm+6arstQpcDRwbnCMvWHr7j8wkwiqWkE4MXZZcX+ajj
9hTHGFkypkBA6aJhVbF164xyeCH09ZUPIxdy5heCFomerw/kzVTbid0CdVKe/T0+bhsAUDyqgTdN
UnanDexa0uo/oee7rJV8BXZoIHtI3B65JVwtggjk9LSp8aXFOkP9hWGRBqqcaeMh3WBwsTjrUzHz
oxBe6YkFx7PautHDFANkBVNb4goKLGJanoy3UOjnkonQ8kl0uiqyAgqaTWuJmr+WyGA7KWafD2Zx
IdXE+X3MsiCQHxrZJFx/+H5+PlSYLmnUADRf9IePqaWk0mb/KX1ynM/IjFFOPUCvWsYd6Ku3ot35
oEFfmpzxKwuTh5zgpvHiZl73nsMhdUgv9AcdL+PULDHov67tbGcvNZqJG2TwfJjf6P8amseCK8Pj
8LrsVPWjzOWSXUxJEBZa9fBUV77Dwz+KWxao+RuaS385qAkhcDsszbJQgaK+B5wH/v1DirhclUmw
DijhYCpg2eqxl9eS3u7rmQWhaj7ZTKVEi92jJn9K83BZ3Vrz1oPheBHiZBVRcmRQPLYYL3HJmE6c
5PlNiSkkRIkfMwtdL5IJVCu3xE8afW+6r9Cnr61Wn+kTQ/tdskfqpeIQe1QOz/Bxol1qWMy/RLfc
QvHr1ZICEAaxng4cmnoB+1WLMkcxYH1PeSC7Xs1oe/dEDbHllnfubCG4UbfCfuBfJCcUAfzYSc6q
g1oPJRXRB0CXUghN6Wc07HPWWYXRIgQuAxnFtiHUZuqNlDcAn5Ch2N3NU+R5kUNjauzzvfGjMKdD
C6f/8JXFK2XKCYP23mV0IeDtWWKJV7+bv1Y00TwdgYHVRt4MIfW3BsguEJFNumZ4PpWfWDeVktqi
hdG/DLrLsVKZFMS6grxROkvJQv4S8sX2dXVE7ikRHNX8VPYYBwC0VvGHoFGoTHBC1oUqmPDxmN6k
QPa7yF+intxs7tu2EH+6yfsqstWAxH+S+sIeiFxT92tqi2THhoGkf5+PCrboTfIDXAIo8m0zMSif
WJhHJP6Je/Hj8MRbsZe2eK/fab9JXEego51t+/OR+seTQ/EcnogyjiL16cEB8LwI9Vz1xj/BSo4P
rF/RFeSAndUAuhwgsONm3gK0qzdFS8GSTYfu3VKlCL+cDeoJcc8rlFEElxZeYWp75MOC50WmeDgw
VWydM7BgepM0uboDeXmMCGL1erGQALSzy2crB0YnYh0Px6P17C+r++BJ3neKlS0hRw0aY0fPDDC8
dUAlVDqsiUauuM/k2QMNUawdocHlkE6BcAmP8wgB2ruvnepdCxEugY9SCchZCvla+CfdVuEHhb1h
n85POhgMb4J2aYKHS834CdtOn67MLqVb00HK3sBy2xpL4zvrefwg2kdF44lZlk8tAGsD8Qi3DuTT
ak8tbPJZZkDsQ47ctdVsmkVqvyjN3ZSgTXjxx/iq+RVeh1mv5lTcjfVcso7Zt26Wxv1hIkmYgfjn
bpZuEDzLOmrl0gGBX8lTI7CzuQIQ0CnLksEWuFEN2K7AB24bFO+k4ZvzvPA0VnT+947P5mXqdA+S
/z1K+3r9cRFeTPgudbFf4uAtoKbDtlh7qizqWMlXX+jZO2P1jwNFc6E34FYhFBWvH+ivTXQv/4oy
NwQwX2++Fkl6gFoGHghRgs2jn0t3p3DQxtfbvBgq/kBPxneajeCtXe4ahWaC9h0KS3ubF5nFydBm
V7YzthKSivKj4upJ/AuRQAX9nhKelf7zHouupzRwmC1K55f/Ybp82if9DNoRbQIdhI66Mw6FO9ey
3nw56ZdxhYMFlJCwZIvrjw0WhvBS7Mht98xSg+9FYVB6QNFpYtLoILjzWlIX77+NaoDWtBS9l/mS
o+EFoIUrbOF4bzBelHDKH80zXiZPRFrUlDCssdyUNpkJkUIs8yQyz6JkInqIBFkiqlZ/s4wTlRMf
nQ3dv3NYpdrLdoIkQw/leVriJ3mCq++Jxrhsj35nwKf05KPrbrGt42IeM7SNhX4bKq0PVTbC+m9x
I2Zpfk/75A3/T/xdRr9pis9TtxzvIbAQUkVFezzD0QJ3R67PM29I8t/IZEocryf/+4fuvMPVk1o9
jvhGDO4AaJ7CSXPqBVKIWmNcNUQKmOQ4v7uxIYlcEhw7UP0nEzXFHRUlZ0fwp2tOqf3Ejb/peLRf
IBX9OazlUC1y/Dm0ZvdQxVDgI8odZzIm7pNcD4tfitPfCkOhW9ukoG8CBlDnWn3RX9SEx2zyaxDb
KsUm2vggCQtILiveEOTNAjuLUjEvhYaxpCGgT86GvqFxQf+z7K+jM+Jd2cthb9K/qClLoVaYP4tH
bIL6gecHEIgMhRyeHSyhpCIAgB1uHm8stJ6juHfDNmZSqqbdR7EV6OhvM6zTMMabDC/3oAEi0vc1
07VCONjP5MTL4KHk6IjxITV534as8gZBT/WsEdj7HYr9smt0Osjgn2d9MXScabkbsBc3FZNuWydo
hN8ZFxdWhSTr+a2cqMS3DxCF7dXxLZ8sjII8/YW1VitXlX4vMUXZjTZMYnrKE+71Zgz8SfPZcRbD
xS+8M3R16Glqp4gtyj0DXNMaD23Q2+WvruOnBxZpM24ClQ7w9Sv9wewIbenzBTi96bnL5FOysFcR
+qZp5mcyg6ZwMHMOxh7q6zP64rdlfqecQjAiFX4LI5y2ZU9RTQPX2k6d10LioZcJ3FiZ6tignmgu
57E79fXhSksZElu3sxiAeqLm8M04tXX+pXWCsteW3iB5MH4K7w4Txhhequd5AiDeg9F7cgZ6oTCW
hfo+bg0VzxCm4QwRUyCb88evzJhCzUe9HxcKQ9JXnx3sf/XdpKoojPJ8gUl7LMHKQmOmmr9xN8Uh
8EYT/1LND3Ezei30yxqTUZpnqxAqH3gPzMI065lGKoifd0joOOlz39qW3ov/V0zzyMfWmraiuFxP
k7Lv3Mk9CdSMKowLEvw+waedz2Q5CdUEL2edkq3r97bnHLv/vKqJFggyfpyC5MNQtigBatCyUi+f
FRv1aLCzB4H/xY68fguewPd4faIEv94iK0iPNeCakAyVMm9qjVAQYP/1o4noVKQqqB6MvQksMTK/
nX/Y+klGQ4KnIqYB+q2kL6kC4ZGsePm3ZQbzMsE16oM7IpLlrujIrDoRiHC9r/KrTmFFd/lc7R93
T/+3SKAihnmPQymNwadDuNq8jVhu38dJdRHHL6bGikWiAtCCxyhWD0bYAPSfYJMx0k56LAgDLogb
7WSwuIv4o9Cx4wNXXGk33Qqea4G5el9AaGWEzaVON7mu2ZYQvMJECIGgO5b60qFm2Kof7BumpqPW
jEmvFCi/xTDJkBdIijdPyfcw+JAhZUZp9IZzH0s2wkc6kT9/SwvtR4FnQp/kTq8WPbKmZWNQpoIR
EmRmUwAQi35PkbR31mAQ+r/xJ8vn5r3iQk4IsducKtRq9P65eGWmAMbE6/IiYAiRNPyARbHv5uyr
ziPdw75qpoj/xdibsUyM98r5F9k6D/h/b2BinaeXLpPSdeyKylnC9CReBsDJFHxqI50jjb2UoYQJ
k9CwQQmF5xONscFiWytut9+Cnn7+NcQMUAIhrjkxPNUDuDItryTM+h7Nn5OlcBMrJ0M6qtvesVAj
ZGun5uj0i9BpYHpqiPPsvsb4muE6MoqQQaLDX7np9CPI0OXvH2ZGUDhiTTKdVWYsD+4rFdonZx/o
QDGYqBPlt2ETaaSwyT8H9mZrMCxv1XULolsP3XfGSpwaiIXBXTsGokl+BwXPOPkqV4hBdFGL5G/C
sR1oPgdtdEBEo0GxqoyyvPVjvCBgJT4mrlbDnomQVdUkxl8+Arh/4G7bgZnYwlMEmha3jm6UHupA
l+a4lwwfNpyOecAkHJVsDXxAJ/Dody4dyjettdj6ZOsh+1Zp2K7awJvFc4rg3s+w+e4buavYg9fP
Ae9wlmvxRCjC714yqw4QbHhXsWkrAul4VoafxBXE3NsavtCzSxdtro7NKUNyBmIBvic1JdYdE48Q
lSMVoX+GvZA3MYsV+GqmmF9kUbF5bdhlIW52rUUIAqUvnFAplTI3u37UsaGlCOwxEuaxe/8WBOui
gHowMd7bqfA9eMFrofzsaU48wNUSPeg09F8oViOTsGwgGn9tzaEvbHjrHDTieacUCAAd6Ksp6lJV
UCsNb6CTQXe7PiJxtyys5bKU3DgJpnqvs6QdeF84QrDH6zKxCcxtsl2AE2GcKAgOH4MV4nLTCo2j
7od2COXkkZw/U9Yx4ZK7c+1U3QBEm/EwCyUzWUvl9csQpF6IYwThFExwbIcWX0Od3vLo7dAH74Hg
Zz7egGaDVpxTn4epk9MCQGbmwi93NSEYGnU5mRxrYKG0I7MrsCoVk+xn/sL7tj/xlDkSm7PfLC4j
Gu3Ms+T5vooDLiIFY1yyNTDPIniwVsy3JtIUEUItqAMvVvGmOSwDR6ARwACgnoJgsh3aC7h+nwXX
hr9TcNUA4KyES27jwRD3MHo/eGGQiFf0Z99g4CWqoI38O3TeeCsN7XQsp0osP3qstnKbDX08duti
aT3QSjv4JNxpJ0rV3fq+bAX44a8+1aFH5YfHYW4MomKxWr92IMhdvpOSzRsVu5OSYs+poWPeU85U
XhkTI1ulHcWvzRvqIRFeeDabJQY6Phv7hIj4xC35FX2hsGN1llbVSAfnCD9LGXN2y8XRiAvsQ6PH
zioU3gXj503JjZLaz22qHIW20IzzWYV8HS2MJIJ0fjI4XQxojb6IC5O28XKEhza71hDee9GP1kiJ
vDppeA5fsXjV850ceUBsX7O5JjJQShxS29UgPOJKH1pXrriQRBbBA7dr27CZnxYeQhkJ1UhHzukD
ARxboC3t3OyJN+xSVnzAT7CPZsFozCBG+rBxqYVquSEiYnNEfKvRsEVLmDX537V4bsD4NTgoX+hk
UIXISvcv2eHzjG1szRtOLJjdoD8nWv3c/1/81/1RIyHCd0l8mKhvwpOz3/uUCzPSmE1nTJG/9o+K
KEaQSb2gonfozWaoenY23tOn9SsOUHCzpSZ0hRH2HoVjgPVTXZjhqWF1KVYJpZzyiLvgEPq4Bg1N
czfvumHgvMkHmJrlksAp2Am7F5aal6WYVvtTj3uu/WROsV5/hy5I8UJPLETnRqqh9rsGyy25glYq
Twtk/3hhxmdJjbsw4NhmOrtyO9wqF5mJcVnuwZ84/tY43YskBLABMuTze8tSp8/5xq25PVCpEWDG
o4A0lrVml5tC5wIwuL3HfuGqtjA9eEw9P9bJOk3wbVGh9YzlrIZsGKBI5rxuL+QogpiMPgSqTdxt
vRHfQ1n4v/D1B9noTliNgWb8BMAQ9unNf5WxRXdSJttVDz9m/zPPMIaqG/+WOtodWDvIl4kXy5aF
E0eAb5SxHxUypYVob6YcGJ2ayR7efiICSrs7PuEdoMXHE1Tn+iXQXkyhvMTz73kTFktBQeIkp+qB
q+wEkrdp2fHuZPu6BmleoJ2BtvoSE9TSzNpFa95/UJDDEoIOn/TYJ63G5DUxSQei1y8pL2OIGl5E
jgcnI5MZB1uj+Z4e3tKjeb7cHkf7Da/LZRwvR4L5gMP8zkDGIIHL734SK3bQCGLI4Zuxib+UXwdC
3Tkp/X8wgQ6Qaosw3qx8lCjv1JISt1pxk4uUU+jhmiQCnoR+mYkTdnpWUbSEvuKH/SSTJ92RkS1i
Ha20+ued7l/mBgKTwRf0J4cMtbQ+CDccyD2DJ6mOx73oJvC0Uo3JhtMwMkBerIsfTdQqQcXDBjwl
65CDZvTFJoD2kWjHyOECrZwKDJMryEqGMHxnlNnOudYvof5JZ72FHn66et8DmRyi1ZeXpS6CqbcI
FTBDuB6fe1v8Hb2nsVDmJo3hylGHNIFWNTd0GnmQHGlthHz7gXciyU/vHTeKeAuFvx3tV3M1o4+q
5bDQSLyh+Onfmq6UR+u58Pci4qJVHxedyys45t0EUknBPuQ1UPRI/GNZZ85TcmWQKtXXMHQ3xetb
XgUK5CQt7QD1otDHkoM5nEB18a0hNoSXIc4bq5brh/FC3h1PY6zdIrg0cOdxSf6ikM8T9cWro5v7
UwTmlIVGIwbF3Y9o1YC4XYdfEdla35TOoFUbLAK/zyRC7HzB4nLPla5rdwHkCB4l2floH47ncAwn
d0DXRzXVWo3zmVlHI7H1xv7OW/jaq/lj9pm8mVw6cusr4VftcHQhj8N1ERScJVQGiJcsSJ1mch4M
z1Y9o7rY2/6E6wIciUwB0DbvUyRChnwBidXuZyjryPuNREG3l8rocTKJVvVG62X2+zgNxn/4+wDQ
c6YBugmJ+ARrF/+YknoGeNnh9e2GhJ23FQiAH9yLRCoRlUv+MdEwD0gZsmkjnv1dTyFCEVo/Wb5j
MKTOaeL+pGzhkcUwb9d/cMFa7n0Qvwd2ze+jC/ApSOsoBrHYWoJugOGTkl39Qyj7dRgp9yCyUPzA
H8ChpamhsYVjPS0lNOn9QG7ivH4LHlpT97e1JlROWPdy713wvjBxKFglCGy1ZXPVBnr0Z4LxfIdm
b4FIkpS5EMjW7Rp0g4jdJt6itM8CpijsYrSgHGs0xQOMKhCOwFSOuNgS80rK7KfymVym9zRfy0Qs
1DDQIMRO1rBVdRIcs5QowYBg3NvcpJF/HtKw4u21/e8XBQH0JkL9VhrCIokvsHrabApZAJZJAugi
yk3DwiKImONg0nu/DNOkCWYwJRVtqC/Yy8UXhNgpjOZr1Ebte/wGi+ZE6q/i4yOu6wY4yqmPqAJo
W7t1YEoNqs65+RiNImXlRBf/G3HkY1hkxLNQRkDm11e0ePQggEjHn7nW0oahuq7XcZMldzJ1TJE+
p/fsmZACvbE4gcSQ66eOuhmI+YzlysM3e8+ObaTXMtjQKGkjUlo4HPlEx9lF+HbGS/Lt7+zmMUON
aOduNIutS1BfOVicIEqIy2W1vSNewrlagzgQ5jFyRCK0CmcNvGoltrtI9AgYZdxOoZS/BUtDt3Un
nfI9nXQO4cPb5OHHlcKqjSQllmNw7O6Sn61INuU7n2E28Lz5vl1yaQ8FSZHlay3jGnAGzF2fx6QU
xjFB4Mc9iPJgft0neITxbXkoHtdFHnZLHGxAvi7EaF8oUF+etEaU6F0GG+Io2Aou6K629udtgTX5
HYZ5kTsoLP4Z/5w+VlEi9EJgOBi7iIWCsBXfB2ae4/IwvUAKaS6LKNB7wJcm7M80TYc38gEFacPv
g73Cxqu2jX3oozZAIBWV7qkNdd0Cj9EyzrT5ktwmcLD4kxcn3cr+2uUazOi7V3Px/tr3yis3cwUh
zBCD+oiiATyrWxRoNP/3pBGloMQxAvXIFPGwMyPONZjOoIGG3k7tcmQ61WxNx1lHqDIuLvkGFYpG
DOx0i2Qg18oWiYtFfhTBZJQVptbfArSl4eSYCLE5oT26zy7AEeO0bxvSbL36ZgPnRtycO00wffyJ
xPTHpi6kjStxhR4ZaSuEZxB/IYiioOMHSnnpEkMWQuMttNT3q6vZWf0/vkBL4LLm8Wh+WLR2nc1Z
TFXwDlfgVUI6FmFAgm1lVzjzGn1O09w3TIccGBL/UhTKIjQ9+989ezay5exf55zASKxtgFYt51Jj
IfMXbrPke4lz9sEw0BvpuMIaHelBdaWzOMRA0CQnAlIUD9fsUgclYJoDeLm0+dQ0kND88/I6G8lW
QskJ5vkpm4R7/FZuItmjg6q7gFWnhwwTSDpj1vljU9bUlcdYbP8LreJQPHp1cuxXOFWlAdbLdMMm
rUBLgN16CUSdAuCZAkY+07B5MDemhcHbNSPW5tzXeBrAI5Y9kPQoyipAbH4mNtFT2hOyiLaaQFYM
ccxw4M2d0+qJQ8OndbxWI8kyuO+KPU+56ibTCmk7kSO30SKljmCxngeJ2LQh7NkUnNcxu7tRu8j4
2C+g2g8GuBC1764OYGuYfS+Yv24Zue/+XHsCPtqi62YEVDbG6YXSMYUpHKsLVSgDc+N9qWyIG466
d7+593tGwM/Z+iNH7US+bW2GWrhozZ3u00kQX80FTtB1hhen15EipNBot3bcTgSb9zc1FGOso7+0
X7yhpDibYOrWpISkglh0LVY9mYUdufhdXbLscJjN4axJ+zDySJh2Ux7BoOfAruTq7AGzlCo1nTak
VdjwRTfrOVYklrn+vwWmbGZ5q82stw6Cno7VY4feGbODHs4bXOux82xhXvgp8VRRvBfFBD/oiexq
dqAvpWWa6mzp3D5+q1BV0G2fAsm303cq/MtW7D7+MydoSLWplfJDtgS5wEhixdOgDtv44PNaLvhB
aAAMGFqAjp+5HGdBWqz8JuaOScYLJSfaE/4aj/v0ydScHHM+AmZiy4n8PCSv7PkRPPsRslXYLmFp
LYKxmuxgY4gu5mT8MR2XCCBhOsC5U30wqiC7d+vY4R2Q2TzWJMZNQQm9h8WHo+toeZurI5j+T4Dy
U527LosBUELI+S78alm02LOPy0XcnXuRkZiFMdDu6ow8iHoF0XSx0JA2WvYw1NEEegvYtIBFIRyM
Lg7JXi92I73+GBEt7M1thFbJiFBFE0P/qMoCKc6anLSKO6GT4ITruE10DL9VQEbp5dXHJL5o3OZJ
JRM0V/vi0joccdAVEJpCX6CwaT9kABsbHJP3NuNPwbdoh6rztU+cjxYl84NnSefzMMJSt7RsMsVY
IR82p48Zp7fcT5Y7UmBo3bQ31CY/SruIrOO8qzCop6EmoPBgDaUTCAFJmQNTYHw6kRP8Oh6/87Ka
5QdKdH2+WHVXZsKOCkeNXb2/sRbr3uXr16CkjIWFeFzlQ+Y9SECPF7dHQCQwAkivX/fyJu1ygY/r
/O5qWvmJJXGT6g0z6LsAbBuS0wB6H0dFmnChAPtF6SCpXWkGu/XS0iFO7qEifGdW6gzGGudpfSe0
LvQ/4UwvIOKM6B9KoRVXFo5g0oC4cB5rfqDjDMzsjaLppLGVIP/FD+1hGq0dI6QMh3WwXrTvwIsA
2Eu7kAFYILCTiFhPQtGQCIoX0eUw/GoaPcblA+QGEhnrL+E/uWw3xRXHMMmrkk2KY9UOnklb7zkc
26GJqXAFF4U82Kdq/mwu+sBHjZZ9Tk/0ocrWsLBqiO+Q9GcUnn08UnvtrxY36YJhONDBVcxNLILU
qxmW8aEoGAiwo0m1Fs4sG4ZG5d/T6j6nsN92GLCxtAp2QRol6mp/y2y9HZkWymsH08wL3yqOCI0O
tlqxnjbKuNORCkWGOzjHWkBo57G6Ep0wofeK/w3EPQxN6SOvCb0R0xBWd21cQodnyucM/odF6WeP
fezeHZsee9sZMniVzWsiZw489iwr0gR6jv7dBu/f1kjdwT3OcTQp1pQCT2Z8MHqQRLTkrYOmuO1b
U9tTAhQWEBKHie9Wjr98iTu3NTaSlO6U/71DNL4r0bNS05Id5MNI3IUtAId0MJfnxq56VzYdFK+3
vIKcEm06t5tHx3LsBHal7QLtr3yIg9kR7ZUAJ1p+QMiQ989z56npUtzAaWNEV17jK4Pup8o39cgs
Avp4WHlSJqsF/HptI+FFL0WaHAB5YvKu7r6OiLsFpsznLyy8JVCrrhmGvg2RXN5x3AeFcIAEUAgz
ih+k0MWuP/rQaki59cvOedafH51djA/T0MkJO/0dVADyM7dthdlcdMvT0Kfx6QiKLgidKS/j2wiY
r6Kr8ocoEElYma1oyI931hSZPikFektbLEonGJIbeiuGuaKJ8rK20pqTLW2iR6ZywtsV3NLXrDMQ
pZET0PnxRh5QW0N15RsR6wvOieW0C3HkH1rinmjIrQFTYcRS448RGuqeuLPOJCUbJrv7PwDsy477
GZa0KNEWe2gmuciLmNVqb9Zc4g0bzlu4mocPzqjUHzlLGdIPKd8LoTg4vNA4z5lz/UdipxXnilQ7
YDB+DvK5BKgzmmtYsd1+HZjt+E8KLSUHFItCLES1oRMkEdSvxjHoVEgOTJT+LF9lNvo3YNKjyRLK
XShjJs/DoROTwDszZNRDkPtKAudvtNIau3Sg9rBccn2flaEgPZOluFI1lHcg3efx9SS9yYngJwJZ
NuPb6QlTUow5xIGk5/rRv6kyHs76jnBxoVCbETJ2gXv9Kxirlhu29noSY5jovdNt5qFOD4obSiCd
xKscH+slYcgXBeFsZit4BWkHJe9khj2t2P5/omtQMnXk50ALTuD5Z7cAonqjIJ9ca/Z4ShDxH2EL
BgFN+TcfES3nu4IWKm3c/tMbGKS5Q57BUssYsPY0wU2ekFCimiCClDocuV18tbB8gJ84GUy/RHzg
1cX4/EF3yK1C6pWzCXVUsG99hdCv2jYGy749Ik7CRE2shhdsQg816H1CA601+p/U8FWKGdOayDNU
zHxBKo7DEUkPo1xZQvfc8lvNHoSSSZg8wZEaxeETgLECs4FxL30boysUTLq/vsLspVv6OfOqVKGP
T5/zXQFSNFwyhyQAZp+28hH186no7P90cm6Bc32WvL4jg97XkVwuR0l40LViXby38uzfJJZ8NfR2
ScB5Gto5ixHOerXXIsaM0x6sdTQ4GHJSqLjngFQYbLwaJ4tZhJV4EHAWIoLhXfZLUu3uk+CO0iiZ
fui/8yl5Wj1cAfEHxshbhL+Hod3P9qGmEHKoNB45+V3QydUV70bCD9ajNpjHyi4RzUwQJ+LzT4Qp
KMP/uQJJsWl+NID//mI3R6JdlVyJMgqCoa+oEP07EQRFa/P3dt0nOVIAYsmb3uKCaiiI4fgVpPq2
CDapj9yh6Virza0e5q3pJ68cHa2DHgAIJGJdoxI3++L7mVlNJo1z/MfAH1a1Lvvi0ee6J/fV3xTg
0EG4psnkBs7/VsFjzUO8CmEPSzXJL8Bc++MBXoAZ8bZT7yKY9aa2Jx4SaGaulkQgQFKuh3mD/rcW
OdBQbHzW5tjiAqgIYTSai7B5HGZkDJGXH94jtyyv3PEJT3+FbHGYBMKHA05VrJMbwJx0nON5Yxue
XiP7gjSWgtb7Y1n5b9e63xI81VC5GCVIi/qLybZEhofKNRMtRhS1c/AyLInsVZIH/Xd67fjjvH4I
JXDHjpk0BS3jGyjwED68vcyB8D2omZ6Tv6j0Tr45u00y3XzpdTi5Mq8uovrgCXa1KWBYw5zixXzf
PzGKXjfnk/nW3vVk9NQncO5GB0ip8aBRGd18zVKbuNuP79Zpzt4gtXPgLNDn6vZy5FNw/5FcTtxk
SmzRUhfePF9fDD0zbf5KieBm5luY5Fh2MUCNCaTNKf00gOVqg7YxbkTLZ5AAvWnRiwy+ZOoJp9OD
sC3GDXmXedOvqUxX4skYdDWAa3jEH1XZ19zyN8s6ySKBYGEX4dUla+42mX5ncCbU/zyno4QN/z95
wMAfDtPRhef1UDm7PsokzLc4GmE9wFiLryYjEHIDktOVUDrWbOi+znYgPHxI/AN9P38NacT0VR5C
UssTIIZfoUXkLLmT/v+fOsea5mulISMLfhnPgeB0gAcPEJtsyEpFlJ2pYmQ/ZIREPm28Y8fMrdoV
DCeCoHw4n5hOdzkCBBbuQ2KXpvMUvKLTWVwzOxNWmzm/lnVBmkHE6rVY8kwZaZJg31rdEXw0mVe1
XKZF1FO2MfauqeKweWqe4mUgeNS986Kaqv44gPlFj45VOz55ag/Rhh6b67krNdmT3sb0USQDQizD
yvtRJSTa/CMUmt1KqCObB9Ofc9TKFB16QTymDjMkVS6TdvTtpyqMn6x4jzTerQQOnb86ORrcbmSx
86HVx96/RkBwhMxbnPWSWdRpXyPlnh9T0QsIQEw8WuNlT3b8oL/PYb1ePnQOIhu9jCVIxKCnuIj5
uT/Cnzo9a3cv4Ea3dTw2q0wDrZEGN1tZ4iGoI3XhSheQxXdKca8U69JasQ6bi+qN2hQSjSUfn9Sa
luhsnqVUNlKi58w6xvDyhw7yT4Rq1QPxp2rl739cAmVbljNmwW6nrExUDcSGdCxgyCt3DcFTdkLy
8KyqChwE/zueJQmlXuyTm7+0DlxHh5i6hEJCTr5RJt1a8+p6gjKj/MVr519CyD07yPrmaGMgEjsJ
VZamqi1+Akfrhc0Re5TrPj8QsQuLSn4bxhePGhjivNxGGf+HEWALG88EjCjxyAPoUc29gIqK1P3O
PtX/qqwzKSqBfMrXgEGt6Th/aRJ505xz3KpYMy/FAH8l/oAB3x0hHiwal9InXS66JMG3N15Lb/Xm
RufBSN71kul2aLnr4QbfWxVpW7brwc6uKO1RUc5S8NTwBjfTtb2sA2zeW9WPbAhKnBH24txOl1Jw
yWzAcKj7zbTkC1fMdnq48b0pQneI1YbQYqmt+531xiZ+kAFFQQTTd094ypdbStsmtdARiDlMz3IO
EkBhNYC3nO934ch4Y5MxjLvnlf4WxwRAcg0mUlmFYLadYyBFzGp9ihWZfQWtUDa7SFRode07w1Vv
wvYSWHilGA2egHvjF3AYFywte6dIz0k34tmIg6yZMuSpFD+JmlGt7jn9hGcbWUCEy4Q1Muk764fy
94LPcsAvIMfFFyJkVkhRdGPJpNU+3IgtWI9Mh32b8swDfooYhZqRQxkUBcYpDgXZVmPnTCym5X2l
FX6l+joXFDsntZ6o3XBkhzydi1wYar3hUZoacm0l9dK+J6hX9kMtRdf27uCdPtcaa15eCTCPXd6J
jlCuQv/kXOXQUJlobj9ICwSeiKtJ2XL197HQqLk5PXlKWbIVebxUmUnOXXjCCap5FCJccAaM3ErZ
ZMylEegsRg2xKcHCSg+OajgU6xay9P2vNL+2gfhJap4c5D5e2NbCzPbcoU35T5Be2Ppl0gNvwMcq
rNLQVFfHLH259lUyxQGiZKaLRn/MlDCPgH8bEBv0IKOwxCn5eyKhVQWDr5eaBD8B9YlzkHUAzrZ2
hsDO0rIoZbCSkaygbGJnJGaF+ORAyoIDzCrViQ5oNwcHTxici5bKZFZU5ANKOKVW2nnxDw575BrD
ov3PryFQJarFihjHLmDUZDUZPs2lHfdsBwaZndzbnEdsveWF9kz8bQPcRnMxvFvqRMg9+Eb8lgN+
EtibHiAcsGOXNaqRt0ttXpqmY73MNYTK9+S3ctHYKsUqmfxjUJ+wvznD4yyaQDmkhvL+bDN3ULYq
U9wgB2f6yy5kz3w3gpqZAjGOQjXE0J+gTB/7UFL+jHQKcpg3FE8ijmzJjWfUlBVTh8SM69vB/cF6
EsjeV0F+Wc6l9uEsB9LmY3JqitDdmxDPaGDzmYG9XB19crEpZcQ3o+pyvHcTp7X/SCxZ+G1/CoDJ
2XNFHu5v2GEWmRuq+CUDl8HtUCzLmSZLhGd2odkL6rMGtp0OuVQ2z50FtK9TkUJCpW5h2VBmTM/O
F6tzg3pPDZJhQ0u9RwZgbe2C25y19dE+SmAAs/WMFk88jBPaKLp1i/lxijXldSa23ct04JLO8wa9
mjztW3Krib4cvGmrMUAlHK0yCxTZ4CmHH8NXb2Jr9jK/ku2T96bMbi2ETxqoY+VwxaUTbRiaPA8K
cVHnph/TNb0bUGhE8g+qpSkxf1sOoOBNVyXJvv8rxhZu77LbtYV3OJ+WkEw2oZ6uA5OWxivh4dKw
GSTUTihBOb3Oiye8a+IRX7e7YE9/nfMFFxq/j8rJFSNTQx4NZhORXxVptCrlLNEO4fLHRvlpjoFK
NW/UstHm1+SaOMUR5Nt8OWQkmfkpX4+aelk96SOaI/hozk/ibrVpb6IGO/D6PLeIQT5nAS+piHle
pEyq/rQMJLoVjnhvHZlhDkfm6P8AjW/ey2ojdWtweP8vyoBO8ZnupasG7DjhuRIpZV0gst2/mzed
ixTLgEjeoxdNNdK96oPCR0diu5PUmX99VRIp2vWPBxx6xUyQhMVOeYWZkj48IlQmSR5UNUKi0o6q
B5ezokDY/5adqPB0Czh4Rx1aUXINhxN5jShQrc+dToDokF/IqWmNHwj4m3P7qVtVABAz6z+h6Nn8
m/4m4dwI5iguhv4A3v7FnUnP/TSCGvqL64F+hntGnQrNtBCDy7iZVMfE8ILu9ufhzaGnO3NJexFi
42LdHp6Mcf5pTjZoOTImyMMlKUrLav0s+Wy8cxXb7olZAbq3cYhik5sYF3iNLdQrVav5fCPP+uE3
PNHsa7YsxSi5OWvOfxQo1DyxBeAT1rhPPpHRhjb9invWlbt6rMUmClH/cwIpkMbLHdvH3j999Tde
8GTFr5fW7kxUnc6JeJ6bgfXJFiRktgvbr6DKeAkjvntIKFt93rykOlnEW+7km1WQ2COd8mDnyYE/
VxDVUEs6/hixVOBf3CKsaxiW0H/buDrpuZcln1hYij1s7LIWM2eoF2Js1Y1yft0QsoHFfzvYlQuP
4ThsFqn8cCzY7xsg3S3xYU+a+W3nU2qcQpLCOTIVHtTBTvqKJZzG59xiBtchdwRPgF2Xgqwkzb9b
h1Ndsnw2r6kYlkJemD5iPWP2ag+WZlh5mfFKCIXsPNWLhMitQYyxAZCXZElHBy7MohVh1E4ywXnW
HjXw0UoRo4tuI64YfzCFdmhOBi8aLLga7ne04qlKpzI/ypa2B6G01XDpv9gN+TH7dU8JaVcNE6MF
23HTwdlTK9QyBWTdUf1YqW4GBfgi3TNOq8FK+TfTfbBM/yjc6vhecyhPPWj56tdyEldy5aGb3sjD
bHqtA15eQCaNzHvkkkrrfhfvUjGUZbfRYk6Lqq1nJMDHsk2nVUSV6xylmlAKpYtE7Rlyt7IEBhnF
ExT0sQz8DLt6+/oDD7jdM6UzjSJdWRsv2ux3mmtauNW1c1xVuAIdOBsXtrQQD+7lmFCYp5S7nA2E
pAUERKQOjqQumXVDdMZ+2uE7dOofiz06f5ZjtKsHH1zEvnXe6NOAqv5EWJUM2Fmz1Zhk/Xs8ZBQz
aqG5ru87rYXq7doEXvpaZNagtzG+gjvBJEHfHGmcGJvQ2V1XiDqzUEFhpgvYdBC/7AVD8aoMn1z3
mAU8npwrEDOuBdNVdirp0MoridEVcCILvSwOnF56539B2E3//UFb06FwIhqa3umbPNEKGb3CEWtx
vpmJGcBUfCA6cBQJjVQKWYKVdlSUUPXRHWk1fEAsaO/vniz6XXZV3d2buPdo7ERmiMsUx847lNDI
Z7+KMVh9ojMjpKa5jEJ9dndcOsyeygEXcbbSDtqa8tY1/ppmUjvw8low9odmsV91DD0p8knNWw7o
Q6bRYYDs8AsC+JxqKTuuZ+9f0EEY1huj2p70O25EkW/ZMe0OLHK5R7wbPGRgdq5bkb+hNe3aBIJk
AvlnjK1WcBWTJVC0KBUPulbCSqeTRRqcbs5meepCeENmlG8V28FdoJXyALekJNUIVSkq+K0Ygs1m
ggsvHV1UQ18v8pOehn9THZs2Kmn+bV3bMWPR0MaY3dB7YpmuMo9mIcQQyfC5U6fLT1wxW1MvTe7H
XjyfdLvVaFlvzgjEVWzqHnafff4WRMaW5dEmQzog3NqI+5/5P9Bz34trFIAxkIhKKyAYZ9jK4vfc
t2vT7LER9+H2lWvButVk8JnjJlA3FS0vT/ZmXS9OADuWuNPdS9C3+nyDbgDLDp7C5E4pHEMX0DeF
mP70H4tU6JDUjPt+20rCSaPmOCH5xt6fLz2/20EeT771HvKbIX0XwS7rnMA+Xdo5/TiiPOao04Sa
wdtTQlgqpOCOoE7eny+NELAzfYai9Er1+bR6vg/q/G5dhkMrSatpmX2cTTE2zD1d0qI/0+sLYjBD
gWFmQq2IhfdY1Jn7wHsaPV3d72oA577vWEp5SEF1tMStdAyp+UKdiTOnIyMmDsK6nzg4IuCKfE2W
mlaOz64KY1eNVZKrCCSykbuMlRwLM4Zqx6sMs2JIlCvMTplDliCgh4Gqs0ZrmKMhQw9ppwySBBQU
k9ZEVJMfvKrkLbG8Ui53E5czmhhApRM/iSfQhJrcKYC9dmMhPzDqllC5d6jK25HY3i4YJBqSKaMR
9dzbR87+PGtV3xYI3o+M+0/WsstHGN7QTdddgTT426K1Xv1ch+HxnB8fXdYrJXQhmTEN868SiTEx
C540PoVBakzbr9CM2AzNK0pX+aN2QDc43oF0q1+soY4WCjLd7rlZI1yD5b6Wyd8IvjUh2BRR9Kxh
1yTtEE8wMtzlrZvFLjdqCIB4fVkjH3DF3vQ0looXlYi+AMmUXJdT8CUmyufs6fmhbbtivas6l2Bf
wXFQrvmtBEwfRKnh8EXci3+3riXlZG8rLfsFqMaj8jk6TpJmagwPZ0HDXLWDvpCIiZHuDgojZ3tz
Ikon9IVdRYIWWSwH1JjwVBHoLz4MTqE/7xa80biHKLKnaViuqbFkLzV7zcWNHVkZxXgKgGc0xnJQ
MgbVLbpQ8C1OnA2Fd4PZ+Eie+I8hOfHv8AK40SkpsSNBgTDPt50zJ9w+vB33riKAxU88YzXfKDW+
pqlyiutNiKoOJZU4EidoRhveYv/qTjFfdLv27zHoYdnlyhwc/i3aPDuyoZkWz+FRORHDlQu4MGt6
hAxiFAhC0higCIfl17UHxj5vXZaV0/wZ74wPhaV+Z0CkBSOf0WhF+SqtRjUYL0RCWIXFmQ5d+7V1
HX7z0j5nF2OXGIeDAh8Ik5/XYFOGEg7RcHWS/ZKsPgpEa5RWEVwB+xHgq1X7M5WxJlHABHxs6+8s
ABdwKJ/ufabeBgWk6xG9uNpILXd3Z1ao7+mxRjH737Nvf9I1uW/pVi+eKJ5Vhwes6olVJL0Cj2qy
FAOZJU81u4V9SqlZOtbOexa47qwzuTqYR9MWa6PNKGNk0hvUR2RdH50Sd9/p89addnxkx3YasXMB
oSGDy5pdiwwDM8f1Cxdgc82D7jqp/26ClmfrgU5nt6EIv0jIqeC+v271ey4i3dZFiBhwQhQoSPkB
nqolnhqkMJhvGu/S2lL7rv2kNx/hs9CSNyrbkQ55JFRyqfUEY3cAQQWh7BHo4NrPWSRcImUgsbpy
WZfLgvePpV/sM11YSURutrq9uLt+uZ5qCqa6ZHUj6ssyA/YzTtezoKOEW9R4GJZ0Kllye4Yu/cgW
R6ZGbOsPBVDPLSuikH/lSs7fi0bawxq1X3MhQmunGqMne+nlIiD1bXfueWuwIjiQe82UYMdO57qt
XdP0IElej1nqOIPDczlChtuiANuDS9syKBrS1wTqzcFkbMFFbXykitDz/0Qr+ZUGJr5BEHiuhVXz
Qjy+gJn7PIOuqly2Nyxg6rtziF7G2VbhA5hhjaXsAeDQpKdlQAShfg5pprv53KP8dz28nS3PCvHT
b/cFddCENf5D5JVRSDiYpR2qnnAgUkQFPs2oEhRD2+R6oKpSPO6ykqqb6pDtTDStKtsIxeVSJrwx
FrcLGFSTzQ5e2C0CTwHg5Hm2lfb63M+qWGzLidTdGSdGJgV2GMbznrYQpVpXYWQT0ysXHzEWH/TD
oXU4/UTRflBvrVNUBL6zyfLtCojSl9qWU7UY6Oc9tHlH+yFGyJh7PhyAUQ0lvoQIi1/NH1CbxN9J
dPbFgpAca1Kn9HaEb2ZnSUIXvY735gATWj9c3bAKD+RTl1Y3EjkD3hxzt3JHocmc+OArMBqn6SKZ
bfj9hhdYKkLv0s4pVoq7sbRlt19mwxyWT17KMC5vhW8pyVQLnnBg50H/5lyhbJRAqv/vTr3/MTBD
sdzfS9nqszmjYaqEaai3r9dHSLY5lJhs0WXP1bh0bV5g38nx+3wKaooLf9Ax9E6bQRMJ1f2quHBj
Y7OtQIVO/FTaebWqdUMErQr7tguEnPIJuCGgi/OFJkJ2IF+/LgdnBv2LgtqBZl+Aw+7xY6jeEqX0
RcZMuo51D/eG2yrWS0G6rKo/gnx4X15MsqK6RDAbRQVs8LBrkzISXOt2kmQWTVF7iqKxymPj0Xcu
/YCfU5qW4LchO3Cr8rIlNdet7hphnSSpg7oOebkWyJFCNGPjwZQk32dbJczyrGU3O9hKol1BtiAQ
eFct5CjwyszZqUCwA4h+iW29PxeuAdVDa4c3NfvQ8rQcesf2g8wpFWeodPpWC+XZ7rplslkmOX8q
ke+ra63q3xLuQu61+hGzelO8DvKG2/H+Dp351zcMbrH59ncTheXPsM6nobbJKrnst1aXfdm9LA2J
4yiPOKuiXpOTX9dkUDmW/i5Gd8LPZi+EV7VPgb6if1affTdsDopXUw+0uaQQtbxydDFONo2wKXRz
9X5hFoOybRki0jDDaZIwkyW3efexFkcKlB2HJfZhbXlyc6mXdO1Ag6qQ9HUY6uB9isPsHif1osTr
YVgJXC1LdtP+ePNClOJxSvpZPeQYqaLT11kyB1aHD25fk1gGxZgGUJmDrNQYpZEZRTYZRZMR9alz
4f9KbsBc2pE+gLQ8lv8QnFjVhUX5vZsanggCUsrsgB+lYuL/vJUJCJLJRl5ffyffvpU3nsQOALF3
wp6xojdSE5nwDtKleIFw7OeTlMqeehDuk0Add3OxlTQlVHltiTPcgjLn9XJgC9IWiWchxSqEwWB0
h+YYPAS07+Q8v+wkwVqBJXw2VQyY4QDXT//fG937snPstxN+kKoQu+P72sVTg/z0MxyULf4NjRqW
dSuhyF5sry0e5QJVkhCzt+gg46C3qfGVD0t48p7teWGz3bIRlZovDdjnr5iyWt8im5ajZo/nBj2D
D0QlzcSoqCncP11Ns1hLBTv4zfzfRBjx5WmMQvmATak/nFeoFfdwlPoYK/FK0qHfXMkMsq89l73O
S/amopu6OeVGOQEE1W0FzFwbjS9xvA8Lx0fK7eEQRJJiQah6XSeZy9TMiN86gAhaXvXjVsLaOOxh
Klgz2sIkLnTXPort2AMbt2xS9jNiVTvUp+LoJ8+ytNvFjqsjFIAh7AEGyHRl+FObaNxqRSOza91+
zOYDVlf5YHn6nc+i/kKblHGQS7L+kVpZd6JVN+QuxPTZrEVvR4t4E6CEPaw8a09yCaaTTdrBt2+P
bTAVcBwoGUfKygUFm9Tu9cRnvhhQHCXlbHdDh8+VRJutB2aMSms1X7rSHaDd+7sqOf32DMypUhzl
NR9E6Bf4m8V4Mi+zFwaK7s3NS0KXG0iH8vzFDKsd/8FvFYmGNjwIp1eqE6O6NsUm2yjbBlNMyB4s
DqLfTyXcNRWfz6zrdFx7Svm1MLfnabr5fL3BC3oYrOxt9f6wDgKSk71vkRGTkgpdfncVZhIgu7gY
spSAzIYIeK3wKQAfK43TAgfmZnJJKBTr2ahnRS/2LTY9A4Ns5FK/Sk+Rw4fGYWXdsWRQE8aMZgX4
8fVaFt3ggMqR3hd0PK2yBl7Yi/MsGC5QerUTml4+J9xV/x03HCHNn9y21OEcyPiadHprKDkfeTdV
lvBbH8T1WDB5flwc+cdNy1lDGi0Z4eEkXDzK98qpoz5m+T8BtuPle1j6dBXONAY1XEoF9+iD5OkP
tDH2HfitgHRPmKu7P8GZe5Ie/O/XLphuRxBJUGrU0fSWEFetibtSW03oX+iGwSv1bo8+vmbT4GZP
ouWof9ssz9Pmq0m3nqz9wJ23JQ+Omzx9tT7rZu6AS58D/5uXW1I8GcP7P/kXnxNsF0E1pJrVXsG0
1fSvi38bqGHrq//3qkfWmoyAgkXuCBHRZXbENZT4qHCQKADvRGgp9h6FzvigiPGTzt/2I57eRVay
RZ1eP5waAxCZhz0BQ+WeGvhiZRpgAv9igzKDOB3C5pI5n7s0sOgKIPUjbQ/u0kzZr4uYxiPwBOil
zWC7QhXNb9cw2+sEVBmd28FduIKEt3Lio/t6FkfIcYHKb6gxOzFAOTP54e3BHG5yX935/FYywz5I
eYNbU2+44548cZXLSjddQu/gj+InloviGj0L1n+jznfTRXjYrVG7hi3nrFpFLVe047GCBeifrOBL
i5EFelFUyv7PH5RXlhVJAw49z7e5QG3bpfSGRLBno+N7Mz0tLd6ZikNzfAZEi2hE/wi2k58tBHHN
f+zUbI5qPyBj9D3qT1gBA4Os4JCpGrWjAYuYypNUldC5bm7zuixkWfWORcBHEYGRNt1b4JbKEzEx
aJQ077EHHV5puRU93Br4/FtBGIhlHrkPzSFubcJrRtEZq/WgkGcVYaPgwJSihmpsWbmlIebScpK8
5I6ki4w3wv72Gl4zwy7zRu9ONwNX+WDNaAWeo6CX+nFxQZHfoeA0UEakw3WZKskoE48DrTkkJZGP
rKg1ubGRmStf696WurImJ/rM37XFEoj3/b56Mldvmk1M+GLuZPlt4syHpJ4C/laNWHFFrte1sarO
yAEtfd2tbCK9sJ2wyrwK0vZHP95unAJu+rfC0EMVgGnIT86PscyKp2JtNd3q11mXOEaIJLX92Jss
D7N+EKCTyJtnL02ctBrhpSBm3j+gnC3up6PfxDga1/o8AQGHQgBW3oB0oe4FhnOTG/n5/wAX616y
wVWVQjkK8s2w6iDO3rKRshNJKFQuKAklB0kgftmGxtHtXom5zrgl5jGuxNT6wxkNowwO4Va1eEVu
h+QhaXXxMRxQi7wbrXpjc65oLKlkCrtwiGVkTuHXsGWbVnyk4YNg8z+eKRSqz7ReqSSCBrLFxY0q
Si04iUksD8rdh3rYeY+G1YtvZbkbfXy03PaPadVWBapLhwwiv1BcgeBy3yiUpDMCGt0Ggg+OYJdy
+Ogm67t/Z3+E5S2lTNkhhZsBQuqnzCwQ84g6p+csk28SZQ+S/DVoPd0yoK0zMWVBGmtS3VfJvfbD
7r5jgllDPkm9XNuS2vdbWOzmnQdENduvos6YMa/CsaFtNf+xo1QqFS29HMlfxvZpK/cHmURxGtDI
Db6AIqqbsL0QlAFOM6E1iPLVTbm/saxHasIdFjlct47SWWELAklJpXSLmYAxqZo1SLaPLmty16vV
Rw2+sRNl4aB65ZSfyH3Z0FWKjCFFjcI4RKN3bnagPEzmbL+BPrtF19WXo1+Pd9zVzteMuEzu0IFX
COWrLircDj4Ngf+ZaNUWRKHnNdHjfYtUp6Dw6diVNG2gVhQ/xa9M7miemGTaKrZX5Fr6maoePGiK
Y10OYtvv+NUmiRmgWQjBIqcuoyAmxVyWBq+lB7sFcBHhjwAQG5gIy/OmfyZ/QFImwP/AK57KuY7I
PnIykblqwcBH3VHC1CO51AXdZTpuhO4rm6wrddeMJm8edLM1B6Ly/XeQR82RNBra2HNdTVaSZWPt
jUFC4HollOniWP8XORWIK/At7gcm249mZPNGOCun4HkymB7XEcHVQ3CTmyPpvO202xawKGSt8Kg/
Nrf1qMbTy6KNJDlKZyCqk2ep49wGv+lnFs6dah2dIlFwqmZWZ3edSLP9vvJ0Jmdaig25UM+jQsfd
49SvTszYnsZPJ70V3xfjqod2rHpClBxAFzJeGTIbWhNXi+7VSSD/QXOTTV+G9EZybU0p2NCGtC0G
C1eBFI6GhNNOfxgHer32rJtGyUH+Dmw5vs6yXVVHEVUyyF/G6HkwtslzeA5qfltsjYTBFc+559nT
U86NahJnstnZ6WeCgQO2Ap5nR0A+D13qzdblLtTZ0Po1TygkZxsz02hK2fS+Iyv4KA6PQk2EMou4
sfrlMnfdowSzZ5pwzgD6D0GjVG/9WQ1nLWyp5q2x2Lga4laoQmvDHG4ysUQPmTycaXb73yM71BEU
VxaZXHQVruWuCZOePZ5XFs7LEso4gaWiDoIq1p0+a14yHMkkSLPCeljLEgsF1KbVgtEGOltvZ+C1
pcCMUjx8eQqY4wc1vM+7SCKKOKnfA65qJ9YNqUOdEXxn0YdyrVDVndLIJJXlPloObKfrZU/zOExa
y7H5htn8JUdCyvqA0/VOstsptV0XeSW0Rn9dua/PfSKMAfGjkTvyArgTu+ngyQH/Dm4BSKlHt+4Q
FpRMRh7354U/fsP//r2iQLd4qrevQhqikUjgesNmYXI3GpkLvPiAmVw9jeQ4Tm9+Oy4NHXL/FBWw
A+nlofyil42yajolvUK86qPeEoPopACjqKrjLbLXyHKaRLKFSzrQ+VS9XYcbt0wqOlpFRRPLSwnn
yCiu0hUlXP9pt06c0GvkSGaPwlG4utdADAP7jWBoGBz0PgSyZABc1jE4iOHZcZgZIvq2F7Z3ZEI8
Uucbgk4ObqtpQUXKp86eVZj/X5FjY4nus5Uhejlkut2pM4PxXoDn21qWdx6oOflFBpx8hyY4w9wm
CcKa5KSMdpwnSSeJ1WXSegOJi59habn/8QylqlbhVb5JOWJdCy+QvKn+s2YP2L2wzytchLoM9VJU
ZXoUthHRo4IVJPigdOPWYUiXr08biWYN2osQF6tEiEIhgyZ6EKMv40CB38NK09ljvRSCTn3sc6aA
EtlvXwcqn5Vs4UXV23otsGt2wq7Spr4hZQbPxkZef09KNC3FCBAvgaSF+JT8FlCa98oK3eqCFIU/
Nzk3JWNTZrs7N+WrzGkVJoYVET5WJMyShh5ejrSuT5L8q8CUM4tz21p1orAEQtIw75qdHCjHbTZQ
azTbF/aaU6F8vXHO40DkuW/itIx/LR2cWWUsaTznJXxQbiEIyMtWlxSBdKYv7sqhJ3l47movW18c
QrX/rl/CqlnF83jvvdDZ7DuBpBinG9u0lJGx7+VQEW3cOT2B7G8hSkkj9iGB9f/Y0QsoGjwx0LPG
49eNSbWqEjL+qKfCw4whMBgru/8dRBGWMtPYw1zTwUViYK5frKmFSPo71KgNXJplIAT4NAXHKsWa
PQzwuT6OsF5XYGZbbf0sb+w6FTMGPjsRrhVaTK8BqNNAFGMRcTSVNbm/isnQr02u5Ri/aoiDINsT
LCeokGko7PGVHc5tc7QWKezAkLL9surnvUsZ2FrR362EJ0xcJYjHCCCmq+ZGoZ/M64ECWng2dCrh
Bvee+o0bJ7qYAiLR+Twv4sEB1NBIH5bnEbUE465VBy5r+qEENkJknY5nwecSMiRj/PcYfv6kJ7sE
bpvUvRXSjEC4IAS2dVA8Nlnlig/55rAoOps7aE4H6qwhGpIuMUGn/bfG3obvJnKE/yiQ6o47iP1/
j7Qtfm1R6nwflAWzT+/4fxOti9c+hsI5kHuec4ILLIQNku1PtXurPZcRqcEUkHYWgI1fVNgWR9Pu
TYX8FtBjkg1a2iUaDIyQnkks4wFf98O59JwCW8C1/p60OgX8qOZFpcuX0+MqFme889216451yWHF
rbkKObtzDetZ+Dfqog5/D2P02ZR/pc5fZQ/lL3ZbNyQ3roeyb5Ly7IzBnqd8d2xhJaXlhiTddBha
x4h+FdrIxvGGSpmjuREpTbvGPdpnt1tCKH3kFMTt7Zy+D7GoMfInXx4u2vqhqSIzYGA4qax6bvoF
rOD7waplC+FGqYLC2mxvfvtBC399OLhDB/Es/Sged5bx/k4jCP/hfMkqsP0ShLRImIohO9oOzTnE
TSTJwOFgbUN2bnYmY8cv5xZnKpmZMZA4DdOQ4N0mJgIFYa5QSILBEXSae3Bq8CBqeFwlKrIk/vlu
AMb55YdIk9EGd6jD1BCFPHz+zRgx80EzF33SK8uwaUOzuhgB56jkOde8yLZEqQdv94lMfRzN9erS
sutfVQpmqnJXeNaTSqBjEmM1Iq20XxR+PENvrx5zyxmekRt0fDg8g6VqTGRmhdJ5G5CLMbJ0Kfoq
cee4pwf4dBeAmqUjNMqye8+f81rHt3+trVDiw/gXhdWIVPgyJD4AfVoEoj9GXhZGbhkIWA2Px0No
Zra8bxEqX9ZDy9K9x+PhvQBwZ50arR7UbPRNX7lVg3svkNeHHpPaYCn8uV4gTqB9Le3WoN9U5gxr
ygZG6Hn6c8Rybpb+Zbvms1YD90x01+oM0l8yVqO1Ayt3PuQ2bhX6eG4adyvyoqcaHrRhT8q51CGZ
IKuPaOuLQ4lgb0EEs/KLz7EE1hKnMiJSoRBSCQ1qAITFTU+b09UwJLVA1/scXjTh8RcL7tis1YeY
KmcZlLfMKaZS56PedB2yajIdAmwDIDdccoWKJ/LAu/8GGmcrUgCrodmMipm9cV0wxqNxxwY/LWPB
oO8O8GTkOJZUcFAKkldLplhwqDrzU+ZYQiKZ4y4CdtZdB+pb6YhdsUkBOrU5QDbo+FFw9jQ9K1i4
HiwBdOVB35bjPlns6nYmc58JxQ2sw/maorBwCrQWlXV4R3zxZ56oju7zE1zVcBoqQskBvP57dxK3
n91RmubALwSuQ6/1yKNHyRSzPjrsVaH52FcgdbxRrnbtaZ/uJBcg/i8QduQ8xbBNl3HjfTs9oYCK
X+d1I4/E4xFGZO0TRljYKuRWZepx9pCBXy3hKYhmzXZZDIP48TmABw+JTl7x/mHVwBJKkYnCgar4
UYMm+gbdTP4/lNivYqECymLZSmWWh4LbPHmHcLC22sENppazqWwbZ05WmH/zgPPwA8JDta35nOdN
RXCUX50AY0Vpz5UC/MgfND1KhqToBT0iIN3eSZ0z4/sMZTjg8xvzvGINSFeZVU98wtRp/O1pjRqH
ZV/QsnWHg1NGloKwuPcvbJFowVDZYHlZNue9LzO47VD/0qTwUTpEBeoyb9nPa4i+1sI9dETEvUgk
XaiIobSLfDxA0s3vCZOXd+yqQr734DvK3Pz1S4k9Azbjon/p0vLxFRiOHhmRjrunZpiYEZ5Y0sgb
WQK7/Kcbkimhx5vzWREBLWgqxdwSL4EsJXT6igivrq5TawQur9WL6+NTkOj6hH0K3JGi4DthjksP
LcGRcDkbXs2DRKiPhkqIpE63ORkLpkhaTkxl8oC0TIcYKK04O5PnQshhONFevSgiWkPH/g/+QCB7
etzi2JrAZek+uAWMo7GOiYLEwMXfvPJryW0Do2HCNFtTGmUqjNpUP+u68iBsW9MubFaTaAGWT0MT
izbw9Sowbd0FFGN26nBLzFhmeaKkNXLRnFUKDeylyLq5603Zt0NZQd3kATgKVFoh7WfVcfGQfggg
WE2px2drA32jfNmt7jmItvKx6/Wo3jFrFqchID36zPCVaOileK4rVNVCUkQNW7jw8he1mtKS/vTt
MJ1sIQBCcOasQEXRLrYOWwILakSEuK+l2JxM+i6PSgt13LJnpY0B65AoMu7iC5jro+g3ESn1oT4f
XGt3n2RpecT9vSeGai/zpBr6lpBC9CN0HFx5xoKbasv/dHFfHZGlzcN/jk77Do8TGAHG3DeOQnSG
ACAnNu9r8RbiQrnr72nvtmA7yVGTl1uQaxrP38b+GUT/wY/TRYOdciMnXNnIr0VnMgqLxMoBpXs6
1L3+jKQ6vL+ntgnpS+Nw5RKxXQ/FtJlWh2lqM4ZA0L1iDEpBKweWLQUWvXuzspvw5ix50L2sCaSH
1RJ9OxIQurRktZB77UC9yVcg2dTqCX6wly3hDo1LaWMIbH6iT2zucgzizD27W1JJZXHhR1Fhz9dn
6M8m8ZKsy4JoBMDXxg7g+UomTZZqMApt/ywh5XgXDaGhDFDEiklKJi5EihHS/6SHKnoyOrFZSdcg
2qgkt1I4/kEmPPqlwTr/C+vZYa9FoGll1+Yv5UKfuM/qdhi/daqRuS3k7iLiI2DryZiK+cjhVR0w
bt5KlZELGi8hw3Fe7NEf1J7byaMPjUjRdfazD36dFExWqJcOTmsEKHtNwUdFw7PiFbINnRxq6DUw
9z0rX4e/vHkoJ52AD238mx4wJYwVJnSCEqlbc6OYrLz+GZVAONDjpkaV42kSAMyfFJAQGb7xSRLO
i39Wb/jOdpI+QxOWPWx0Wgkg6as0/kCyjCVI+Yb36+aD2D3099+YMnUoO55EMqYF99f2PDfOCtDv
UImDmJu2fXQI0B5zqPxDIkiFIwrmkt17ENpI+LXoOY4EIP/q00meE0cGgScel8jvTl2j4vKvukfV
MLW55dz0dFCNpTJtXAH7nwvTZzGP9iCA3dEWkQHuowAJFp9GEVdIC72c0zrFs00TsBxhn3KToBZs
2g/pDLKUb28LJK8FmDrpGHd/rVI10zfTYlbiXxYElS/g1+Xdcs2+LYo1zo0zeuO9SuH0S/Z0sdQQ
Yo0iP20C3XFATr4fgxChjGh6fR8jZqyJ6LO5nG9PejrBJDNAI8YjP2tsUdHDSWYPN4klzcL3rCuK
SBe2y/nmaEbCFVceboTs5CafTqttxg98jkcxUKBMDMaB25dhBs74N8sR7dvSAoJhJQFMlhnfyARo
Pr9YtjfNzeOysogLNfqcJfmaOv3OjAG55337X91BWtP05cRZaG9a0URsdwrF5euJppx8TbdxUVZX
XZ6pKmqPufbthWUKEQQDwv+9A6vx9PZHlwlRYNqq1nzJ9fv1kwwjAeKMiddhKux/L7VaVhQZ3xEi
xw5hc1YLAB/nC7GY8GLrOpf5iiC+Rq40OvnY/KG5jzYAWlRdURO4EXL0JuQ81waTbnpTmAmDgRWf
kNICgp3GKwgbpjn3A6h2RkY7/QRHRDHFcCpNRej4QIB8yQiqUI5/G5jQ/+/7Dr2NJuvGXZiP7rNb
oXcQLFtlVg5MxmP32X08qB7QQJdbbHe6vm35gr1Zy8i+adFi+SKjEkwcNlEuCsyCeXPSMNBoPd4S
qwXA5331LC/p/l+KyxVdmqStbfXzEIpCiBsZLAJV3z56LMOJHxEZf+XfqKT9NuJa3Qx0xYl5fDTj
MAints3vzNylpUXoFtZDoTMqnXUvwWtKleko2FUZSkD0NF13Pg2WXtin4+ps7M0QM2k/F89d/IZM
LFfxEaI05aREZwhWureaIHTRGHnrrFuJ716k8ZTjQKqOiqVZacN/qCqFuus90rgoP+oxH8BGN7y6
i/zhNM43WLqKtViMfqxBQCD5EqwBiy6zCTPtXzfByN/nG5uBybibD7Y4g8phIwnh+uFqEMClBSJg
9BG5Czvb+sKA6ZqLNS6nK62gQAItjU19U/I4wjyEN3tL5wr9TSTVemN1K4HkP7jpF4dMNpxcYkVy
1D0lPunK377EkaSxDCEFLdrGBuSK/0nt2DDPlV4cNHRARilguHrop5M6n0FiCCfGcO0halvIIRuT
6oGBOaGTQ7kDGyFE9ufsRiWBDNdbz1elpn6mxNxt+RUB/cmgf11UAE9bazpzaDvLLfOSV07OgwzU
MvyryXNKdtYgV5pMIiRgNRlDVRDJfj3aQDefA9xToJG94l2xDLRcg8qrr/+6dlt9i+hX7Jnh5hQe
W1UuMi7MFHnk/v2eyJQM47DLkNAFToo/PMfitrNma9cbfJnPw2vf8ThFD1E7ikZZTrsbFqVi0D+u
X/gpvIpv++oraugpymu5g02cuM9efASLebHTzAbc0o5ybniNbpc5uhYF39vWhovGopaJXhYINE5p
mV28Lk4HdjZgxPX3+CqSf59nRyUh4dphRZGmu5OQjIIdinvjoGIdz2s+aYrrT7MOTAghrEsr4sw0
9nsOfUUvp+drhgiXN0m+1NZbpSPMoCz7QfF+d+S9aOxALhuzCU9VsA6vty0uE4fU1jv2uD2NS1aU
dtPRuXE10x7+KTCF14eIvPt6UzpkN+gHQFDJc9kXQ4PULF/h1ogeYHZzwH8/jVnb9sukgJgYnJ4E
ZhG5WX+dAbz7alIkmKhy7WiF/0a4m4WOfCT5hILkNhuCd2DOd7QX9KsRxL60aM7RqLrC8HBh07FI
PwOabOvIbsPqNcAmdovdwqnRC67/Wr3YCxGBTHticqeblYxWs5c50u/MbocgnHr3TcE0rHVK75EH
l2I8nw3HUp62xISCrY0ZSl18qm7DXZcG7mDoj2hIUbXepZqK1W8VJrzGhzxGQO8Txq+dQ9sWtoQv
nsvek/t7j/f3yPsod9uxgw7VJ8Dsl2RwEgqyPRa8eAeywC6sw/6lC+bgxMQqzxsWwi8Q1gqGcFki
fYmMWkyjp5i3cKhe9i/B4dj4qOjjhFVk0ugTkEyT4SPoOhRwjbVYIkxPGh1L1jJnoKX7lNZBey9S
XAjsxz8Ih751YPBqASKEN56tArjb01jZ+kF7R5tgf+CAdNyLfIyZsgUk20hGuDnzbBoQVRcAaZbB
jJNoiXXfx8HbvTy46YCaq+xc7lh7Zl1Apn+LIL0cG27UXwvUOXUcFHF5LCm0dI2G+6ibE2zwMftq
sPYVNzNlWV6MwPQcaIWu7JxZr97wFtHY3oxqQyOclTB1+AmQ9YRTfwymt9sLXKF5eimGMw0mLe22
kIzmrbd+5M1+gU0g9zlT6bDMhDPSxlcHBpqlOC3cOOLba1GkbrU6Bg6lnr97pjr8qO5Mic+QKHmz
RTMJUUCRHdl+fdB3E2bmurdGtjMkstc3i++TivPFsDQheNOpgFiiPlGr4+sSocAdotJpXX3xIBBH
esmX7V0bx771mwAEr8v1bj7rvH/2hNOECV9QJl0U4LUx+GZ5f4S9WJ9WXH3/3nvP4HlpDZotYhBk
kSmFC0kTb9wBs8TnZVTG1e9IOAYVG/QEDCvv6CW7ArLPX2eLLjZHIMRSKeaGYKvrkrggdW5ftaZ6
EmOIUdS/KDUj/TNHStmmVnvz2PWLk7Kzc/f95nsaUHJ/R5y8xUXVcTqIMvR6ARfiV3haOx3FmFzL
DsTWnRpjWmPZRUPhwGE8oMblahcfngyKCSItxdizijVX4eV60af8LiCeYRLPZlZ58cqqv6ohAxsS
vaWjDhpNQjqY3il8Ich0a4G9U0w4rVfeuYldUbWJHxvRTQMPPXbExviWMESOn8RmtFKU4Zqv4s8Y
uJKCxL56UpYWRqUfxmePvR9ON7pnFEnq4xLduE130hn8Zr0T62pWBHp4YGPJCBf+LK9JU8tjp66p
lxsnDuw82cgFUKsphcoH3ypIH2AOdLaLxWw/MY3Qw+qiA3rDw+bu5nbX/Hy4RpeWiuhnZ0VcrsQR
REvzkomtiSV6od6imDawu4/bM8t0ahp/VLa3Kkrly4dfJWfXx5KI77mi4UeKR9YYgcjg7L2uPyfO
JBmr5RZy+Iqiqkfw++geSfLVOM+7iUy9Ln1qD6+gNi0MYt3EZdptMYOxQASTTXjUx3hb0q2y/bEO
yW60+NaHrjm1GdNdbpHYcqr5dMBaUWx++10QBkeiSP4hw+DaZ+NwqWbTbFVkwEAXkyz6/HtdxbxU
5Lli7o27DaxLNjHf2b+NahiotDxU//WnGXIFs+MuofmiMZOVbkcPMcSxIGFJktsNYhbLcE9HioLJ
rwGA8Vkpl4q3P6AqgGYVMJ2w0YtcV+DZvNpVl4gQp8fvkroUxI09QhgxCNPFSyzVTsV4+0X+pZCd
bDOAUb5MVJebE/SAPXiS94JQp6O3Nbs2dIqhGAcbXTDhux9duPsvh0zdex1IEDn207/HbcOohdcD
cLbgj+0y5D7oJ5KWQJ0MG5XyAyKyoxFmi9Rey/3L/gDpWDZ3f6IV97MlDFYcJ//0LBLcW935osBz
ixmzmn7dyy0mzWTtFZkKAq2hzH0KV6ro8AF4+o3pgWVAnRrs7owx8NWmOweeC+BUukkvmIqTmuwD
eu+DGhrZ3rtlHvLfEKgVLn5ke4fCiDzUne20JEm8ErZryyQgKVkxxc8g8OBTbb/BM7aPfNBgOGm6
a4JAfzipXXFA/kIdNkFeWOHrN7NxueJ3WkKbPreP/8jnsv//m8HTvTO87gBOM/xDYyWuE3hqE0tO
G/QntyXrC2y/wDIfrKuxZMcWSK1abhcuFuKq9mFmQ06BK6mzGl1CaD+407xEMIVElExCmUcw7oX9
7iIvx4lXylnz0TjhNg1aEddAZMXE1gzINNg586BzL0f28P1GCJXIlJr6Fo69uFEGxrShwn06wlHQ
/JeFMhJfM9F1eC8TxTiJarhsK0qsJY/krds91YAgcRCjz0bOG6z4rAH/HltvjiP3jFJP5WJSGcHC
m2YeyOm9lj+mPsx/M/mn0x5+2O7OPwXLV/5BgexDz7fANwjOzgLoto+UARYI26hehVJgzMsYnEGg
e9EWQIQxKNbbrXtKMLwgqrEq/5+5SNtGjs20z2jszN6zt67dPPQykgMeqUI5tOuY90anlbxKCLm/
ReVRCISVukVV673QnaOmpxZtZHwM0QiCrt2jzRoE+r0onFFtH4V01bcYeYqNKAONQyht4rz6gsl1
6UNtkSi9lV0WfCMfeEP8cV0z6ya4K9XnF2wRrraSfAx04nMqQpzUhwfp0nXCDwOPHwOIZw6gmRGq
0D57rm+g5yBIGTwVSpvgnaVOnpNHB2MpRRF7CSvZMuD1P5QkJUo2nrCRscbG7+WrsSZh3KBcDLuE
L1LdvyHvxO+PCbthWG7RGP8AJ55JfHYqvSnD/RDptTv/GuAT/+WkLjcYsTtnv3lsas68ydPkqUJT
sHrOokNfLS3jkyGmsqvgpsN4t3pHVwVQwKHTsnAwaGuOu/aMu4dNCb/olJveJ8NY+FGg6Cyhim7x
6zh7+L1ch19JvLVT0wZv9wiJzqV/p1SC8W+x2OxWLfg9/bMOl1lUn+kEN2DPWNzXzv2QKknX227+
dfHmgl622vPfad4khZd397pivWN3LaJQ29rwThsbr+1By+QnhLzcI+7yfR5ZLxiInG4SbFPOCCYU
jCwxkiHFT3lAFgwplNg2tU7OG3ygQM6FUgQ3qXTnE9HOLLgLPhHHgxtdFVdRGeR2Vl3AaewiRPMh
3hCTukwl+cXgZNg11UNXASz5KU2S4iN56E51u+JYJSw9H0v2LSR2mod4s5phWjs1tZBA8z/d6OMz
3fJcE/94k6HDm3GQqsevWIlfF/dn2okl5NuWee4mJ3JmQgXIGzsWY/zTpYLPMCmmLo5NyXg9mASy
QTVTcaIz8fhWinbNSi0PNONT5Nug7wusvkXX9I3MiIBRHAbBFFtAl5YngSvqonEqnC7SJqVudn97
L5Z5ZikELM3SOrApqJcQ1abZBbWfPBtbzC1y/mehbq2gJ8kWeDe/6O8cjvP1KT+3H2lgOeSoXBkI
fsni3OaKgR2i4QES7NeLaoBm3ijbgZh2GgCr4cPkiGVn2FoMyfXgOCbGs4DO5OrTydXUERLenRE9
/5ulk6PukuE2/LYr5PnGaJ5A0cOekRamuQ2ApoFucYAcZ4HFLMJTKP6/PHgXo+VUUmOqOWBDVg==
`protect end_protected

