
	// Symmetric encryption; lambda = 128
	localparam				IVEntropyWidth =	64, // TODO rename either EnableIV or IVEntropyWidth
	           				AESWidth =			128
