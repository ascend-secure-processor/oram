`ifndef _AES_H_
	`define _AES_H_
	parameter					IVEntropyWidth =	64,
	           					AESWidth =			128,
                                AESDelay = 			12 // TODO make this a function of the memory clock / AES clock
`endif