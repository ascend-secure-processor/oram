

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
btBp7uJIJc23c8c2NiYvs+4ogx1UOm/KTe20ZKzqKWRh04jaU1yZooKOyNXrEi0VxyoIMUEgYMVO
01IlcwjH+Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y2Ep1DWEddpf32haYR5DVY1EkiH0kJUDFm8jWU1ekkljialzV8OFrzrbGY8sXiH6+o6BRjVfJNuf
kvrSPrDuXiw50EIAdduC5ZLfiuSdsxYM/m3lE9um3ITt3Gg0CnM1QXZkzKKkgRX3U09Nvxr6rG5u
N3YJfgeZKjfBhyaTf+w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k7YVQg9tdz1tsz7KOSJ9JM/tE+jcWUWidSE7NTVyltqrLB+S3IcZaE200UI7XiyGWTk57ezUrd5t
HtLTRULcbqReIzsovp7RR+/uTJ+rdpclYznCdm9+HM7uRhcozIRvamidRZBndVlkUxps+IOFiHfh
HYJFwMkH9HNFiIowtwllEVDJpfW5zpAx22JkdZpT+3nzs2BljTao/D0qDViqCHTuUuXq5E1oG6hA
92jY7mYimYfu5+eVe5sC+iEhS7G9/ehXcTKaQSGfFDHt0tyGupu7cy0YxFbAguU8307mhxREfiNJ
TOYBGReMmRA3YxDz2KKPjZIHEtGGTrb5ZztDcQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t+B3e/sHBFsIBKWLnr/k+sXqoBpVvoem/HIUo1UCMeqxRKOyUU5uZgx01WUuJZevEmGClB0kUE6w
onluoVqBfU2tpcIEsYo6RpxmyX9783b67c5b8lih2u4rbfsQcWQCcuRjnTXxsnsSS/ur0youXI2Z
7RHSQTOZispTBxyt/iY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iAJxXwAkKuHyQfPW7jLsYa7WLRlZmkvl8M/kULbBuAJNjlDv//QIzuYS9RR58RTgmSTjFxbLEKCJ
XUHXyK4FhgkL8bYWPmQNX156O+Xhpc++EoaHcWjk73k/UvudYlqq1Cwus9CIS9NTUTuDB3/YORp/
askwFhr2icWLst73FEm51zRac4f4WqIa0XkGulkUZzXM8kyZ1RLIdEAFfxxcsaZALqDauH9Fzxj6
zEkUAmaJCEveGEBWnoULewySDXRwRt2byU/8b8EJQiZLkGRgTYpdLrIkKSpaPB83fhR24RZWwDJH
5EXkNccZkLCugdrfeViFe1tMI/JmmrJYzMlYHQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6224)
`protect data_block
HLd44yXTHk1IVPnH1pNSqyaUoOpCTdvL6cnY+yOJWeb6nDfGv+/CgydM5k2CyStNelh4atc1U0Pu
WT0P7WzFAzq9JzwwBPWTryMc20vvPP0SgI/wislprPqEVnaxwL6IHIkD7AGU74uaD/P4Me7INg3b
SxQAjWpxGHNElUG/BvMQFyYDK/8wH6MrliCkdr8BttBj6NCE0vlFgE0Hqt90NGNnDgdY4OixSjvU
yImfOEorr19kxo9dQfRJOLjdK1zY1SsoG2A6mn354YBDGgl6IUmeZ8ybe7i7OR+P0jD6t27Iv2w4
NE88QJ48GZCTj7546az58fFVt6Bf+gUimoEJ5ZK/cinVw52P/KqDy2lZ+ukEgnO6bYbiJq14Hdem
fz1WgqxWMN+D+CacAf70oFpybWizwZUIBkEdIJ5V80twOmZ0gJiVZ+ST8wAEzyS9gXWrLPHpwTfk
ABLMAB6V5iqIXetqlM1x2jr07H6e9u76C3mVmEMNVAYRY6eIiOuoG/9OmF4yrLtVF8KOX7WE4a2f
NyPVQaagqiAfLji2IVrpfEqdzgfx5/JbPm0f++BYc/npHRlYmodOcGdEX0Zq15XcVl8VfXWTtbDc
zGjSc3BFNs/9D/LRkgJNGB/fiOqtvp8klV8zHE4cC393QxROhoTtKgT9XK9z6qdZkKtlRWr+v1W4
6ZYhFBxopT33LHS5ywEk/1Y5ghlnHOCHmmXUuq4aEsPj88X406/AxWsNJhfWdifFoMuMkO1zCdxh
RiGcuBvOzOQCDj1wJU/myeE0gfuq7eX5/4HZxFZv4v511w9hz6cb8lyqFsVDWyaS61RLgbVMg6pR
b4sNK/pj17Fd/ETF3/XWlRLHsXy1fqfU9xEEhpmwHSq6Iu9NTOJ8jHJmn+ncIwAHYZlvA+yvOgmK
6aIo45kG+4/NmdXHLgaiRRuidFU9Gy+QYfM+gkEp4cqdNRzxSX7YRwZZY7eBfp4F7gXFfNKyEzD1
hQrSCDUi1U4TwxjM9hPKg9skaVb9lVlMUexjNRD3ok3AxwTymaPBmJnz/mIym9ghWOwiyR9WnVmc
VNhltSkjIOA/Ec3Nbz6upVihJ+bf20x8K7JjbBAEXMGjzKxUbKefHaBomDBfNIglstjYn0WKGmvk
9H2CEe3KFJxmOBW3m1BG3zCd9OykNo1iUkuLY43FBY79P8IYWUnqe0okHgxROgNh9+96E4X6XLFZ
67HCdiN56J/95D1GX//0ZIlLELaQT2VpH7AOoabOj6HrPU9dYikUIBN2OcVg0VW0WIKKzRozEe/P
OxmrAwafV93sb5YzlvtM8jCTyR8RBVAe0ETsqzSoo15aWAZ1Fp2qM9rBVs2CT1s9JoQWDdOKJDKa
BaEW00tDVghnNJn0uThRJEIWMlxodUk8T79ktEMPZUK1IclhV/9f0hVlBX6UP0S2ywmevpoLwbvU
ll4zFqNMuMXa0VFrQR/QBKMUUqZtTmjTU9RRp3dlHCJcWT0bPynaPCRi/aXgxlwGSo0EBw9a6CT6
dDYoKZjFYLBFVKK7B3f3XARXCmgabdTF9eHYf1ESvj6l0tdTmNGQuhZHrWJJfce/0HwKBcM2EVa7
nXnJqm8bqLRTL1UKTIIJmoxYEdXhhp6l6HoTuaRH5BTSEvmDS/kuNfxN300soCILnPqJ453+3HuP
C+GLTaDOIYVrnyZ/ufTN13tToPj/Ta5+xB6UkcUHjmutqtM+88cDgeoOktj89xgvXrW6IcVb2F+I
eFtjBmyaAk72dJTCwO1SCRJWgQw8bOJcpOd/bhT0ROKHuBzJ+vwlhw4ERwlTU8w7BqcI66zhHAC0
jINewFtwuivXxjMH5LpKNfZG3GkrWSgneWrDw3udmgi3W7dO8U3frtnRP20B7qWoOd+3JWde2/zX
U0BpFUf/rTDU6xo9chmbTcWuDurG8H00qAyOON0Jetj5h6dVTnu50ZAnXxKWG98P4K+4oe7Q9jsH
Hu88A4Gj+Wigq4szp2Dl5849/yig0Fty4TgtNvqySFI/1QQYQG6bb0byyxLIH8ccVba8uLExuAoB
VjIrx6fBiuNmLIacBYxjG3w/mLd/LlBEuET9xYuomTbXSOKMQSWxnWFCCJPVXDMLkZsEQQ9lFZKM
7UsE5wNxY1jhA8mHXYipasLi8C2p5CHOMuWFvCaVDSSUYfoR6xqko+0b+wLr0ypoeDjDfUVxqKwy
GUlmD/Ru4H5fvnxJ/HHTxMzsQmAd9qeaCs+9mvM7Mv4oQzgHdnBwtOaB2cthclOMPoJLRvN/gxpQ
IGV2koh4HAnVDBHuiw37PwaER7ue6nsT6PlSh+NfSS0VS4zsgXRMT0BypQZXVtwdjMy4iWotHy88
5RCU+b/MGfeGInIKJo0mxT2KIpQ87bkwQYyo6ukD4oLu3JszaBYsrUSczDEn+HpaAJvPX6iQ+GBw
bczXKKBwEZWLoc3e2NHEm7f5DkbETWI6slAsoSsOTNJZlOKuBM6VNW0FC42RkLairNCPdcagtJWM
2zB33nn34OAPgqfipkfelFu9/zJIaJIs4B1zt5BdaJv+uN+RH43L/L3dZnD/5ALbeHPXQGJsEN54
8vNujh3QsvNvsjk3OJ1Uxsv5oDZ1slYSexkG3Oxegcxz1HQ8XGRX69WrCMfuRbCOHk6c5uFn6fU1
EiqD3xSMpy5pys1aOxVhNyTAbw7goB+CGQ1yNtRzY/ESlKlY9Pp6+HfH2sruOQA4k1qr/RSaT7fp
/OJFC2SpEXtjv8h1RuVyk0JnzENBRSyOc2tZ0PTVF1Y2jvX6tPIt7GLzdjdR2OdkO5S07Iem90Sw
3CFIhCyg4R3OYGbZTUk82ZorSrQKRrWlBwX2Q4IJcsaBZlwRPnFTVaxyTyG8MRQQxYoxvkL5g3ka
6YaJcoCGWygitaeZkoc1Ej+DwdafZxXYcd35jayy21ksZ7yCbHNbBHojkelX3KoUJYbh5ulzHJaF
HIkTFdbEhnrBEVTFNJODDwiGOtz3hPJpYxENPoVnZok1z8wuNiNK5tQbdmQ9EQE11eE31i8+tpZJ
3OnrGkVfbAuy77VwDOJjBbFv9c216oXIFthnwjJ8+JTRfXYW8EtgJ2YxtSxHj78i4O9q8sufcLhA
fXSq1Ru5a9pWOYUVSTKCdYube+Du09Y4iAOkqNl2HpWcKHx3qLRmPxTl7CPuAAMkesz7u2dq4D4D
btAuRL8fVfSQ9qVHRfOb8ZATv/Jr60ZdUxMwVqGHYwSqFgROwKqv9TjpuhyH3/c+8nC0GiwoBHbG
YNYFB4Wjp5YqNqLfOF+Mzr4+IVMkg3gQLUJE92+v0014GTebA5+AzPi0k2xN9L8Gqx7aq3/OlTq3
ju4AuDMRbNQ5REnA4JENYxEe1nKsHFxQmhj55X+XM3eDx387vRKgh0wd54Y0CXi9CUBKu1SYChvN
S823eWkYvLIEiXfB0st5v8Iivf93lnOXjvLLBwGYA2cAp9F8dCglUHGOPjo2VdD52exlJc8RQmzJ
Dj+pJQnXoh/wyaixFoxWDMUw9KsiYFUXZoOUuhQd8+DWVfn+FV8QGxfddciaTQi+z7ZdxXGi8xTd
rqn0iygDIgel7YyFtlLuA8ckztTBU5/EP8BW+d5V+hpyHkvNf1RGcaKGKP64HeGHcFYLNuKVt9re
/7WexbmftGQIq6QsviRFfTeayoHgUbn/O0UKF5enXzniJ03fZZx3ZJMQ3vUjhjN31s56EradxfGL
YzzJLa/a7q/AyvXp3E0gMn++4Onv50i2Mml121YhqF5G1kMqEPBIsGisWEEqnDfyKToyOZCAG/l5
U53dPm37xQJbMq/qzLMb147oxTrHNvI3iZHZMUET2Ob0YUVK4czcY2bdAxZVpWysOXczLp3kk9V6
dYl45NXLF8U+Abde6nbcXSMJhSUwgEK6zm/4nUI40q00wi6tqkOcdNA9/+BaNIDueNskGt5Pi4AC
rqOfYqqIQhAQf+/VKeZMrqRX6yN4hJsuc0D75PUmfuBYKATMvNUoUfe4dGxPgh8btPWWGbX2cdGD
PO+DuLxODL7oUPAvDVEvLqX/1KygVjVNCpQ2Jrm7SCUg6F4D89BAFIYBgbpikaAQjPHKP42hXXUx
sZx4hE5lAaS2AHiX/uWIp+MplVDNMD3VfW9tfRh3VU4r6K4dbXyi5J922dGrs/Bh92piXHyts/eq
rsdRQ5hgB4m42f3t78qLxcQLVVAh2Tm9mvBYV/Wb9+RHtk7w3HrzuLw1cvczxCcdVNT35saIjnrv
wMIdvv/U3zcIZa9kO10hFAceWXOUGNCaKqJ4Qnqoh8jQFZT4GAvlKTFGs032NrqbrxpVKYMmw1fF
ANYH+l4/xQ4kM3S8FlSK6TLOnq4oJ9ktFbom8OZU1o6qThhod7pzGLj6ecJxR+Jk7vgbJMvcTDR7
03kBQMDYDNw4tJ//fCWO4khc+mrg5yFfAjv7gz3yjgB6ioDGuU6I1fARIcOES/wLLGPBeY8TCumF
9sAJiRzfp9pjsJifoYUhZKnU7CgUrnE0HMzS6FCk5G3mZMS/jmobnkEWAijHtisYEtjzBuRdb8Ft
6pITZeJaVDpoq336YrK/dXAiKHMQzXEGhyI0/AAkW6yqyJ1/CLEx+YD2rQO1PxlCjOqPmvGZVd6d
K96FycuKL0xdfTvnITqvs+Xszpk7sdpswFfOOugV4rXcKdASlwV6nZrKEJ4rnrTQ3KSTl+Nt9mDc
gpMNSIS/h77JnsNmdRUrcuYzYKvNQ5vJbDkINQ5T4+pUWpoMlYtha7mM7zNFX2E+32fvLtN3bPqU
mpla3KGANYb4wdQJolzfqUV5mndLn3S+TCvHDlEbN9NsIbjp1CB46p5yZMZ/TXFsO1wXK2to6Sn2
1vFgJL+h+zUW5rho/z6DKm3Nf+lWl3PhOTaHm7wRthQVmwkFrSacViexRila/0TvMdMJO51p6PP9
LWUM5E/wIiz7v8+3MC6ncl/uA1LM1Vb9H9RlEPBowNOpqkMBREoH3gkyo76DTD2p/nLISJ6dz1db
xgTMibK7UsN6VPz7cLnJ0nHqPntqLS2Ae7ZJxTo5ChlH8lS6i7YjOgaPVX7mQzI0u4WvGZQYESzj
Il6RHnBm0c4EVebjLYW++UEWbFArUo01A+aozLJ4cIApyH4l5skY6ZydZCRKyPTRGpfCaZkGc/Xt
jNy57JpMdAXK6C2h7ifNSBqXEub5HKHW98QQEczetaxIRDA0X/+sltnZuoTkURLkse2oYbbyCdIP
l4+FyKpPw/9hQr/43X1s/RgvzcyVOYyH/TGEhrvQZPDaBBeMyHbR5k3ZmlSTNaXc6tPaRP8H7f7d
ylgMyMiwscamqaQUN9xShPMatloylDyn2lMO5lEaymjC6JXO9T42oBD6bEMutzEisiIaUiPU3IPP
OMPyPbCiLjHwglSpwDRZapQFPpOxAtbwM3BDAsTdx+vKnhch0D/j0eTN3cUhrtZlZ23dk6qfHqOt
wQtlzi+dZw0HUDFmU3WD5+uSZ/ueM2ENooDjerUmfc9mEvMabUTa+wnj5NUf/NF9A/Av0qlNnRmR
qWsVTkui55rhPW8/zsdha69rqK+oAxRLvQOgYTIGPBjHS/1YiTCwgFn9m/9sNjGeqEuxvOGgMat6
aFkr8ZjhpjttRpJ7h4xJpIQsX5wHe/Dlt5BCCoXirBaquMDo4mP2ln6ZWVZ2ZRDKu/icM2v/Rrfg
rwxZpP0qQGNooNnPdtlxjrT191O8b4FQ+hujHwhia1YTWNgkQlUQWAzj1SlxIspCVmTm2a1uL2zc
D/FS4yqG4+2wprVtCrKsXyytI8AouJOHLFL0eblDfwgyZdiCTyE8+hPFC0bDnU5jMkj5f3Z3qXu8
ySRbKZq/yUIsWXbe9supePzGERQ0NzrC+jRE7OgjFVa/jyXxsQ5Mk1Q8hOnOHFC/VD1RgRyvkup2
cFQEtI67Mxil5qTOk2CWvTgp0kEpsnJMUFiArVw3aIrLlXI3efgyyvakx/4d5hb2ISHOdcXixDNQ
26F6BLsPkg9R0si0Nge5/49yX6hLF3vpz0Iov7/LdGfiYePTBikvlgGwYQUABtI8HDo4E1yUIjcd
gqNGKoFKHBNsd5chfm8QpTYZwb+ed2h6Rf7CsDRlX4KhUV/G1qtboXMOhLPs+JxvuoVdrMSKkDed
UL7OT8QamcbJ3/oqiRpKN+jkljYDFtFw2TWwzm5djUNcFq4OxfHuQnwZY86gsXpVkJdD9eJOWM9X
cEVfF8hCjpUA/bw4uD4c/SifHHw0WhoPBikJ0WwQtDVUugRBhLRTrdPGl1wdGE8DLuNvsgy/sfyj
47/QTzZiGZWroPMkKyyd9UlrB5hgnpCIMmOk7OTN9fn2oKbb+vXBADdhIdO8QejogdsbGnfcUDfM
oT9nofy0tZlzJI87GBDSkR7umeX9imykL+MqpTX4esFbNcfyF5JVGHq9hnwCbHZbnOLBhURs8umj
SKcCH88+a+CyxHBVieAXse35h5gl652UBXnNPkMKdl/UuNyG+w75y/BKQPIxO5G3UYgnDJKTNd3/
soO41lLGdf7wO18qNRzAcSWA7Hg7jGuXeovNPgDh7D7SZ4is0OCG7/VzG1DopF7bUhUzVqa2/JsN
YleCeQDKSo8fhM1XMkpZKQFEbJgY0UMUGplgDaBlwqIozQw5hzIFVajoDfkRgH2U/4xeXoFzGuZx
zhDcJDEaYeYZjbI9emyzv7z+NfRb4Xl+sCdPKNuQdnmvHtJKO0dQe3fG4D4ABNg0FHV4xrPHzq7c
3tR3VsJ45JwGIZXyJELiQb5CjIqknuN4Jl2cZZhHEhQsKz3uXCcQSYi/MXrtwXuxXCivEdv0oDaw
KK+EW++haHOEaC4nwIxAYFe0LL5paSdMHCrA0gn3kbF88hrkVnMosPOO+Cq2W7WyP1Y8L2ebmaXA
6LADbsOuqumxTeoFyCq9eLy/5VHEYPp7tdyLuBkX6gQAnCCdX5IYnrasLD+Ks4auB5XIN9SWIWJf
ln3Kc3dphQ+6UKw0wPNj93CkPbLimQ8iUHgmsb1YJZ9mbJ5/oxdhkkw8L8dvar/WhbRJzcTvBWeK
NogSUfFZ2N+PbzHyXxBTqMY3vqKiBETYH/Eqw1knMPj5EGczNqXaVGPOJxjdZTa3OdfzSVMEpD6u
BvJ0+MZFMHCQkXDqW45+MPlBCpetTc2/F3VxTXxnOp12YBmDEKheR9y85Y0A+MzK6wA5KpS0VRW2
LRljIPmq1rvGlPWZrpM1hDmUZ1TKWaXc7C5EZMywAiQq2xpbPaYZRwqiFSC31I3anMy6pWBfVT3+
4rdXLJ6TuD1MsRP5np1j0JdJFeDXi4P4fUVCQ1Af5q3cMRy5R7IvqU8JgBo+GcAm7sv2lXuUaFSi
WklApakYfLsJZDfX4L5Jz8FxQAmxTtKtHeUe262yVZtvc5SS/zacfNG3buJBItm3cOF7n8lvhoKz
IfYFcDS2IN/omLZ0fwMnyxk1xF5VM/Ck1x6kh8FMz0sDlOO+jt+R3rsNjeYCoIIdPLBPBtDDPM4w
r3TIFjawSGsGMHPaiKOZ0hyqJtsyLhTfNYZKlwKA/qbutrQFjkUtycpZBS2wZvLRcKywNtKxsnSb
4tBmJ1OWL+LSXUZnXZ5/YCX+v1PF2bdbSbHR7qwALdH1bGSjQM0iT9Yqvm2SEGJNYrpb2XY44hma
x2LXDKyje1oAH0fLuBI37YhhafvxVkHCYQvtz0V6O8pClgoJ/00r9VnYLagL/xwUNUrmj0AquAc8
2WRDuOvkZ7cGXwGkjV57rlXEshDQQF8TP8qkpEgVZWOZmotGlGfbJ/ybzDjo3JoBtTnNYW4xve91
Ga2a5EUHFcqbZKKEYEhcwkh9jJLjl+d5PerhFGcJfU6FzkWE3/3hJvl+BK39D+XFoxcmAOqlpaxo
qD95hpjvfjkKqDrwUIGBzwD4SWS6ZHFqYIwBlWO6iaeyJMo0pgD6/IxsS1Jva1As+58/t9VeSH6q
TuxJLDabo8F4x4mh6oUWh6tPLC9WpvOiVRDHRRtgMItacOD88GS2L6/77x5U2fLAs4v4eixA1zHf
eZzGr350REFMBBJKcgWzR3S5C3w2FamI1x56PBmKCZh/qX2PhK9/FlFIt3epRsBOV5q99SBRjnYS
SRexhmsRPKabVqJixgoy1fh8/N0R/pLu5YI+y9cE0bP5uHLdcHHLRXn8yamZX9Abo7GJRSkIcJU3
3SywnlNd9P5JDtaaO972ZR9BQ4QhBN0cHvqkDoMfANhzVR0zg4NgaS60VlA7tXOblX4nZjaIhmBT
nlGnoFcWZ9iXdH8=
`protect end_protected

