			
	parameter			DataWidth =				128,
						StashCapacity =			100, // isn't restricted to be > path length
						ORAMB =					512,
						ORAMU =					32,
						ORAML =					32,
						ORAMZ =					2
