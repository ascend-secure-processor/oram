

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RXzjYiAuFW9ZPRdJt+HwKKvDiZKOOS5JBj9nI3uhT2ZD3RBamqgYzr9woKSYklDDNGrYPt3Vz4kg
IoMuLciFKw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X89ALiF4NNmpknrwaY8kdJdFSvAFb7jqIAoHM+Hw3LRQolpRULqj/QwmbTaA312hoQfi2CQY5HqI
Ahl06JTL56m8wl/ntTv2NEoRSYaZy6LWSQoz6MN7FwxKH1CvgF4lxJ90pA5HaNCvc8/lQZM/5KJf
PNnx/1EHgCfhzPd7vVM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eLKPxpfhEiDRKuu9U/joqisAyt3gRNu2CwG3pWV7lJaLVj/R16rLY6DO9ikbZopbsmARNR4E0B5O
QYsWknng5H4M0diIXVCheMMQIhwVqmUzmr86AxMeMF+hph6jI35GuhbWxrNXnqczuzUXL4N21+Pk
O/g428xB/CE7P/d/g0lqX7Isq+gRt7SQ1K3BJwUyqRE2+PXrB9e8hFfc0Ud50fm7l7Xl8+j0kkHg
SBSgINukt6l0ZPOyQruUtifNOvjQFcQWJnuBN1HCPTMQ91WK4vX/WzYoo0TmKVPvjQo6yHKWUA62
2r+AAvv6nWa+8+hf8azqERjz9t8fkx+spZPrbg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z3w5n/ViwTWf7OT2We/wm1Pr408onv0vSDLVWNGbO8mmJA2K3qZNfGL+pNCU8VOWtN4FHYIKUko+
B1Lts+Wm+OEVYVIE8ZafgYqo7rjbySlMHHwYu0GHU+cG9grGKqv/OYI2FA6UG+yFmHNb9WvWwrSp
BJhJBcvgmTnRRg1BrbU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cx+av40gzEDGhpSKDGRQTx2hryoSHgEzGoDn5+saH1Ig8yg26yPtU2cfQx23ezlWFotTHjaDjnl0
8xFpsaz6yIKTJrsHRkDWNWrSFhNeTmGiLXHfGXJLAkNGSmmj+CfVj5pJGv1R7veVznLyONKgzc/3
NRy5LZxkkN0VfQGbzYFnyobdRDhQqlJL2tNJQk6lXUvW17VObvq04qY3wAku9tGocAsj6zWpKpB0
to4CqzHs973zJ+R39CwkFtyp7f0n1Cihhg9NaWOG/j0fXpmpIWB2UOAiZwUWHX6j8adc2APrnnhP
L2RShabm3V7IO0IZJ+Dek6dB5JL7agpUbMi5MA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15200)
`protect data_block
40SLVmb4ADMDZ7hZ1MKmNeeZg3/WTCnHX73F3YiVl0bZvjYDQdc9RnawKnMXyAz/PLcE3Vj8DG7u
GCAJKPCTw815VOgl7zZyXKw4d3Hl5HYOrC6JEgReSChp4dljrFpHQTpvaAs7+zkq3FXNdvenOMot
NylB4Q+HzSzVw11v4ol/Uwx9fw0B6GVO85I7RAX6rX3V0kcodY83HiivDao9EuNCo24fqzTVysEX
Sh3G7VvDAjBOCp3I5gswYeGmSNFlHmMxrCT0kmeiWYU8JQVglDS7/1uAdnl0pjSf+D5u7bqLsXYv
Ch7iaHQPi5WMMnfYqlJ2K0o80xzhTXd0blgekRf3iUnPLeRUtnsUNdEcc0d0LUIMw4rwEANXyTdg
Fyj7QVUluxndjgv416otIj4uRCdfD2p9ZZ/TZB+HDcI3hhOJMYP52sfeCI+Dz/wIIsOuMqXFUtLJ
D9GcZVovOr0tn5VXSPCqFcPP1ojzIxxm+S44mmHXyyXvn+RpEZADC9tZNmOCC8wx8qD2Y9hklZgt
pJootDpYZWxIo9zpfDTtDPBG1g+4hzLB8fy59wkRvV7w6abX3chz2NimrMnun2wcZyqit3bzrAwt
+eabo1R7PQGq8Z2iTSnAIs2tUoUaBz1dREk+xRJN/xwgeZ+i1MzI6HoaN+k9FyEwJkEgbxnBpaqT
uK9HkACgBbdTLdhg2px+65Q/xV+Pa8BX5v6sPbK5hjGi1+LRWSzmeK1o2H+rMIUlZhSYb1Zs2+xQ
CK/WNuSLwZ7aZ9x08s7GKSNOn00MPXHQ31wHcbm4XLg31XK4fCmTMaiVU7Wki8F0NAuBxmw8uNa7
gajiZEp51aOsFlEAGdYDO2D9A4c5MhvU3V4VtGAXv2McS4ey2Pjgt8ESYpXn7+xjUioBfdgQkBML
aLtHsMibHXLXOhAC97gNmWi6fO1ZvmJ4m3JZSWlSUNWsalR5J72eDaT8V4TxYbSWFEkWiZUsEtIS
0DQtCaiFvuJzgWrP/9NcDjtdFjafoTwzMLAfUTznVjoBLCaElxSbg61XWVH98jlN8aM+3HJ5RyNb
0Cd6nRIIm9esNhUSiWwSqQ03FOCiGtfjlPm1E9xKFIRDMbaqWzpRPL8SM6xcyZPkCS3JDT3P0mw4
3wZVUr6UNW4Y0BwLTOFZS6wk1OtTaOwRrMvZma4uT7s/bc1Ns55VTjWPmYXIpN0OifDDd9GCcTc5
x88aJ8sWiR8XmGpFm+ydkdnTAIkOjy3PeyYm6udf7IlAeDhDXwyyM0q0B/Jpmnr4oFM2smlCb0Kt
8GuJOgrqpl+ocMxJ0/wsZI53BfvQIfiTbUTFtotvCHTWODd1jKzlmkicmSsjZZS1tGtjR6/KKyMW
yPI0Fn48xJjr3ZMVfM1gCDQpO0ZewGeB6HihUW4tvTfxCwHLinOYpL40ysiP45nFvg2MNaa3colh
ATdVb/yH6QiYNAHE8OGWBRqFCuTB9F+w1BMCvQ85coXKrEMzLrvq44PlDOqlgTCbeZ075GiNfVP5
nsPJEVS33AaB4ZjniqD80iTvB7s4NcTLLskbCSFAeYkfx6vaEOG8snWniYjvkCQO7OjME3X8XFYY
Lt2DnahPVPOKl14+aH2Xprf9JqfemZbfrkstJWrPHhRd/wLf0GqkCAbCzBVOIV1Oa/kyHpKGits0
lZf1GfXdNT8WH3YO0oo5HgKn6ukFVP9ZdLyjO4GhmWYplHrE7JbJJ2lJcIiSoTXTQ53v1qn7wV3E
i2Zj8yt4vtCeV+6kFGw0rHAKYobuLU7umyH/ICoFgMqDoeU0QSO+60HLVCm405nI/+tpXSMSm7V+
VSnG0vYAP6XfrZkzpXUyDt8vRuXAMa8HbcpCDmBmg31AjZNeQjyflrDwqB3viZWB+PgHhOSsiB8B
4ofGmDHiHYAEGSe5ieqp/6NBF9Jtkl6R3iabhTcgdJFtJw44r6AztlRbb6PO5KvryS4bxvTsFu0C
HeUvbKpGbfbXZvgwyAZUz7gFKnzHIfHdah90Dxtqpj/up1JSxpFklkqHu4wusF+NiGslLglzdpX2
584r32mQNT5F1cjvn7FyYzQKnuliX5ziXWsqf6rNaG4ue59oZnqE0yGXIa5WZxmYxHrwLB6MSSaK
vAYyPBGEReh9ESZd2fVVOq/YfsFJ9V/JPpXrO9z1B9Ae35XSt7Bj8iP20I43otDHhjgY8lOowOeC
1M1Q+ZmvvbVjhS7so+M4tw58g+mxPNwHuOPMawr1RezVCQxfcpf2tnS4SoRwctOeYVQ6nmbadEGs
qoJ0OldXCOKmO0UJNnz11CC2UFPJ1o8RHiTXKIrJ8IjFZTgI6G8tr8hGSSOmil0XnDwgDTqnXtj5
1fWFxTbzcC6ZlKqO0nGrUqkyYvx4ZVKQ9nXf3q56u4VvgyuyHH6eVZ0BfZv2f/3Wyme7IBoRIlnK
y4vFdpY3JrpL+rfEGsezec469rwQ9vWQHQSN1GMhPky+xcDCOilyvefVbMa4tlqJAxY161xpG7Ts
+ZBy5z1stv0h10E3tBLoYYcagTHovkdEBYY7/Anh84fFtqpMclkMaWYyg+uZqGuVc80V12GW448N
dUfX35P96fh4spYqKwpAnSTyIxURrKm7E/xu6ULCt7y+e30LBBuzoePGsUEJmpNIkSMGtf109xnT
7fF/dVhJmpE2Q/vCjQ9WeOCqt4Po6OWN6aeT1LlIDdcBcvKJo1+82eBT7mNJw0zVe82R91yX/s7M
/yuhe6bd5ehV199/5+58bmEtxTYeCdJhbENhpUlczX1WKi3BANH/5qOfxJxnvMjcqX8ENbyKxDfz
eUw80Bwx7uVg7O3vo7+fRBlAXC7v3udBvMJK3PfLhXo6njNZ4X0VWMTwa7J0ztjSUKsezi464dwX
x4cvES2xKxjvgQQQCgA+1yovzGqwo299meTgwyuR8mlwgPnMLBYGTijqbjh5Ygv1hD9FLS6IY1VI
ikJw4v7Nym2nxDH8k0NUnvzsaY52oP6sj2up4qFyhfD+tM1DnYd+P2i+PJy6F1cIYUYAshlYHVJ9
UnCqJKO7/qkqAumAh2oFw0bvLgF3a8I6fbdjfpystxLyEvferNDzua8DX9cYeniZz/rAbdulNgkV
LfKKfVKwSabbHIVLBOMMoqydq/KG742jyNQdb0y5J1uDpG8rFjBkRAJRw/YZym6tWX9Nt3nfwPsq
u7n9X9UD1agm0+/v7bBPARMGa49Qoo/W7NoRxee2+VvRlovouzO3hqUMD2RHmiN/T+NRW27oGQPk
UOngBWkzL0pS0GK7bjyXufQtEngtfTC3RF+8xhVnUWZmgmVGS9kh6EFqajqam4z0AOHQgKmi3LTM
DOvXTSrEZIrSFRiw0c+ksvtE6F0xItf88iNwSfPaRQTiAja7H1vuE4g0j2sGdZVOFcdBvPuM7oJE
lA75/JVBpNpPDdrzUB+8xyIii9Yhrl0AWYBzrgt9e5kICSz6B02/GC6Gs+3V1AfMuLjrirbeMZqe
Z1zdoFtYlPZik+ZOcUXVKX40cZ7ta1dMoOIG7xAikRMNMgavmsE3NZXgRr5yXi56NF22gs9C+5bg
3YroByPUu4QgIefUJZJQmxuNCG05O+PLlH0GrmLtrMqU+NPIrRWmBmJNT05rVCF/F/Oz+ZZhZj5f
5/yt+HjKoHlLMsSnOpd3PP5Tkc2iU3KtIcVFtMt4AxNarEdOtDafQG/4k8Nho+k/cx+PmhjZOaZJ
/zoC1ZxjXYsn9uhOBOQfFh6dGRu9iK5gh4k/5J/O1sK9vW2CkwlDMScpIPEzOOI24b+3DT7qZG9a
HR7TAf3laP8aoqOHBcoTNor1KNe9zcRFaaikr6juk7xb+ASLTcf5zsaV734o2/yK8BMvZDL80Aw9
YAfsi1B6/TOWWVsisLi+Zh+GJnrLtFYcfMhGBFFQMo/JRK6QjpKUPTCAalBer2KeWLpo1hrJa+xL
rljBsopS5VTelBmZKYPM3vP71oFN0pHMNIBIOhuxcNnh3Gp7XXcvuYAHU/PZum1uhgvDRWCf0x7t
FQqyOlhLNo3x/zQkxPsPUAyoXMMlBY5k/mO2fm3aRZKLpp7FZTHPrNz6cwzHnQAHcjUnqbVK84nB
hTETuqN6Jg6ByFfjwGDtl/NYvzIpGd66YDoYSUwq2wuFb8rWZ2bAZ2wXJVavs03mfVarwJm0e4pl
EEVVAeew4Y+qAFhgEglEBRFXr9TIxAQ0O5GJKimTjo0L9cpqxw8zoChSXUum9TP006SF9n3quAiC
puPSeOnVJvBb+AxjwLNc2OnOcTtzucStaDn6074ZruayFwfiNpW9vYbssLAoJXg/plUvQ2y3Er6U
IfLGiQwLzAJX3Vv9L7L0cs++8IeCsq69obSewbiWXJvBwVUnSLXrYnkp+sVfDG8KHUTFJIGZvIBd
ZlYce5DtIflO9s0rwzbFxYRNhyM4brxOMWdtZ875+8Gjm77saKucRLYFdJ4gMhR+JLoEsULOy/El
M99NaUmJO/YFTFKV4DfOqQGIfuApHUhwGWIrXEGJcxzDqj6kQM2UBXBz0d5TcoymFaNaVJFHAyGv
6wo72q0/Kr2lRQycAJqmC4tMBTvG1GjdinSRGfMcYdUiP/YWolq6O4XiI/nzB7SJOm++80zEGL52
DaGKPwbaPpXyXiIsVuV7iKrB9dKGOB+OmeK1PJobmH0jYYNk+EKQML05CFWE1s3H5Nt3jT5/zJNa
qMq51/ox/VOzyAoZRlgd9/1s4zLeEobdFbrAVKv0Wt1d4ZW3jLBe7W3VEUI78Yx7PJOtI6PgYljY
gzoxghw+RDaTL3c2WpolxtvpKrdcZERk1TuH76G+J3LhQbDYauqRbtreQ1OgOG7qObQfFrCMtYPX
NJkqiVjE3SsBpc0NnIGutiBu89kdPDR/jsyVNpe/ffJEDyH4TOdK1JdSVw1PXo89pGvS2C+ENuug
c1vbFUSew3EleXnE9in93UHDzRu32M/dmmAN4Blsk01MbErmkZBK1XeW8BnXRw/L3Cquo+sgJbHh
2flBjmT/72mbJ+F3VJxGWCYMi6V6ee7JHz7IVJI0+p9oqmZCDKSl9S6wQ/L8pqOD0v4bTTYLvt6k
HR77y0yuqC2bwxKGj28aIdaxDnaRxHB6PsVo52A2WTP1WAlys2vRyg/nGZx989LaIBzFG6TKH6Zt
pcTm0LwYjPQ+ZMt1a9Nj3cw5XrUgTBJwCIzUIsDR1sxYxA4jPpysLLc+0k6bh+iPn+08t4dsI85N
a0S6ANzTC6CwMYb86IDYbUc2AbUbcbA93xETwdLtjnATC+wfOJv3AVl+Tln5f5p7cEWn3N3RqmdB
yJjcHdzlFv2Cp+cUrkF1z67Vxlohg6hMstckyGQ62iotIKO1q6NQpT/5SK8gV363OP3noQFc27w1
6zi+YE3ugxnnG/Bn4lHccOpJYAzOukmmMzfjjApS+epPSmZMWWYZeGHsp7bBD59T82Dv2D+RbRrn
3wsgokbZ8zAmcp196QF2ZhhvHOZ9H11hqDAUXy6ExLNw5YYalncaEv+/e0Y5WjwQ/oBbVmI7TxqM
o5oje5/67qrEOxktWNG5Al8gpEvIhXvrI2zVK9P4tNY8oQczsgP5uQeLu8H6eZrw+h9VLPl5qG7T
Ssrz+tKMSbs7Mxr524UoINVFK47eEq1CWkkY/CnH66z6higXRJETWI8ZU0az7vYNZBTg2qdjEaUU
5ypU3R5oVFQRYjHQBI7VIvWELVBEVGfX5hk5xxlwiQnZx+sRRWGMUSaZHQOxQXut0b2Ivmif+MVI
vc0IFHaem/L4TUj0hQx6OFUiP9tA4G/pCnNNHKbfT/n56+6J1dGxuUmmCif8sWyUQX+mPFtDXyJj
U9baydXU6E0c81nu2pyiGGOK3lHGQSDDptXZnIVCQbvFsFMjoQx9DC+UJpdlrNjCr2i66gIWXkBV
WvjbVH/pYerYi85O9EEg3Kknk5OvRfJPAjBcUSC10aB+Dy8zOlm/Kod+P1F7bKUzn4Dho2V/nw5C
d1F9BeGiGRdKeO1nzA2IygfAHoX5bdFLeyoE+tE7tKilakziZU5h5WvO5o5xY6uAcaTzsGIn+XXX
FVaBhY0yLzMozAi5xXEvHeyHVVP/ytwc/48MDrx29S/AvJvSMgjwLVut5OMOY6eIo8pgFS1fSi1q
fLPAa/HFaxoqMPHWoCyzA8O7MYaVts2+/dgR5xcezykEJxgvOAa9aHd4hRGrrU5bYwkECLfO7QyL
TAB1qTc+yj4gm4nt+/d3L9eNP3gDwfG6sMmhrhNWpdOk/Vym+avex0WrgdsWhR8kNZFKDawrMBEg
9KRzU9oFGw9MeH1DrCgO/+Y/UvaQQS4j8NBMwJuC7FzVZLxtj1jbYRKhsRbSY7iMfygCHfQZlRH6
Axa42XZzDcZL/7uIngglanGnU85DGDR6RAOLTNsMtLCmUXWGrq+ezpqBgdsINyTdsQVoY75oJTOu
kEEPz7LLdrkiASmuBmK8khYIoBn8Zecl33XjtaLI+uDOaAziAdjHb/+PvWvwI3UAkp2ec4qY7+SD
PIakU3jw3X99lLMYphkiKyAbAvFPywYoXtlVrGiBBPvTe8jaLtmeXQP4EkviazvvmLOW9dZ3sDnb
C6+U5CBEvDAEjJKHuWeNPhQvytA4PdYl7AmPcApDI158nQc4VytlscXP+SbvqSC0UvnSTjXOz74Q
lhSMuf56aHzgjEKwqzvRrxXuK62k50dfk2KKsSRwPvTXOwxCDTvuC1QtzCrlT5BAL9BYw6BSCOtq
Jir+q3PsdN9214gdjF34cycS6MSGLCO2fwvF9GMtmFQiFZpr5V2KwI6u6+rLIyF85jAlsfzy8RDz
zwRkC0WpE2BnWG22yXKBZQ5b98APKBuHbl8QUDDUC02Cm5c9HPjI+BnsJiMZ/gY7EDHvbA+HRa4l
lTxcuNtZSMlGncdPzMEx7e+bhxmq0ZMsHoz1Sx6BGT3pbUpIX4NfOutdi5iSO6FyKSpoR6+CXIa0
eU2UHMv6fpSu+2SaEIQQf6re9FK8U7ov0PPOu38l916W5dYR4xWXIoV/Y2XKkMFHf2qXdEFWRnp3
Y+6Q9EbRb56hGt+D7D3EocKoiTHj1hWCCrC4JwzHQ6nTdoYEYyb7FJsYCy7cF8a6Fzam91HPaypa
ln5fLtlwOfTYJ+UA9BwB1YwQQqEAwXanuWU5YMewR/7Bz4eqL+42xDQvdvuEcKCMIIPUdF6Nw2Kr
fwtuR2v729t73pDQScUCSlADnY8h56jAIOMqOWdIWqRZaK14DSmYOtEnDv1ZU0m4iElHs83jamNe
11gGkiXdz545Ik+LOOsbhG+PSTcMxqu5s9i00p/0Z8vJmpOQWMOw2TAa7oo8lEB7gXEMJ49QR222
LM9SU0YgZpcFxkqCo1TuDRURcQUcWgx59Ed3tIFL5Sid+CDVuhhdu/+wNXoghXcRFoom9HKUxCb7
wQIVgYRBdgAwwEuO4+h7GDaQeP5axurFmOxawQZtwL5r/Re+4YPgnrr3L+VRibnh3ZRDRivKy657
X+YJLXcGssqXQDQXHp5adOWMK8Po4MsXStXD45UWLmWgkj6N0iYDTPup4dywPY9JFKhEh9cxEgKT
uKbl0sP9+X84k/kZ+jhukYHP1muvUlPixewAyMp7vAMvtRNhxpYit4nESExF4gyY0SdYK7ygUnqu
l1Wgp2htdMjkx3z4tPCjcPOdqrFAl11gOrhTV5apA84z6jRRknXt2TUqBaSchowdbk55SL9WfC3t
m1teYEhwAqgvpl2G9prW7mEhQZuJPvpgmPFKlWuvc2hAShyO2l9XQejw/cXvEfks0JiK5bHkuTS3
Ybm739q24AlZuJr1LT/RH9AeCDlFELNImgZMzDNZw/blgX/T8vvhaI1uS+O2m69oM4j4RTB12dNk
hicrBSOQ55JdE7wUiHWb4SBmjMAfL8GqinTysoqJMbGcNZgb2eHXcf3MxqxeXHmcCLBs6h7vNW3X
Ujb53OBwxQHnFT14sdVRF/EK2V6N8oK89Lhy2qOCvq6z25zI87jRtIxw8oR9J6BhgvRJoGYOBCP2
8Qy76IR0Q0HvMiqL7qS8IxjUhHG8bhILb0O2dzx17w90cwLLrvirw655exI+kX1KJn4WMPd40rJ6
ZDVE5Lzv1PDIypUkf5y2EUYQEzFyWCzCATLhoB5pOvAQ43A9xeHMv0Doxix4hUpf+klluMZOqbDV
XzWj/NPWgBGLGklZOWmIUzFow4aPfg0V/MWVcFl7bpqnJPd1USyqDiI504FPwsoKHbRiMjkBnJN3
qus+5a+BrK5dUNu65gf0IeZFIrVQjXCVpGYEGI7FwfCwG1QArW+oQ+ST3ze4WFY9G2TJWS1xTHQa
NzwovB5zBFLB8bh+kD4R738AcarF0xLbWnJVd64d+yVlTw4SD9MZ7rBPq1/HXFvRX//QGMt+mQY6
1q74H+aj3EEHyMi98vZ//KScfV5hrbgMXGnSKxuRwgmkd+/nq3xN3vzZ574NtmC5rPoFoarhi9ia
WbKXGlSKpV927Ou4Gx6Tn7KrYhCeMLkw7mgifJP11DY064/11FWrY1bH0Yy7zSgPrzOOfh0hFN9R
Cv4ZgelIOUM6g1w5OKjpJNB3JgvvYSSsSssUmSQxqXUG+cwBHvwvA2RK3kdbO/p/U5kUCejhhcqn
XcIhPGg6iwmQTpoVSn7pb+s7BB/pqxBZw0uPpKLBIfA0y6JhQ2UB1AUselAInt2hpdlCFY4t8Q3q
aCV4KdFFGKlfEvznqhpr33wP4gHQlFHHxAvQQ+P9b2RkxT7uJOaopfg6ajLWD1Sxf9cwIiI7oj+N
kmmnUy6Nj6H/BG5pUmxi+NxbpuTO+6qO0bWI16wglT9BqCT+G42VtzNP0yfJeu/4MTzlqzf5yL8j
ezxhkvGrHseP/5Hd3FD53vnK4JyAJRguVArCmGrK2UXwO6ZRsmCD/CEOWA0hmb8kFYgX4vI/6N7g
ymSiECaGbTRYTBfXhVeq7JssbWWUNl4axA28XKtZO/e5n4pUJ6I8ap2xJqcaCTiqkXdundTOuwQn
17jBs96bpwU54lk9T14pjk3S4Ix5ZxfvrZTgi6RerGxuBmKFFQ64I2lDDdArhLso3oojcQcchyd+
/E2mDJ6Ux8mvsWmZ2zW5BCVRszr3ptP+Bv5Lkpt4kXrBv3rSmKck4s09f/JX27GT6pS/9VGtHlcI
jrF//vts5AWXVndIgcTmpL20rviISOow881L4qJVCQUcZu/uOEXvwyve+lrcs4aKLwkOLgEsnK59
dmoJvHaeXeQmVrbeGzMqNSWemzOTracVATwR0d7MDHrf5dqE/YVW33V6q3jen1QNijVQTvwEohTZ
pzOTWrnXqmqfdzlY4w+oMaP5izoUiv0uTOFk2r1ql3nbAGPLb7nBwbYVi7biMXxo74PfaXHEFgmS
S0hVolfOpHvwYP5YpnOi7YFSQzWCKq/FjfbxjpLG8x3Fdpb0rtdsNFxz2jRtc2OiYqLifSxVgwXu
Jtneh4PjoDA7ShKCdDNVqSJrvZuD6iJYTNnb+3cGTqthy8i29xPjKUh6rDQFJ3bB1J70jgyJEKLd
UXbmCZwh8cHXLTaJTg96GVuazc1HGU9JzYTNX29B4fSQGMIqp4J5UqSNF+FWzflTw9LkCg37qCuY
qv1n7YyyRdA1nzljla8G+Cf3HRvWOjq3HOCN3fK0JjuILeI0T1eOe/0Qk/eQO0XnMTLlALevtTmh
PtYWsnk3EaUFLZHXJnoaNasyqfXn3t41aFmJ7TGHG6XWhtpC9Or6FfCX9lirwc1h8ByxLfQPhALP
i3W8yeCsjIo+yR+QoNThI1yr4YE46RNT2KnEen3FsiOcRUD9w9keATJWMY/N9ismFC6rZQQ03k/V
Kg8UEaTpHTEvjjxXcMGve7oOsFLP83x9+XdNj9P+RdZdjV447TT3ipsTzfDF4kVtbeY+98FiKnzI
1SJWV4YXQ8rOYO88Xw90M//92ZlBADNuHquJj1sfrt/UDEn5LAdUD0eRjV3zYu7V70hTZVvqRRhJ
UuMMJdeYBkE0YOhc12rdrg4rcaOd6SYce1+mxpusIS04jS5dIrYvIvRndNDEE9ObfDm2rWGJcxPb
3Ob9CAHXDHKd2td7ZPpVqNb7CZv//xUtJ0eT7jOP+8tsd1C9KF3HRQHDazHpMpzuXhPNGyrWYx9j
jr+EM0UvdOoVaL365GiTgXEJB7NDtuRG5OSCE1tXq/ywwIVUAuMrLkWFt4mmevrhs/CaNZSpdJI+
ap2xvr+l78QrnYEZWPuAoLeZcX4hARbMnDFXmnSD37mVCzFpGCtwIqRNi+TOeV7tntkdMYvLVmhe
g/TZ52M81B2wdFSDydiunM7/9O5vJ8XkvVhsKTu9CU34cbWz8nKzEBGG3ww7xytMSteDo1xwv22B
SnSN5WwTr4V6tIJmAo1l1/8tjNzQE0vxcVojFFmLVclIsjQJENzl7Mcb/6/0f+KgRbHOnTs83JOc
xiPc5TnVSr0Lx6ZukscmFL9yU2LvmbG7tTJoro0tTyAh436qkwUiI9xCmiwsPoUXdaX36AOl9k2J
IGso8+5txNXDUnah4/O2KTgwpGxIQ/YB1LdlKcRhckTd7TiJD9Cq/CgEJy4gv5I4zalaj0eDA6cB
QgtobmtM5b6G1MXojqeMNaAImU5Hvi6YR6CowMlTCXA3LMVpIwCYz5JjyGB/E2+dCmjvRDuhngI5
QSJAapxkgd9L6oP1jYIOFeo+0Zzv3FsC6RWBDkVmgz6UthrEWdR4IlByzoFwfQov851CzqR+67k9
CntXn+YWIKu3Canl+kGEMFgIeDNqIcmCn9s9qMMqrHtrcJkSflr6/WSEi2pzHh3lxj8toECreyob
R40zZ3loKGl010/3g+U7l3Cg7ZLb/UzhUQ5GobuxZ3Tq+sA1Y7frRFRGsPCPBV9mxMMjAc9sX3wG
mH106FJhgRK3s/uPsZIJR7SGC90kzdbFQIlV1rEtuRqnPwd5Sm5QyjoDRY8M4Xf7kKKByfWs53UK
qX+wXn3bkKgrB+4WJWDPkILyRl2ZQawlGAp5Sw4DTr12vP/i+PizxcYk+TXX6s09/BSZmIaHqOc1
zjqQnNvhdNzm7Ey4qAlQ2peDtresEZuzpUiNunejepXAwQcG4S0Lsoq6NzxFPjSyemFIC9Dmz6Kw
on6rzSxxfv1J7n/XsQjxxSGPPKTuo351EuJyybdHW4Cr39OcZIn1xSDdobXFZ9AulejAjezwaolL
vENGNJ18a54dRS9VduxfWR36ymrdCPCEoL83qQiUyuNEu83I/gVV4sN+lQR4auolJ7DYkBMo5ARB
4I8fS3j4UqpAKAYPu926cCJu4IsL5rdKnSRCdQnS4xo+98yHxrPaSloAm2zjKTlptQQOBPdEuBMu
lSD23QPfLXnWgiplDlzqMwcAAYvdd7WoNsbKubsr4lCR4haNxbRMPTmd0gRKbj4VSAmflcOWxTlv
FrS4XEox3GD+5Mmt5P0IAmrd9mSzmNwUwHuVtzyknWb5k83AUPojp42iDwR/p3TSqOe7NsLmoXaM
nUOShAA6Z3o4RqajkGzO/5FRIuYxfpzZIOD8OTwxCs74k2xK9EVpBKcbq1M4xQOpQxfOr88PBCZS
qGppcI7ko6EkLKDlOkAoP4tTO+Gqf1ClhZZL6eipjswQZnuI0VU++qJyOwuW/WLhtUecF33QndTm
FUDPomemw352VCqNxEATDBetPTMB0K7h/e25+k0nVfs0PfghbtqsSJLmxOmJd6kv3ZFXUzimbBhH
uYvcCwlIOlx/Z5eSXmA9EMYN6OPK3WYf4JHqKDdyx8DPdcqwfOgsdN5DXzLTxKNIBat5uN8xs3tv
VC/U9tbWQTaAqUeFMo1FpAIW9616Zo+LLySE0SuuYk8nOI/Wktxj4PNHEiPHcwmXGe9J60+JwT66
0yvzjtkLOQ/k19dOfIkVvmmZZUV/JF7pTrOmm4Z5r6PcdzUb5xCht6uZYdmcC49GsEPATYC3S9e7
nOvuCk2SBrTaDFEzAUeCjWnpPuHrNvRGOwcsBRTxYuO5TakzZQ7JBTdsT4sxHXqmw0DzFtsKNXZ2
f253q42ir1Gg/Pnjspa8N6etP49CYhdFYZRZtTPPz/SYfS27S7aCHM3BIoA0kZ/4t8R1Gh8smxdx
YC6bXwqV2ShvRAWQ3k0IWC/ljP5abSZ1b9SzFxBin337dU+MWWtQj7ZOmthYXBnLRamelgJA9mRF
TLhGLPbh9ZpPFqPJYBsjhkQ67SDZoIpp7cHde0b4ofy3jcbNOmkPOQO9PEjhbY6knE8By0ixwZAr
FJ+iLEkQwZKQAhF9CBVUkR/okU7l6kAzU9/gNMSwzm71sebM4jhhduwOdivIZZ3hBVqW+QHVdwWc
Z897s4oWdqmzm+4vZljZgayJaBQqVe6uX3mGi7dW2rnrsQek63jjzz72Lbm8LY1MOtw4nfggQoiA
Q1zoV85Ox6a7w24YrPO0KLBP5uPRoJwkJr6bB08b2xNDunkb4XBV+p4NfPIT1SMGEq9MD7CrPDvf
vUd6P+QWFdXoxpyqJ5jqzci8Nt0O8sNfrz2+vFFVXTCnKbTknauM2VKcXIRsxuHw/cmtJKyt+PN0
jJaboWfUmnPEiMsnU5O13p7qyOr9jxtd2NPnd1kUv1qim/Mro6BC3O0NIFFT2CpYplio8Ul1ZGvH
g0iRMKMw0bFZRVgmfNy0usn7hoCF4Fmih4CCzZpzsXtDrkU8bf+u1nJ33Y5WH7h25b59hYagrLXk
X9Kw0Xq4xGq7hFU4YxrVvuz7a6mwRAWRJyHfj9NfZ0irRHkeLMKJfC8lWF3CMA9/tEpyfdgS8xwr
xyiaWv2Ot/p+SLhLrmj7Of+wTlDbzRGVaZcVLXvSlE2tMxKbf8WW2gJgfzsZAkrTZn9T46yYbKiP
ipLj187NE8XZXiIC3/2CZ3+gzsmB9GMnjAiyadFXRj6UTGJ0/kYfcaobZ6QrhI5S3qJfYh5UnTwg
LHXZ8GxO7POpFC3b+wEzn9/g8D3SZvZhW7T0aGnrq8OAFEB5bTwt4kVK6YNYhtf33vOz0DXQ8T1b
JSc+NUTs8c46SkO7CJxAe9qvvhzh7VmietZOw5Rzl3UEOIEjpcZYOhzgkyJJFuh2/EZcpIUJrx91
hl0BTF6WCJb/q6kc+kBhxpSk2dGCF1DblSHY5lotDvJCEUooMih3m16i6czGegro8291Sy4TlzO7
PS2oVfMSwep4W4S2c/OP2yQiHoHxbnmIRSq4btINP8ePt3tbH6+C+8UpR+I+wmh4wIGpOtRYyrMJ
FjLBSOYeZIpI0nIB2bg+4zas92n4BBU8ek7qtUPLaHimKvjXI0PHBwYjgfbnGZ3bGEsPoBi0YMPj
Y7BoacK07/bk7v2H032MgHV5RLnYcDBhXk0rSk/h/BuxhubYw9qQ0ba4FKxOhdZMFlUeNgE0+gSh
eN3mLF/3UO+v4T5EbVoEJ75p1GS5mTOFUH1gVxUR4N78nsVCkwLYVEQeYGi/ZpZ8z5mqyUiwRP/T
6XVk100zyPDAz2K3QQXpNgwZRxcohLbdO/QTajXY7Na4cR5u2cBHOtLvuxNHIUyWyY+zjUHakRZZ
iNLf7e9VBtjHd9oc0YAf4Wd6OkCtDpws6fye8PL5B/S5VcxgyLag/kGbv48CO4ovFF4L9L6s8N/M
9hxIteQqAjPRR0SH8mv4sA+OFrJWkWIcdsget/aGHbRILF+KSDgWdDGh94pxIUXO10cl8UFT8sCx
BE0OhPkKLxQso58Vzj8r1owAUgBH2lyE0/lfzrQrOo7hICWfvdWqiVKCPZ6Xz/KTOEivlM7GsN5D
alsEukzSPszvN0IEoiKYO80EI9OOMF3cxMDwrtEgh2+1cWGFszlMNgvhK4sqnl9/UFg6gB/Erbxs
IFsBPNtqd2KmkySHtfMpvbFCkIZoV2pbsJ5dqNGyf/9kb0gdfwaE/3+GRfcMQJA1HHz8eTG3Nr2f
qlulx+tVuXJaCM/Xmo2BNV8xFWhKCKxtM8dOBwvYb9DZoqUMh+nAjTD3778g0NybvwZEO2uKi13b
oa1xrXlEiIfILWlJhEOOH7bnG/6+k/cQBkVPoLrDOYhpYcDOhx3Az+Pk7a56Zjb/ZD5u/QBSM586
kRZRiIIil1+1whYf3QI+MvTmI8jHMUR/tNTqqp0CW6GR8/WaP23RjGSNscgzxX4vidjHzJH9ZHdS
ErY6xZGC2cj5d2Y4v4yEf2Flc7Sw5/IPOoC9gH6mOZIEQZT/vKWKRv07gQ7mjt6+INz1oNa1/KB9
iXin/my3mViNG4AKppQ1ASsFaL+kJ3dygIskhLhbodsaTfnuvUy+IVyuy3yYkeYguva5z/x//k69
ssApYcVssAc549/c9ebpPMnFYt5jk95J3DSxze6wcHp7BsajsIJgZsM63FWyIYS8sAUtLTIRJqBq
JUWNYJG8vdP9uBmFt+cFlz7WX9/qnvOawobaUsWl+Smxb+XU7k/M1dFpWDp4vxUQjmcjGVJFsz3g
PvTW5ZSnLO4yHIMC+FSog6DRMGSYaMz9XnSoJjVu90ghXgFx2IhaDkFl1nD1rsWAE7fRM/QB/8We
1uSRctytY2nKa4Qr8/j9QqPvT/7331cH2fduNxoX7f8J+LlGy4KBuI4Js3KyZ4YRqR3+GeukSsLn
G0kp8TIIUfcmtUOkhSNAIiUTGQl3f9FGj7imBnXr9FzeywHJohpXFsxQYQaq+mKtLRCUhMfwQrsk
zydrLqdfAPXl/zP8jhwyhzOw7btAFZm3Ab92COz0yQbM7Ky6/XkC3GEVEwS6pkGGeytBfLEYWtah
8PbOpgMROWFDmiDXfI5jWX1EzWhNchQO6zh38zNyP839yaLA+xZulM5/bFCzOEO3A+siOOtChaN6
CU5GTyXU8D07tYHroHjn5F/XP4iHhDI7zk/8Gf+NGG7UcnAbRAzwYozQYiqkShAFC39J/O6iQlna
YxxGfP9uLIf+Ch2zw+RdgQbEn7vZFbjng0f2eIwFoE2TN5aFGiBodKqQOpasQdZ3aURq2WLa/UPx
3VIjlYO821GLyuaBqSvkqzFPNVj6WWSfxXOBO6Z16MiNSiJw9V0bstulnzMsOzcau5GVrgdQHSeO
Hjp40hLc+eTokAwpRo4tjjbx0Ja5YRSCGHjur+2i6+L8u+OOY6+YRANc6ERN//Y75fg/cWFHeAv+
48TP2OuJVIxHLkV0Y0Qc0gUwP7OJ4fvHdf9fcEAYeijHm6Wst9WZzEee/uFkI1qZiaOc8tioWtk0
l7L08NXPyfv4Do8yTbkCHn6DhsXQTiha1JTHLIK8a7KQFrf06PxxuqpkDLCB4qPS3D+EXmnKlTOY
wr7//pL5aym3QgWR622L/Am8w9cdG0oVOc6/r5pecXFU1UqwGakjC1gsOEkxdr5pBpI/xaBtfmrm
l8ErxxQB4PWpWkoamyhz+xhlKv4feV6VfnDAViN+upLaHnO8IYj9ZQ9c9A/ZFTiQG9jNFzOTpKrs
UpN5576T4ryI5d2i+YZJ2VUdw/XnXwgEezD3PEsQcE1GpSNBO/Xai9T3vNObTrrwptMOCfO/Ebzg
TB8prYAZsuHBrhwCb/7Ccrbf1aB9U299jO5tEtgPObx7slBUEf/IKmbAiMG20ZRV5q+PojlzJQj4
Y8hlYDrcawXtS32C/jV7JmC6OX5X01dxeL9su2Rvmw1jvl1hNtnQwOKY39YO8JAiq89Bv2pEcZZ5
zAaqkaan9IbHyDE7HvB1Dy523dBLg9p/36pqb76ivK96v7KbHyNHMTdHA54WvbTS5qX0r++Eu7Ml
MW+GMw3Uf34s5jWs8nBbIGyUOHasm+a0oyk8tAEGgswpugEGpcptytjpZnzQKDDvOK7CYrhyjdZL
2tGB8xR45hWxSLEVljKhT0V6VtoGHlbcURMM+huzvBm7UKzJo4treJ6HRo4B1XtGAdKpr5zXw00A
vn6snLyR5/TZzwgRgSiytvV2e8+QTomq4k6lUggWIgcpFK7YHVKtvFzKO7JjzJ2w/xyOBZ5mMwuY
iAOpMcb7rOoITAGSkvC/apQYExBnx/OKAfMq3AXH4ItXWndBMUcGIgd/XDa0mLAVLCIduSxnbfEM
oWHXwhnEZUzdDOuN+zWz6mJlSu+ikFqPViPzbrKk2KVHqLXBXwhZUQn0TNpTKWBaMCMt1drvwQ+a
z9cuARlgBCS432wrNyON78liIqaiQmIkC5wI6BT4N7uLVwIXy0kNuj1NQdbvFOr17mXSBvbbUXbN
/Avg1DbmEtdlPROu1RC3d4u8AnTGPzvOU0GRr1jCaF0ZvOhpegsGuX2MBLL7gD3y/RTnoLeDYHno
dy+vk/5DHc6Gl67KQsusOsBsZ1YN3BybRhGIJKjFJzqY9tAmtKRo4xv4ELIYthjlH0PTeyjApezE
7AWMb6Ra+A3sQvxPq5Vjepj9qmBsjWZZ1fb9691tjNbSN9mUbnrPhssi7jFYivmD+mFPljju/Tqm
fU8u+JRZH12AP6A3KIfJeTeXW52KVURomuruD/CpP5T4ZgmYv4JajHvJSR4oF2NiyWprnNu8RHRV
ZkqsbzZDqYdnIc1PaGvRYhHsK7x3qJhcKlP9WlXhzOTLbbYvtO8oY3GHGNJebl1krCW4xntyCrI4
TX5ee9cz6wJcZ2gIL+v0wV5c3BIvVUl/a1hZbh9PRT4981IpFoAGc5Wpiy2+k6sPqEQQbeXYWqdc
BM0VDRoq07uIdlKqKyeWz78SX1CJKg69PxAxZYpjl1z0AyQm+mwtA8BMLCyW0gJ4k5G4zSZjj/al
rDnxp4wj6sG94iUqs394XbzgPUrvKSIIYmc1eTZqIjYpTp7feKhhjM1TKQAtpd/xvBbKGTv1iNeb
j20saagSzJq87NgWXVPedK4bltPPmXHFmUr0X2LU7DwYTVQjo4NG3ksVy0gnqzeiRo0dTVnWQPe2
0MDWXdcRVfVZq9KnCQZr9WfRyoOzhWZt8J7MsM+WPOHJtWKjrzbnLma8FKp3Ez7jbf+jpt9SRllU
9KSd+rEq9eb7zMKmbw0n8RIKeD6ctiy+JC+lhCDiWsZIPpvOpyiitMfLJ6fy2by31jHWD7O9qnLU
em2PUJ8Vimp6OqGVgCy6Y1cYSoIz8mfdaYFiYyTlPJ51Mn7dmp+VRH6TMKd/shPmmr/a6WXq+9Wg
DAuHWnZl5Rrehx5ZwgB4yFkvKiDAJ8+nQ0JSSHRQJOc4EzyHjjOk2puV2UABtKQvcVwJ4576wPhn
2xewlQTgMvczvXo/qs9AHev27pgHq8CkTmmApyAS+Y6ccWacESqiJWABfkg+HDlAeMf/OpVF47+d
uXrtrEx22FlVz2slui30bRW2UspZfvOqMwmoc6bLGEougvzqszLWSb6pW7dE/UzkK36tJ+JkPPEa
1rn51EAw6wLBoa+QyTWtgXt1c2x+2qmOEbNbzyvPALHWmz8zInKVcOzFQ36spDlkYqZ+LFUJ0zBc
h1lahuBsZyyjPciSDLkYpUH3Foo+E0AYnWzKYJSjO4sD2Be3X7m6T58nZvSMRGE0Aq3LWh/pdpfs
TrvJ0a5Vb0CKaYhpFyW+0rq4p4mL+2jUw6nAg+z9Caq9tWLnFlKa43OuMlk6x3nfHnAsqAa96S11
H2Mv9d3D287L2pyAVSwrhTLvP0WWIkDwAPmyzvSpDI1w765cMiw5z0MCACeaUGyCEPA0TB76qGsw
VIgic1n2ouGF3Evdp4PuEswgvl92hBNXRnoOJtPIyR/5Ca48vscH18rgpSJBdz8/VbYqGxQ0vwx7
r/bBcuz4pgtJ2pf6zFCYIiCaPKI4/3xTP3EtEWZgdrjfDY1YdMewQQZIN46v8KHNsXyy070cA0+u
vtu1ZgBYABdO6fmyx2h//pJxN12PVDEqDZqNTKiScevUnY1Iplz/xm+HMBOy4nxR1ZxWK6jlx2Li
FX+jhHmg6cTsEyMqXKjHjEOAoqv0D3LF5MW2FJq7pc9SWRnHdrlNlCjfQybFdrMJuGuO9FfjsJZo
6v66SxOk7PnebQcL4qu/XasFVpIkSiRuuHRz64PicE5Mr9Mg5Lnr9YEoE01kmtwJkvaYOcsf1TCv
1fHTmWG63bZYkF+Zi3JqswE/2QClVpTGD0IGsU3RZdkM36/QWWMLCJzSmNEvEy+8j/MUOlMZ4Mop
fnvX809TugqFzy3hw5VWPUB+dmq1fg7pb7C5yLUTLvVetGAhCCFZ9SJM05vmqZgaBB7fAPv7AysZ
92gVvCVz/Rd77RjpKCZD0GZpEGMgrz8L9VFyvTWj73oY3Q0y1FjP4auJ0LgvK+pRhlEtPI8JXxmt
+yDhAXVomXrSM9CtJ+gy4o2d3bXAZHGlOC/6YPiNt689XiMoRNTmOXKOkFPnaiQ+Uh5nqGIjl99r
d1APl0B3qeGde2qDA8sB/3mXeCzJVZP40QwCKeoJhpEBQRqBeM6iBdH3Sqdi2XKJxoBnBsKGwKC7
BHpexeLUiQkuvYTSVnOJIlJmknf+PCUCN7KfUlXDUqDbJAA/0UthcyqBDOMaseFXlq8zXUI0VVQu
bBIlo1H28J6nS4fuR9QA7IS3hPmQ2XdXeHVMgBa8+PZqsh4+/pl6Ji17BGsod7SSptSH99+0tfkH
9f/DvWsJ+LO0G7pzo4Zir7Mkh7Bg9OKhTR9uRt5hCVXbBLnV8dPq1tDgZGyEuv3hXyVoXmBi+61e
CBCmrEnsbn9BEvjBJcgJsWlsnRHeRW8ZPfAYVqjFu6VraUzR5v1fX3cHoO/Wo3mL3rxfXSuX+awO
8t9E6E8Er4rtPr3ONYn3vRQVvzfrpmZgytabZGftLqzY3ESO+xrKQ7HlrgXJQcqVviix2Gta+BNl
u0K7fPxv0pHF3F1Rv/y17myKZNs7Rgl2ReuswY8ZJLLgfO+oWwhemiBJ8LKpW+FZP2ojoppwsGdU
xghst4tKCm4gN7UiOVjar9Pq0jQqZ+TvJ8rPpt+PK3BjRwgRYCvnDHI1qlk2Z++eYTmtYIxXA1Gm
4zKhztvNT0xT+ZjexfyNbf1JrhLD8wE2qvJSOpop4+eVH7epUaxjnIb4n3eT1ystZAVB0EIAZnIy
RgYb9/Llk2b0sqKIzL7cgfrIY2RYML5ArDlP0dmB3IBjA7DYgrlACHAbj+CYeFJbduKp5f3WjaC6
6F4iUvsU/4GrxnxduTRmmva47nr/OCWHYvUFLCY1Nx1mYqD+FtroWci3I4cDuLO1gNus8zWD0UCx
BhHZogyTSbAwYs39R6G1Fcyz2YFvnxaUD36ao+F2V1gTX3f4CKCnGYyfkUxkeEKJreSjfZb+Obp+
U1F5fCyO3JKeGN5B96MwYoz3Ww2A/yTEElHeaJiQvXguGLei8yVvLtmM966FWhOUevLJQoPZX/ju
oulGJS3mOkwjt6urpzgupn4MtlcTWoVukig0BXvhJODpy702syYB/O4xhXJqye0uxm9Zn2KsNoeL
as6tUu8dUNlNOW2nCBicOrSsX4sK/BvjMKowYT5fS2LoU3/r2RDLsmeG3oZhp7u6xdhVcKr6SIJr
fVH7dEjnDADKJwHjfnhTkW58zaNTg5eukJvYtdnzjEazZX8CbvaI9M3PNDoBRGUexpOci9OPFj0b
FDjZEmIyK5Q8N9IgCgUb5AOlhxrTNr9Xb+qyMhfIoTqYpehd+g2Cl7ScTP1avplWOLg56yr8vMz0
nC9aj3wDbb7CbOP31EtyFNofYkOkuEh2aITR+lXVnoTyUWVQeIhDPW1Ri27BDvo9HDrCck72IxrK
eLx6OtqQOFx1OxEl8eNFAn+XErB+Ip2bSu1pkALLWgGAIZhv//JPkKqCF4gTdfEKnKf1cN3rHUqt
dlzm2C52512qOszitFvUM41UtCgSy8ZXgbWlZXk+76Ji8WOPxS1YvRFCxnz2zva8O81CMlaaup6A
GxwpB+C6bqxMJnxYhoav2G/PtppxG6pFGSzItAP3bbj2h5+MF9AikYcnLPhkA2li7EsTKRIg5k0u
vk4crlmGQ5rpmABktS8UfJvt7JlXUj0GkBOyjMFc3tmatQnCkSoO1AsXJv+aw/S1EAUgwNn/kVbb
1FC3LPjTbW7kdB14NmxYHitkR4MiB0d9diUIB9Mj9XqEx+rx6PQmlUttyIj7zga+k2VHUzyA2kQV
qMBPi2YOrpLjWTeG+X5OC+gnCgfm+AH9PhjiTPJ32GPlE7zBWvVRN1mCBqm1grziR0rthxStJsQH
3KMkz2UanuUNm+g9zZVPTOr5n2DKr0EwSHk7Fvi0YyVUqAUhHcI=
`protect end_protected

