

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KR2hDYVggE639152eMCgLSSMtTTekjXPZWOzQNYdeIgytaWoFmLQqGBShykbjg0InpCuHtXlC00H
UBfNgtEi7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YaSIXzB9EYuDVZzTYz22LglzuIzmUizH1/qutqnW3RInKTEZWeFioWlV5Bnz+AM89vvTsufs4hbR
g11zB641D0Qy0ayYwnxmWy+OATkeTu+hdImJ2up0Jbuc4y35ZVttIP0NrApkX7gQ9gk4t1YdO9lH
k3Vwu1OWZOst9sw0KjM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
2M9u9gJ08cKISkgO/6/5OBFK6/lOWflXkzM3CG5/xTD0L77pl2KQKT0sZuPlQNH0igw+BrFW4rSp
SZO3xZ6oka57ikqkoxUG3w/fZQxL6KpUPorVhKtYhFPF253FMXcnDgJXLEQoNNo2d378rxTANreh
iWydtIA7sQUDvbS0R7XuppqxO2WYhwo8pwGJzmzDSxp1j2cJ0HXEcPKgECpBBIxfhehRwwIf3XRp
RNdZ/xe2XRpBLxXbv8gtnQgsmeyEMhe2e6tFwVOQdHdJey6N5WfTjd/5lsCGuxpbALbQeZbUa0jM
yxt36eaTDaE+FYcxVRiSGBC0P81d5IoxtQLRGw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AqXevnlXYyOlpiJW+WiUuFfbiL7odODr71IO/WBRBfUdWAlHiLHWwJNGNXEL6HoCbKY+WjB4+yXK
kj3p2HBaARVxRZ5E+V10L0Ja3j69okSNEE3h8F5BgAFzb803E9D0LW852zxQEaq5XT8J9zsI6/W5
RNBhH+inUmnz39+NfBU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T6ATUzG0mHz5ITsZ+4ZTnfNDuhQOIgqIUwpEoajh/cBESiMACJ2YDvFSTIo0lhnXGbvzOxpwUf3W
oud5pPpBmMD2dFaaxMEm0EcFSeiVwyX7yNRlTWyn0sAE7uKYzMySv1t7Jbu+C97OQQfRaUhEFp3f
Yqyyp5zoeaTDqW62NGfPL5onjEN1C4rWV6nchMRGbSdu5eGGGYUQ7gGIQ5+XBzAPlL83EDWaS4IA
NFILH+mLrn7/QcvvDs2CpJZESojwLlHEeWmB/moAuQ6my37M9s3MKdiHhvZLeQnZlPnRF4SkQ0Is
jh16D2R7Hj7Wbio8lFRtNmmMi7Q/M4KkgLl3zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3744)
`protect data_block
U4hqJ7NwTHQLDFCm7pm1J1g5BUobgFPi0E0tpoMcWqFXeL/wgeaDDaaVonpTnBhQnE+7n2KANY5v
a8kcj1vwYiQm7m3oTuyTXjUbDwiR1KZd5mWr1AMNzJNmwzOGHgEc3tZEaMJMoUlha+QPiY3jEk3F
JEQBfB73bj1AX1Om3yqvgHlbyYPz0escerAvK/WsBfgagoicGuQR9+EGzP4/CPH28NN8iyoOOnFC
IeoL8vB1Ru8tTcY9/wt8hObSOXcMMtt2GimtdIg6gFCIj84Ey7DE79ZfQAmxEdTzO5otnqFZF9hr
+C2GAOm/tGslbVKRzwFR1lhFPdb9BVtEFSiw7KT1wix4Giqk5/Ayb0NMZBrBXsrL8WxTTV//IBof
Rie9MbvORgcNXIE26UUhWrQGastGov37O/pGzQWehmGGHj48zjE20a9AMRgHNaeqikAIr0OnYy4R
GYXrUGQMWc78bpqgX42S3/04QAbaVkXmMx4KSVgp2lDZYWhSiYF/KEw145fSeEoxpwEbf0aVmHf3
Ob0SB+6anDLUOAQN0Emw1rfN/r89UAur+Tntje1sYDcYz8Po3XPRHS4hoVfb0qxihKoGam5JiSpV
z3zwA7jPtuntJT/t0a1jmZUxcKTSMRLYhDqm5udbnhILHUoK+QKgOmyMC341/pDS84/8wWxxXAm6
CTp5opB6QIRusKRZEvS6IP+VkxMD2gX5DDJyBSZrcYZnxRZBnSvObrZDZ4axsvswjhOYQau6moFb
so8JZB7iwbLKGWkCMvkglPpyoByBKcAynI/oQ9RKQPnOVXNTRYYkrQ79yYsPdQtbHHnIb6MUA7sC
NjXFsUVrhESsYMkAhihwLAU613bhKTGzO7fxBcszk8hNITsP4BYvnZzxjyYYuI44bRJPEAMVxMHS
/9yyBVr9741q/TY9T3/q7nzY/DVwMm0wNoySKwVjjNUI7p3qDmA909U9OCbKxu81GBoYlHDe1305
gKqybsb++l/hwhbrfJJC9EyoGoeGifVVdyufMR3L8asY2uDbamAKbx1+WMKs9873wbnS2HeO47wt
m2YXONS61Rx/BolEbi5vnorRWaGcDCyJ3n8uxWedPVV2WpOOpjVz9Bs+kqDdRrsW1TycAeAjkRVE
HTZu07xm2bMOrT9m5rBZMIk46kerRGctFauKzy7kHeBXbEG7ySwfa7SNX/DfrP163LexPK0i4J/h
6f2mriqtAxC5kkqEvBvA9iVYTg84XqsdZOXFmLJUTDHgWLudgzC4pCuV0g++lYgQhHxJM1sZcDu2
YgVaOSqwCR3tDLsNDnmYMujDWPu9wyKYa4Da7jH2WMdrz+AEpj5FcTgQpgMNwO15XWm70ZzX1xIR
FSCT/LV8sdTAVrHtVB1fWwnHo9m55AGeSCKT+dz06JyF5UawPR8Y4BX2qwI8/J8aditJzG8JT4yE
akkPg7BjjjgRfnonoPacM401SVYLM39e5VE+bIgar/k7P4tHNrRBXTctwsqaEN/ZyNoxLLhUXtXJ
5YzpeCJUwKojz87ONkPctQGBubJd3ubGb8VU3AeE4Uy5ylPYW0GJegvzTG0Eo2+Gc2B0WBhYuGn8
kZevGY0MXnY9NXubLbcwRJNKJ/9v1zJHXojEnDUN6IbjiqcqH1YEcs83DRw5aP0S24DYqamxJhwV
GFkBnhw3blseN04E9puEN9yuvWRx0HGCGe2qMN7VhU7VxAxdgSsLZbMxXO3MhmuIwlj8euEemoE+
1100Tdrn06+D83duq9nSh8QNxByAoxRLWsw4CY4s+Zfgw0wr1Oxij8hBo72r4C9ul29gBthAMNRy
I+/HIiT8Loyu6BlfA0WDvPSPe1dTQrzF6vjAGyTcq+dBIAn1yKDo6H7wNqYmMHxgLunmpZspX32A
CoQ6LqeSrt6reaujyPIGe+6efEQZ2mUonhOT1POUQ0SSpFwp+b85dPCOWgwtSZfgBne0gDqEv5R+
68V6/bzZl0Ihjot7KULrMn8CN+r9pQQah6Z9M9vCeWN9Y3Ypvfw9fhpPfEP9d5cQ0XDmQWWqH3pp
TOKhori37iTH/k8MD+uL09aBbKhIWoJULAqUuayyyyWIS+d0mUySFXVmT+K724xKK/VrU8TlF3Ld
b3+qrQz1aZiHqgglOZvlQDy6Au6X681rKwyANbPD29PPs4I9uMFrtxZgp8iIVX5OwPSHPUZLnm73
t9mD69OLatiQYyUxFyhgjrEudtL5Kjk7DkFamuzFw6s90GqzI1wyNEUX//0geLMkmb1vilj4rOsU
suYd+jyQgHs/d3QfsXv1KquXVxOBpML9/JXxKX2v02QuXG3dt/gPL9WtNZxOed84pfIF9CLWTl4k
MoNGLgcx7W2XoE4j8EuO/bxIs7mpZ+Ka5h+hKBx7vEfBotH3dKk22iJeariaTZOpVB4oeu9vRcHX
zhpc/vWVCBBd0slkPz9zughJ/eTlVNe9CVWMG1JfIi035PU5+Zzhx1wLsxza1+we/Rtk/SkSUJGl
NB2rJ+0YpPAsNh7Sd9j3cryMXr1fdMbjmJCYngbpApYUXfpv2e+6ymuj3IV3yHVQ7t1dUDBtrcsJ
pI+qaul4vqcuig0obWWJ8SxnP1FAuZCSSNptIIGg1QMvAxhJjr+MOpjV5kD/FD53uWy8A1orCaPC
LoWw0J0UTtlu2dBkWZSBYYhkGZb2QdLBFrGbCJacIdctZCXUjOYlH55UJ5ISM7l4uLJqSQTCxF1t
5KeUf4hJaNj1E1jIJJgEIScBbq5ZoMOimN3DoaLuxL8O/gGPaMQGY/KZTqrEQkEuDYuBZlTJ1B1s
CBqBRIpsqSVybRuFn0f6Koi2th4XSbhgH2xiJBADCTGcrFD3jqcjeGJEwdKKilnE9G3B4YNr6am3
QsLtrG+RP9vFdc2iuknNwZh2kB8yvyglwKHt/gUOyZSgbB0/YDwjqqjMOzDTxe1aFGN8CzJz8c+c
pDV+Z+P8TJZnM6Qg1dYMuYpLf2FRL6EKLaYk98VxBkEjLdTwbqJNZ2UFs508cD9R7GYQn/YiR1QK
/qAfMYfRx4Jkpzv0ekthbDh7WjRWXinzgsdMzNj/rydXqfjXmI8MUpXoiLyO5N1ntstjWmmXugav
uTdawxNwMFl4e0LmKQk8AroICz/d/MIZ/Wqr9RRh9L1DmjDSTQ8Lw6CDZX/uUG0NS279U1va3BjD
6yzuJYUgi1ND9Qejo7OIpw2KEoGAgm5qemaZoCR4SGP2pMMeZYS4dovucSqUv1I8rMs/51tIixfI
2XOEF4WS0kc4WaqXpi0Kgv3LjXyTz8DScXSlHSpVKk0jEAmmlhcXolMh39muzp/dJR32n2M9zgun
q4f8b9rYyl8UG8M3a5Iq8l6FNz7QePYtiJ8YEPQLf1SxezqEXYqj2n5TSUgUBBSydPxY88o96g/S
SXDGHHZgm7EKtnEX/j/HuAhOC6jYvnKJoaCph/8NGqegsS2VLulae+c9OMVmDmUOji4igHPkoO2h
LM39A5FjHDqI9THUTmkGIj1nvnBwOa6eaDty4EImclydDrnI40nVrTs3tH0BTfv/xGE0IPyQ0KCE
jEVPX2A4OlxdK2aiQr2TN+dqevRPt3lMwD9Efebu/S7blHu9aEpeEu0amJPspIR+gCFKFcrgEBH3
87s9lO5CDcYsz7J/ck1noLnOvvoqlh1lh993X32koWkK7lZpA6UzfrQTeYDx9tU8wIXorvqfrOvR
0dkFcg+mQ/73EGZjZaIqM4+Z20GAwIMtJpeDOfRfUMOzLyhiPo2j10ochTm3qvM45RLkGJomtZwn
v7LozFHtOT972H5fU5pGLt5UxZ/vTSqUc8Uga2YbCtQKPTJqmkx/3xgdOvYqAcqPeTUtLmxGmD4p
Y0FEdT5KSBIN11lR/DTVTyrSHg+dm4+/1MRJaZusBz/pUVYwMtlNxZAuhGxmjOxa++F3UXzxn7/c
7LmFrqFV6XLcgmpXDg3oz5U6N3Ln57THXmauORF3Zr+xVbWroqvuEcSpbspkYaHcRqwSfYcebajW
kaOS6MzYWmAMGUsvAwaktm9YoSFjCg4RzbdMoJELXQECd5KYdTmGEwaj2k2+a1BV8O0WL+FFhov2
C+xr6G5z0Q8clZELWW91aYtUPe/v7dM/8Zj1DGmyqkVVjcAIQDY7brlmgKwn1TdK6bPtolaBk6tK
Ro7oGHWzITJju5wmHfP4WZyWDUmX5Dd61rLfmr8r3RxkoEvOpV5MsGHhuuj/YQ/HSNZPVtmRpxda
UJQ8QLJvg4/PdTNnxgIvUaOzCL1mvkraXnCDBS+sTF45jznVcFO3uhXaFcASy9ISh0AAJfa+fRet
DyijRkUyzjeB7gTgVrCXolf6l9vXtJe6eHnt/+nS/RAbH7miHihrFp0DcrbiJ69qhtLEIZTMDN5X
Cmcz0eNXMjRsBFHTzyKciZQHOBohmrUKjRhTjQAgIrrX//q4SanqrrY2sBjrLC3Di94TsWQNH7Bt
VtwS06ABm4Gw3uvdrRRxYwD29IBOzMql2Y3GYiFJMOmXlWi3tYOHOXvvcLVuQpT0HvhPGQITGK5Q
CfAjwPLKcRZ7bHn8Y1A9+mCu5uN+5rjK8GBsgpFoJzpPZxVY1I1Y8EJfFpk7U1J6ZCF2Yg7E9w6s
h8th4Mq6wTToEIpVEld8TPWgNsKxAgcPxhdaXWDc3C6XXdEtGxBhMsAr8TxIGL98dHFGCgLspznE
xK0w7qGRxQztB6M36B1XltG5BYvNMPlS2slZ1KBhbfq8hkMrzqoBlUH4sYXeDVO0pp5xKJJ/7rY8
AzjECl2dsBw27q+L7hiz6/9InnUyuwTI3ZcyX4d4aYzrk9UCR7k6rbB36sewXznB1UgYoLB05Oxd
SWgnmaItB4yikv+MV5UXEPrSeYUytB7D844udU/He1qIpl0b/IrSTsCOFoDO4g+DOR3pPfv7FyPC
LC0wwBC1V7Ysw+9+rpZAW1/JKY49Vbv8TDraSMTpEjC44TC7kCPe
`protect end_protected

