
	// TODO get rid of this --- merge as ORAMC into PathORAM.vh --- why?  C is a top level parameter!
			
	parameter					StashCapacity =		100 // isn't restricted to be > path length
