

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l8Mm3uT6bf5K1wGbID3Q5kSYd5+xy2fhZX/Nv8oZT8y1S/Ad22SsU4vZRhFuJqL/nyC4p3y3Lth4
6M5+6CdVKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HQSiZb/tOXsBCIGXz7zZ3qbVqe1wQnY7qnjESBe5HHywzg+HtAs6Tmb3hqv75H5py0vdvAVHDEZF
pHukrgjn7a+NUmMmICaESWZFlhX4r3lFd2CvK6UYPnW4PY89l7zt+4UEi7iQYYXgnc+dmJQkxKyR
czFH3ewJVCRq73U3rgw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wX0o3JwnbuVMV98ncE1DqqoDPH1GALbHifxbAtDIgSlbh7LVfKEVlDmNEwaoRiPg6Nzyu6IaPV1o
tRn11RTA5coNDHw2t3WA35Vo48MPMVGSic+VmYhDy/ZyYvlcpBBiP6Xv45DRBuP8Pq0qarKrHWmh
gtDWMv1TIlCZZkPtky0iEexTjqyl+o4QN81FaTkY0xUvqtatWToZb/sFBxggHCdrOKDtvmHdgf6w
nPaREcYqdEf3M6gbK3AMYRNW6UxDiBEmDPKzzl1CfdjQ9dHw1yN9cxFdNDa9hN4e8h1J6rEFukI+
kktc2YpkvM4GQmA6hbbwHkTInaxwrxiaAeMXVg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W4VsVa8BcTl9eT8qdzHRDe+ckZ4I82pki+wvcNodjzkYHKkeAOstIXW+MaylRrPPSOhRW/VyObP0
lDqvu6u2d04AbflXMDF3NkxcaVwtkPbaVY2l2+HAZB65Y8JPgUSiSv5ETyA0SkOdG1xglgR/dlrq
zUudXoFN9NDVP867A8k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HyVkAaBVS0MGm+kFNljOiigb1aU/hKRqYUxH1TYnpaE62cSIAQdoTEBbpGN4Wtkf5AdTqZ83so8e
AspZF/2Iw9WQ+jss/fF/FpSjVnlNko7e5IrSxrDLj64zJLsoiwVpoHdMYOhhpVokbjQxaX2cL+9i
WX47RiqhKQRRpS2Riw0u3fc46KDAcANfhYNXWNBan9dFDZpk+HFWfrWsjBxO7aXfxmFROZdwfm2c
btLOsZeCPHCcMB3TXfvD0iSmjTPMVdwsWUUYafKY+8yskxKA0ZhohRB91+1ir8Y8/EF10S3nK9yx
Eud3AVoWKk4TMyARjT+Hk8V8zmWsBIWLbZTThw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 157312)
`protect data_block
ygAv/wnLcEuDZQLBSMp1RO3UV7SKCZYQal19GJ94I6jy84Q+8s5ecvUT19eVz1s4qJi6tRq+S5df
Ka5kZ0NzE4qWOfunedqEB+18szU7Wq7vab6qqcE4qPUhVtY/gE2lK1YhqtmV91uNYFtUC+LehjCt
DxANTHwq/AG6+myd2ism6lLNFrxZBTHzNDktvQ1el3gEPArjPrZn6c6QvgPvAJWQ0YxXe+L0Egq4
f0o03B/UJ2faKA8tMAiN1vRrPMquaBSTW9SRtkPY8345gmecSCpvyMXJbAS7smRAtdy7aeuhaeMm
ALrp8qb/wREIwve2Pkv6S72vLdvRFsSAeWZMCK5v0mHaUKy1Zgc3usgViH8tIqhK6c2U8r5WKThM
G1qzUEfClYeNSnjOGzVvKeXHM6tZn42jfQxdE/Jpj0ZmoiDvFQWR7yOtTxKB7DzjzS2SeCNwTzdv
6qHQJIb+Cjhlb0VR4ToJV4fv9HMuXYcmQ+iXf14GWmkE2toKcJhU7ShXxdrQcluoN2dBtUIGdfsm
3i2zEc/2QwPSk+ETwT341RqaEDE09ibO8V9hs5qEutL4tMddMIkeGUxiZmSRoGJFFIpfgCqbnEYD
+lgSPi1FzQ9nKOMXgiqSGgEIISjkjDUSnQuGoAZTdTPkmaSgDCbbGC5zE/TW9xuKdrmoAQK1Nj3M
QW7ThPesOh65DtydMZBInoEaE+SbG7bf5yaZkZ/acIR3xtsTFSX9kTZlMCcGJAcZT0DXrDnMLrGC
mJ38avPs9TpDgS4Nra01n08nnP/NOWY2Bj3Ypn8ImGEpzIlibHVfGnnFxVIzKlJlNDmP+0il1esY
kpOeoIHCi037KqtUqUdB84QEW/suhpKMgPRpZVfPJDS2FT9y26e/HvVmYH2k6yewEoBgZG96Acjg
bTYJTLxS4b2Cz9B6i4nxh9V583Pp869a2pUnG5cpnnFmzeHFgWFYe++qZUavzJshtpzr3KPyVZBy
Lh/VrCJHkF3dlc9COaANxoCQ2W4mJ/6HrLSxCSgsOmHLRBm068lFDXAHA4tx186gmTPbMlrkWSVu
obsVDUpcT5APL0erHYByqZbhLX7YKlQbFAsyrIEpQvc/N1P4GjqEbRKjL0f7aiC1aJWN9TaobHzG
0YnNcv+m+UDBq3xX7YgTctjFyehDlVS62i+qpiYMelk9DasmeXAsTKXiTXaz/F7gyj2XC4+V6bop
VUrmFZQUZdKvbFAsjA/FLnE2Uf+Jd+NrWT3d0B/dOcwd2+m/62dLW1C3ldu+wAPTyw0Z4kDyKtmn
RhgMvXIgSFRfK+8aEOesMK83SP6yZvtdP06guyr+bCFPDu/KvgSZBgIKABr5p5CHzosMtielI2Sc
wk5KK5a7EJBSE7u6Vy+JPqzQ/o/78ol7T3W/ed9daCFAgqZ4GLUN3UPPdcWQBo1YFO/OJClRYcvx
9ntI1ti+TLfLEugvynAA7xPaBUWXJKOgLc4PQz+lmpPV/S+eblZvB3kyKtFgi7KqxceRsCeu91vz
0kymPbI16Ypa5mWEe1Sre5ZM4DVpGluE/EQnC2p3JVQk0GEpUxlVbVoarGvN3izm8xiTshGrWDql
9YTOFm9lLxsPK1RySFP7isqkiAqkZAqIxamd0KUL+TE6i7xCJL5SZTwNl/01QflXKG2MAs30QOkM
yWYFsAke/yNhJ4i2/R1M93In8wS5y0EQsSDLhLGwcWd+czJQjYZbMF5QFuUMd4VVCVxWrUbAvCt0
BBZSaYy8vVZOUCB1dNUQYW0A3hoHFUtNjQqK+25GXT3pQ+eIUpKCZc1ggylbazoPXOH0ib0BhXCu
rb16ijstT5gRAgU0Mn/N2aoeNrR/FbO6/jUzJZ6/sgC1O8cLgh+r8CVVTJWMPB9d1VHoHm1pBFQs
9/E8R6I669XydsvHFXWe0VWYfeowyVRRUN97gyN2DumyYaGPDV/1IkvbhQdaUsttqbyqUIUG06mF
lx2R+d8yEHyrE6NLC36pS/62od4MU7TaF+8B6yLq/mlwOxtaSFdlYDwcFXAYl/2DE8TzJEC4UKQC
yKYk8J4sVOZGp2ThihTyO9UPL+7Bqw5hMHiYAINNux2TaB1yHq3sTUN3To2rJAvZwdtVsvK8JZNj
+8XGry5o5K/VzHeCwkLaCQHexMvigqpp9GkEC6jxkQjnvWlsEDBSod1OcWacWOmSe67B3qUnn5+6
WJ5VAHw0whfsFocffHU8HpbbfNJQo0DIy1G4jMjEz467AZkH2KeWV+SM47wYOW6QowYQ8k0wgrd7
8jbYxW1bKTMDdCL4pddEABhsR41JEHm5ZqO1HqY4BWMu17xKQcMQGkg9+VVEveeNCY8Y4vYJekzn
+zSqxx86T+Qo3Y0b1jQrMC3+I8obSDPx5DqwlHdxHlECZHUxtcpZ267PrYSg5HA2qEz3jvrXrGYk
MRiOags6v7apkN73FSKJTLkvzWCb2LoxgvLFIvPCjDYROyCthECmLy9bKuuz7BaxbHsNU45ZpIKN
U80KMfpBrycVBz8ILSnzOzi4uBFW6Zo7cfLNRpx5XG94d8h8GXLjKX/oVOwe498yN7/Lgu9+W/pV
+c6dFgYKsNygZV23h2AuUJl0isH16azvBPzWTxIURIezE0eeD4irPIr7BgQsYJruUrJKyz1P3wr9
5zPqTOj+SeJJqPDBJArCXd+xrrowYvjIfsHlqzdXq0BzEBNjYwqLMWvR4UzDe1KBoQ9ZPIBVlQ7E
OVoZSsGw+lDWYHqXpLuvJEG8ROocYTsxw+WZWbul/pCaTEI1pK91Tn/UOa1mZ7gqIfECy6DOg3wp
3VTHwuLvBtnmi9panYYqet2HdTfmtZT5dPFa/JbAdKYRrph9hlcLS/+aetHDFQtmxe55/CzhCMrI
SWNeFqkYyMvY1gFZf++G73IxUwzCeCdI4g/1ypES0wpjYTHuUUFQyLi5O/uoOYxLSDR/bIKVYQa/
6j9Jo9pDlxo0QLF6LCn5t1KOx8F+1PhVugrB3KYQpLjRahaMtp63rn3Qpnsjnm7oylPDPMEtbtoV
wj1H+yTY8lvpro8boohhwgUlEJJF0sKboXJ8IkX44wElwJ9U+V38tFzwNklqAPUptiIheGMzME7a
PnGfM3MzF4NdNmZ3F5d0JCnxJlv6Lsb/z5tpk9cIyhIrp4mKppje/R1yflEkAdFEAPjiiIInDKb1
8IpNa3U2zEjEhYLgi7p5DKz1anZzVM1D3FMqgSH669g5xDAlxPCHjspSlaWApI9fsvSMGsKOAtfC
0fmKsjIZtrJzP1N9F6ud0M9EocigwmCUOGlVKkQFLTsZwtujXptuShYlL6rn4JM67sQkIITbtdFl
LCC978VRd9xYsiVV5PxZC6gGqxnwUsX4rqrtxxjciIQV7YaiKmATqVXdVi+eSxXKeUnHsgdt8Cyp
cZkqfjt+/54pyDq/ebCPpzFZIuKclmSRma6BMaTMDozo25dFvkc9h/N2Y5X4p/JEUc4WH2oo5EW4
d/51bADucWoJqA4pwI+T0x5f3OGOoWi5APn0rbConBD2zul/OWWDIFa3CrCxGVkfaBNin18eTz53
ecCSLJu4UttQsRjEgDrXh3lXjZrp/YRxIKuHP70YgdhFNo73vPASGzcc1XQmEpMgX+HriUzD+Biq
c4Fl3Ja/beqM6g0oBbsXlPeMjrBG6lrxTITJKbqfQOeTjzuimclHT68sUc7YzehdWAmYw/PxMjHz
rt+Qpeisw0A1SEaENpUrJ9fwx1SbyaMHL0Ibj2t9FilTjGYUNHDNFfcqsRfvJKp9pD5kPqrvibMd
pMTK8pv5L0J70mXyFlfL9P8QadKMMx1NG3mrtCZlZVpkbr/8XJFEF3o+CslhfEaCQGzEvl/dQvA0
E9Se1b1Buia78ghtwZHes5iRhImFl6l/5+DvpM6Pmz94PJOT2s2S9+I1mLPnHfkpSDkjUQuXJl2d
9XPYcqFny3JwXWBkOTMxo2nHHs3f8pz5/r2bbFP3D5fUg3R9EBJZeXnSDqHKYXNYA1fsaNMI5bfs
X6LjjjZulU9pAiLczobPR9LGp7G6ykDUaN0YpTcQsslJLVJ817pecR2VnD6L44XxSHsOJcHE1r92
3sWdDxqi8wwOqi6IHuqUFi2nl5m6tVnlOiXfZz4JMTO5Wnr+pJr745kEsaRahmXtQRqrro6XYVIB
GYIMBZJ8X9SRzXmV1SHePN2+Id1Q01wJLM1SztSTmdncOZNsPWqHVNO3tUwl/3IJmaDao8U009Zh
/tVxqmAO3qxmDTcc6UE5DXR94J/GgbbrdbP4+Hu6Sa7SKxYidTrNT3dLEe8V+wKRKzYmV4OvFGu6
BfaH4Pl6jejveEpL/jvcnojg9nKSPGSuSECvS6XXGA3fJwTma4jxBROrSU6tWtWsg4GfUHQqO+yz
Xra3sXzbXZUqxwS4cOvJc+HOxfG/N0oRc9hhxiYCqkGgapPgpPALksqHPAeYDyjC3e4QcDcGHOhK
nUvQThn1z35v/Y1Y90pXKhSN++bRRPWhjyLXjxA8HYzS04YX/iC9pzG2cvDdib9ZJ9vE1qpO1QAg
L7KXlQEEQi51rsvM4aOmtPcCmAgNMCuyChk4M12DRKx7Z/WfSqqU9mOS88+qTFOTRUN+w3NTQ/47
77Hvo2pb2bd1nsyBxF4+KDnXkjqZz+WjGpWA2/MQPbE1f7/CE8lGj+IFTswF4zq3hSjxJ7kJXwFu
GHsQgnX2n/KWPLVUkg1luaPzx/Q4p1aMp4E94gGLIkpshgwF3l4Q1kCHsZ1hSMJZmXIN5x+4txPH
wQCMLJjnF4oxYUxdxG0R1FD0rNZ7572YrwXBGGaN9rBpEfpg/QnyKcOvjMj7+MEcW0klDguIw25b
1Mmv/VSGfWsouOVdZltWovsjFirtbasweXKzA0u/GtoQfNGGX4TfqaMPDkSNzkG7KEVRg5go3HYt
MB7HI6x7JqXtZvEaRIES1Aes3HFjSDrcbHp9XW2wegeIFg1N7wmpZMF116123s2JRw+Xs7vGqEem
6HSGSo+HtSSdBAsX+c3kmv8en7TPpdHe85gUurLwwTL/1ar3zLNB8TAnZBCiaKsu69KBmtI01cyn
tXxzKlB0LvrtJwbGnP4BOK05mVjMeLlpIAMMphwA99xnN1q5h5BBaf51prnavmR/QvexVc5gyLRp
FUKqf/KmqrvIZxhMLA/h1bk7hpgTliSrUvrmEkq/QI6e9rVK4SGTCldhi8rMLYUaxXHKTguR3ukF
eUF2ARfHxLMj28xz6wf/xRZCreZrNuSCAjszDS5t7GKh0imjdhVAfvSycV8V/5OADl3x96BnKbWz
Gu1GQGZ6uNMeQ2Ol7CCJYnKKRsMOXysPpfUQYGeE/8glJqf6bSoT1pjz01gASX82tQOLQqULD/U0
acqDaBg2GaJUMIApv03oSzWIsa6ZJcRNdKulg6/Ce4oIQRfSgNuf+x6hQaGJFlZspx1++i2l0kjk
ksUrxljBWfsdwWTxgdm6VVeMTclc+Ou4diAxn6weH9ehvZOTGSlaLrtt2Ccf05gvSJSGk4WN/kIV
Z5Q3stskjGxDaqMmJDltGlM910DguN9jX5gOTEYS4ol0IIwiW9jm6Bmq+wyY+hxi50o4JNrLDybY
01hN3H18w7WO6TKXuoOZIv1LMYtUgWU8M6F3YLo98L+VsqVC0+/5j69dlarAxga5+go9pLXCXvIZ
28ydZeEd1px65W0I9CotN8qzaejJWeSnS0eVDeEdkv7+eGxvDfp35v2jOzeTcoRqLQ3AF66McItn
kmajUrDvIPV1jJBr/Vv+URRgm2+muOB4G9DAor11KEXNBcX+i1dnhNiGuplIUYsiuHe2zxixa9Ql
nd+XW0gAHoYygtHkJrCJ2qjcNExBLz6X8kBMWYqLm8nv9LVE+apBaVWFRYUHBDoPGpcLejm/HEu3
LeLw9QTIeZ1wHF4VT2hkhfeKJ+vhAXoZdk8JBnvO/PS1iuemzxfKKxPJmHvS9hIpopawRkCg9mj8
VFieycQYGwWx6ftMiEAtfzMHvPoIa15TSFXuH8Sd3u3mmT836QMI88lOzrFWGpZD2sbst3Avxj4U
NyyM9jADNbbHwjGCcJdhDm0Rwj38twFZtwL+MP0yKZJBMemE4wS/8ti6NcJfak2GmvkBe12T5rph
vRZhw2aWdt/LQPEtOqeg+ymOrb+1ES1hOAcMN4Dq4h8PbLCtRJtRYzwe0q4zf/dOrZxvCEsZMJUa
NW2YQ2Zh569sVPaUoAfhmoqVBRe36iZeOlftFvnyNcLBpgzB1W1mEVgEzC94UYEFWLyzmUuycZ31
4aCqRVM4/lYYnTJGGQthFhJESitM+fZzFqYo9T/hoeIgCH4qYQCsNzQzAJ9ltEK5yat5QxbQPc6T
nyWei3j07XVjH35EyphMxTjp4Mweu4mfEvZXO20U/rq3+6res+y4L0DMOju+NqRIVYTIfQ3cAaMF
lxQk0PI1f48w0cHzVtJ8+pLcMddA6g9wnEKQFKuilCckfV0LuQ2w8J31GZMoNRHqw6omleQsPZCe
Rogcaj7H/2PD/JfHvzMQusIsjCAcWhMY6p9upPCJvyALBHyNH835Fdd+dooiWhWXVSz8BvJ1CwWe
T92etdrbJgqlyZJkjc7aZmqQkj9LsHT9J8rGlezEn1zEz/fFQ0GPpJBPiz4DoLXgouvYnHm8gvV1
7Jhh5nzmYaPREj/nc3f61N05QJw81gYuMcuKd19PZlRA86r9D04iaPUQmXkrqoVGE7zec0aWaJsc
CukQkLW/GuNvAbdEMdwUKlG54FXXuFiV5kpIEMi9XFpwN9QiULMbQwyf5IxrTPAAXXyOYW/zHHij
kAS5rjcS44itlN07QkfJ/EyBAXIXwTWVhsGMQN0S3glR8B/B2SxROdoCvfk8wl0ldMkrbGzHCdel
3SR26pQqWcdFOmLGm+EfUY4MfdYYJ86B3gEqgOzi/TB0DgDFZh59ee4Rr/Kk17Kon9CP5t4NbCP5
le33TTK0rnakJ8KaPDDix2fXcOYORX+xeH+cT+91qCM7Sfnkyhi77vHJi7y2/kQ6JaDKI3P33zfl
fMifYqIQ7yUsIveQK4MO+t9ggPgi+lp30zxSfsONBlwEFMKp+0X9PtYtdJkE/ufkpUBW9I/iIg5i
e6V/mVebEFD+Tmd9+1hueCXtMsbswXIEFIjG4fdDgzBCELqtufvEmX+25jWxTNzqev+lSqC8jyJY
lTaOkaPqUd0ZvSEZnFdNOx3VWxF7li8gnLOkmduzsbo5p4RgucIGrunB2MrcWz59F0XZPv6g7GYU
OxyWL+fmmsVn9P4acWtR+9PMwaXX+I+69B/PJgq9z8NWc/FhSX/mgPkuw6g+o7vFCf7o00nEkGvW
GpkYMxRWW+6+M+MkWHmZxfN0XgJeQDH0o16ZugE3OtvEE5vrjJy+mLuxLkPwZ83ejwa25KrqieK6
G+s7ZvgkAkp2ZO+PXD3tOcPpMVkhdV81TaA/OjLoNnluLWNKJke91i0jMSuJzRW3HLdvjAuAfvZJ
vQYrxIlJCNfCHJ6CK+QIrAUPGye/+p3TxItJHjW7aLq3J8W73PK2cIPgpyOPT7jHI/68H7Pub85e
Wtabd523JuPRIRiJ1Gh2JwY8OnQioqcLtNt2vFWbMKoZNoNU1nqIJV77cUCkM0XEj+UBnQI+eA3s
OPA63kB/XvEdIFuDRBFPCjbd9e/ZoPQsZLOTP8nPhi4S2HR2RrWAb43s/s3Heh9ykfGVwsfmZ84P
FDIPEjfNCyXDQpJ8jasdLS3ebZ/sC/cvqlyYKFU4Nq89I85jFS0eQ+5Txyik2p7EwUjijhSFuNZy
PxThQp27vglQdEMU5acpLMMAVTU4BX1S3tNg8iruKYq5PvvDPcP4aGLY9e5hjc5VGbf1HeCVpjpN
N5W6WRVYdR0SNGYQ8rTl/zX6lhB5lTjBnoOjWe1mBKhWquyg4+jeR1AZ4txpQPiWIVf7U2KGqxwl
0ELsY6XDfYdCNshmDUTcWRwREwlpIKx044+x1LpXKYHcvKPZKp64OkbpgxSFQpnXt5gg0EgdbfGh
th3jN0i20OAP1bN55ILJtLzwyj6AQVhbvGYeqgCHQIpokgSynCf1jxhZMBvqslI+SCSWuu1SEdvE
hUCSi0vJPVLxKHJj8YCmkwSu4yC4Edtqbv+Lj0b4W5OIatnUXBRPWjoYsxlP9rOTN5R/hvm2Od6C
2ORiFSrRjfG+H04jmJUNhc58ArvQZT0DSq+pxiOlDGr3v3fq304GQDZHJEuCrRbjsV0Gp9zOgLee
Q3z/VhTN0S27/MMzfay6RNFrA7F1w3+V31gr061hYFLHC+C0iCzaeh7Cxh0qWiz9Ifw9a4h3AGC2
lFSXHQZ2uynJGpFGeaXJpeL5+u1CrPCVDYUrSOUB9X/QqjAJ25N7KPsBD1gUyujw6Ec3QXYNGVrL
XPwYNcIfeEueT06x2e+zWmN4mWA/8JPLsPnFmP00FGUEs2QwlxudySOW5Pn3DEJu1e6DwW2aA2Tq
VEIiAqkwKHSqae60i28J1/jtZij7I1DPjMqzaG9krKzOvMgwooQy8oyy8EDvVIsRTvVZCKvjeyLZ
tW98pgOekBJb3ubA5J/Ax1GtXa9vMlbbkdZglTqeP8I5TL2H6KSNJDC9xwGfDvoFLuXEtLDSnjar
YGecGtlRpGdYWxFAalZfBmUbPoDpQQ6tFN/PY0meeKxQlMcFYQVdtrCeq1z2WDZD10tDStRB19hP
K1yz+TJSo/1Nz3Qzc0aQBhngp5u4e1xcwugKg95W6KBp+4VJGp6zKLex+V84dnOd9hu9OYCEIUWd
tu32s1vc5XwbsJBSUfzDj0ak0Yuh+oQUYtC1sB0VvpQFpGy3hSHrw0Y8Go45bBVOH8uye1BtoZcd
kvKErou4h4VWQvg6T02SRTzAWEfyXe63Yo1Gjla94vjKGQFkR1pogY+TgE7Ar2YBi11d/vn4wdqs
AdQE+AoNjcg19FUZE7eOytP5zZHDN2h3GLhmSvwPhldUNG8OFYcS2geQ7W5HY8qp//jTrj2wUtVQ
MXaiwZAQ/5MN8APMj3c8Ggs2UnO1/lUN3YozXs/3q4NPy8eWaDL6UIzooA1QKLtGfQ0pXioE7R8/
HDkeGX8KVlwcDC8kVSuquN8Rxn20TgAhwubaSZAsFZCVWrnNv/wIy4drCx2jJzMtg5uMqEzIyg6a
Qd1vkaV/mzEKemYEEkVuYB+yX9cdW6tc8vYGhxFGkIPUuhNlrM8jQDJnYfuv8gVNhRqiLcD7sc7d
lB0E4GkeI88mbAnurvku2Fzcm4LsVX+ErtKKMS+A+619SPsodUnC9oTabcyxr1lYnOhX22vKOhm4
SJEMoGmOHvfJ48ZTj/au2wmYC81aQ0+e7NLJa4iXmtkDWkAKEr1aRUvWaqS+GaJ9CQC8D+hyzVUC
x0cCIRrp8Pi0Vdvk7SfVAd0bPPKctnOtpYRdlLZlqP+lFLIlSpAHJDLCC7sgYsjoAcO36Jg1+CaI
EDJQBWItA6F/NfuAZ+KYNTZHPy7L/2xzfX0ud04xC6aCTSqxA2sXwocUx+vDLC4l+TA0HoT7bKRk
QFrp8rj2MpPZMaUvAHv8u/wk4Ucs1Fk4vfl9Jwss545MHW6g6xMBQ6UiyGg7G3NXuaz5QSsaMwF8
elQ27cq8eNgci7106xU7ZCefi8oZpi4CQIhRxxJoft2TN4o/KtVmUBKsB/kIbGP7IcEo5NQfsLfR
oV/Ra0OBTkJGg8vKLEpwEWvoJPozY0RTNwPhoXxxg9Go9+ejzr1u3eY/vcd7bxqKmIA/xJRMFD40
L1B4dgRDmieOWCBSftEM/GCYe+PiAHnce0wDkq4wrz+GQQeQcMaLDedYv5ZOHetoxilxfSt27/rY
YgeQtH91HYGFXjr7g4/DqxgB5YKDB6GZnimcKpKDk+Ny1xDviXNhJFnjD9EYjyN9UVqs2HLL7gFc
SAOUtRwCyF3u5dcC32GpfIYT8svqzvw8w5vrxTENvUhDThHfBcdySPdnOGzrkhs93j3fHQmpXCmv
bEnX7oehR+ZWlqBNSIKchoGGZwzJNKtcwkwhEt3vh/LwiJkRSiyybO9PvJF3O1jg8t06J36isKA8
c/TU9yY+4zA4ZqKSjCOxTD2sLizoQ83Hcz8+ap0nfBJt3zOgdHfIQ/0t7AEQ+6Hp6nAq2oF9auTw
rGKCErqpKFfmOfjYA59jeWbnF1Mw84GVxWaMEk5/tH7xcmzVttJgi/IEcHKqPPUDHOVf0A2WQRVk
Hmx7xcqq1WdGzoVbrOHAv0Zx3cPbTMBriVAEsHAo40ls8AQUe07tbeoloLvXX0BQgQkJLlEULfcW
4ccOESfb8YZPc/heMTzBpW1gw5jR9clkUisY2NtMXpiS0KGea9qQNQC56+hSUK/XSq1hrA6yWaCg
9LsL6NYYvA9bmlHU21eYhaDE7wl9T3+B6qAhX75ojvO5vkZ4ljm4mdoQCX1fq3B/5XDUnPTFKfbV
myLsyx7k/t8ksEthFJGtvOH0KmjMv9A/RgiiInxtNDu67uVRPjp5CfboDuVnSEQ0Xlx6dUatQ4FO
VNwOqTczVz4CF6n4n/BgmjzWMkjLf4+S/WcIuuaRgLDwj2TERFwITHVvk5IEYgKGfCWu39OI6OeM
FzpKkQ/HoDGlqxewy0Pu8HWHc4ZWYPBEPCY7K+cMxhq8YpdU9plbUotnOQ8Ht8wNuvd3JO8bUbbs
eefbwLGSxkc2qTYrUiR1+FY/pKBwQtKRoV7rb2Ti8yybP/x2BhJUvQo4rTIfH/iRMsvkuwjN1tR1
Ik2clIjrWJxcKj3o1CJ0cFI1vm6JWP2Mxh10BnGXZG0x0pK4hCgzuUQ88yaxWoAfX9zUPM6qs4Qb
gzJPpysTijBdLEGYBAPRa/eXbSNV5k6m04wna+Dy25k0qxOMfjKZx1tc7TAtXNPG28eAlhRVVJ1h
WRW/qtrCXdbq9F2kso3reCwUSPExFn84kiVwlCK1Paytr0e+PmG7y478l8QzdwchBXCNpJktmwSw
qTFyKqMeDvG1XqnhRta7lsglYWb5+3zJf2RIbYoCLZBx1f+dyR9tKd/5s6KGwgJo3fiHuqx3h27T
Ipz20DUJ6tp9d0jv3M8cKRGjw68vRcZV10uRpRCo9UQPMRyMld36lTHdUxqnE/BUedwnSsl9/iYZ
/HSAZC4+gysw2PrL93XHOQ6yW3P0XOgF2m6WBl1OwpuaGe5ENiTeZONO2mkKKXloJ4ahCnOzfmq+
usf4RJRb4U6x6oqUgo4pb6LEcPvuCFuCVv3dwlwgYFq6u2OcgwFYphS+t9UFQlv2h0A4gSp8dOtr
EJ/eQe1PuRssYstpiq90Ri/UkKedTNR9Lledh/Zs47DfGsIrIf6v9NfkWHj4F8uZalzrpCo5ErSr
tthopiHaAaNVlN0NJIUeT2htuklB0mjCBuBzgCZMS6Z9tFMDv2EUxaT/MrZBTk9pwi9q0pCiw7Ks
HwgTUjJfPGVJQTjFKnroKdID+a7+vQzjtaqwge/YHrXNjn48wJiDjSNSNyJUhV0W3mkWQMgkFjcY
UKhV50YmvDan1R3dg7teyCcbTa/wIkyqKBh65NAmqCapD45fR3fdfFOhI+db3b6Cyesb5dAGajKw
+RNOX31/jf6QhshUwGtuQ40nAU+0EVb1DRJ2UKG4U7bFJrCSC5apOgcJWY7+DTqeLEKAj10og9UH
YZ4OmJMF7mMJJcC0COW7p2g38s1Q4D8AAAWRJzCSK6Lq+Hdgk8VDXgvhyT8dsw0U/YwnbcmOYl0n
71rMD1SkZmJuQCaTdqmXPXO7iXg02zK8O+c/FXfOzH2ICefcWKbUhWJKZt8Qv8jxhZpPzkKWOpeo
UmeYdJrDKJOTWpNdI9I9QBFBOy/TiQeUN0+jaEX1aQohUDV4aQAgcvBpfx/kNS6EJsZYig7p2p1m
0PVBMP+JTXsw6rkg3rJmv++UQMb/1g1RjSydbzIBsdTGnXLZ/jIfe0XD29RYU51EKI/3+4pvV+nd
I1wGabVlSGH//UBdzQTm0136sJl6ciJwp8pb+/6X2JYUOHx2I2wG6zVH9hPgVzriNVZHvFJtsb/W
lQDXWja7OpKkr8KMFe6gwxGPHnjYt4NOwl+MP6624vUkyvumyK4aH5I332q3PJb5m1uD2OOKbLkt
1PGk0+LCnfyisOzofiixfwAF9n/VANPHyuuSnT13hwc8x9k/Mopp2IySeAOOjnCCJsG3VyWV04r/
V/rDpBdJStj4tyk5jBy2jllG33aXeReKZB2D7Kv4EQqFsWw7Xt4ApX2XgLic1j5Yb0bdbDxxIEEp
o7opUnt8Isge7ewwjLDM07mJm46uva1W98F5wInpZauOloZv3WrvdRALvZWJrQKmS3LfIRcJykZ2
Zx9tFHEptbK+uvsjDaPiW4dmQbUzLVLf/HHXI0f5QvMfIca50lEUUTkYaX1YHH4MOpEUiPae8qmq
G9esJclR0x4vbDKhQP11D7PTPApOWBe9+M8lKBHR5yUjWhLIogHPRcCZ7ECodZgWL3e2NzE4haf1
t0fhDswB74vJodYHlZN0j0XjLgd9ltQai7DyKvwQF1oz/BRnkf/CM4cwP5/M3Iq81oGXXxZ9XVQw
XbF+RFe9R2zcfygiSn84yWaOxG5L5ybBvqFisFFH3y7C9YYD2/jShxNsRgGVjqXVVeAGWPndMfPv
q0ZKWArVMFVWMm/DrQ6sqZgo2AgOjJW+8QknkparHFDW54vZIJ3txSD+bwGdP84wcB+UXowa0unY
FJCngTzCm5Rx+bR+Uv/6SaIDCLP3arBSLYOJl73uJ9OhQIh70ARBDeutqEr0F64LI3xnDyN0DejV
9z95vSHplyp2hjenm99X2/SFIjijHMSORR7ABFZMHVxy0BrkxyOVupVJzSD5uH5r3tR7FIGzCaEy
QM1CMEq8MmZsdtq2mRup13KXN+t4LP/qLI7G4MHZLBCoCzRCpIwV+OyzlJwka0jAc+wUL36BEwag
b+TTHD8jpZQdcRpUoVyzuy1E0WU5BAu436RsKbQAq8Enyh0on2y8n1OveiFFxW9j5E4PPAA6YNNC
fl0zTNzgXA/MucUWIxmrN7hAr17Bz+M8aZRYy984OGEci/tFubZW2y+JyLMPTcDy74/j1RiJIMmN
NNrFBE2sI2sWPud2KPj8M18Brc3lZkkjdgYiwT7RXTiQxZryqkisT1j2cSZN5SzQ7ELtKI4UTITs
++hb2rEUkSOwbxbFTCyS7WfCOOpriIN7bZ77zP+XqhFsK+h84rC5mBTbu4eC341u+9h5w7KCIr+r
dYp3rQ0thSeZUrfsZ9di0ANIKSGf5nDsG3VGN6F4YuNirQqax8KGGoIKeqRSmRlodF/nZivrxhxe
3aYMR9scHhz70lJerKLpYRiHh/ygyoSWbVxZgioN3hwPRUXpdA4s4ovPoluuaLIdytJkQtAgd2k7
Pz7fkC7lwsCbePV9ZYHlJmyLCtdt0XWALHPDCMrN+13sd/yWCZPuY+e6NylbuI9WZkZT2yP+grE/
kcdGFsTo6ZN96aNcgZ47yZOHvd0X6jVxrPVqV0UQApstIrqGXbGHtikLUBTmW4l5+yi3+I2RyylQ
3SKvN5Mpe6dPeBE+LjouQDkEO6tdvfo0tnImhyzewp4D6CYVxH/wjLHzy+cU9e03CQSDlz/dXkmP
2xPGPw/C3cxSUcgiph1zWoEoEJAuJXrBpEyiITMDO7Qz7Pp2axbyIT4+ftlySurZlCdcYt3Ux3dY
aLzLFRjO+OdwQqloKo8R1chrd0rG0mqM4PRd2/jzlwrOe98WbCowGyvzE8vBGVn3T2bgQoFfm9IY
gpntsUaRQfU0kgd1N2IaMog5Dl3EdFQklx56DAq6+9CCxeqiZdq4T2aaAceG8hwxUhfE8vOtAjaW
ceh7Z6iVbk/6ndPDmOmstnjdF3giV8oV8FBHbVk3HUGTRIKV9J0kTRn2sRU2Vu8iQ12l7FRanglz
X+Qa0QyjjNMrtAYmCY+J2yd7Ha2A6zsdjafZnEF6P9iL4xsFCltaNvesJ6EgOgrcznsn14K56nxH
7PCfTEwCzEdT+VWu3xUuc9kmHXjorthnPdz1aolTj2mIUxbCJRUq0cwecmFHnhwqZ3i9iraYjKzK
NH30L0e/zZFg4nEDvKRoIX1J2W1fVthlb4fLvhvW7eZBfsga/JBY5qBLFq15lMVHwJF30HqnTIHg
Q9+f+IcaKYi8tanE8OneOupiYD233c4xZxUF5uPfsQx33Hrg1nU/GVYsW1/GvPK9w1puvSFSwERa
9A96gzAyaNDoQZFB1aQVvHln//wI7dNeBF3FiMRsofPxG2xoWEpGvk99LPoyM3Wyy7vlVWcOsYlF
xhyjgUKCrBXumCnTebjxZGjKp0dJFtOQW9MqByX+CgR4jNqP7ds7D7KqUsUqPOGDAhBkfXp+JJQO
RsXeVsORGKR2KEWqc3BgZKBVeQFX+vcv3RfyKf43tkyXsCT/KncAJjHh9a1aRuSIj5B6OyQPwNSi
52uFIROuNsd2LlgBifivLCVdfUkq+rLAubSVKnZ+hISP/piDkHYHez9vLxFAxNDPr5irj5siQ7fM
J6mpRim5WEWRB1eRNx0HzzqaK8JF+VXyeW2pXttWpL6xk6xVIEW6hSGsV0raEGj94u0mAtzvWqqh
PRg73n2v9R0QxuILx0JT1mlPYXf4ghqjCEVFm2qrCyq5kfUq6HgS0NEtb3bLss7L4KY1x3mwpvjq
y7Zc9rMcXy4c1KrFXcaWZbPmnMvFLBE1WwkUgbZuqByOewJ6pv5mlw3fmy2O5fjOtBCppVXtemi8
Jav6TEfLNK5yFLy+pqa/zxSwoSaNcsIlFhsg8/4wxwCew+mUgny/PooT4JGunyixpnbJDHOMpc1V
Zfjf9WU6/VXohgFTmDnJkaD2bEroQQgc8wkfze4bzdt1TLAXujg9+uMXGkah2Yyiv0FUnKACDC56
YLxEE5qgGtNkdpufFLXjuN6CDmBazBlrdA5S4BgDPapD+Sl3k5jp/msWl2xOSTBGo4/NmSLb0QFw
LVBw7HehSxokzXWj6dlWnqJik+vIJZVefSmTlYHuzPbtStuqsP3fIvROHMdsZLqpeuia6IfYQT8G
s49nEhikGI7jys0F/lSGhuWDFotjmPPtcNuK3ih76kPCnJ4LRwYGdUP0L9iX+8gXoxP4YPryKuna
ONMstUhLg/2EfodqGhcFUXsZciH0Z5Us5vPzTas0nT3T5uytX+fkCa49LofUlMXWb3GkyUCS4zoL
e6nCVr+WRCdSyiyUwaKoz/+u6A73d6x4EqTlih61uNqm7NmN63JNXFb7bQ9HCvsAE7s4uFaG/B12
x6MYRWTcmEnEFIrUn8DMSaJ33QGiT0nEKuuAnTriqOvZjqUYPWniuS46Cb0WT2JbI+iedMi1hYdB
RuWp79NetPlcZXzAIoAIPCXm8HbCi7g1+Mdy9ExzBb6+gvPwSCDpZtbdxPY/WU5KwRXAz7uqRRNh
vGUKVh0LZzdMakoZXDnTaTz/f2B3j+huwmDLXqUHm8QO2xa2j7Z0G0wp27kkcDI6KQOmkUTB3+x5
UYt1ry7zWQSNP+Q/lQr6uVzNXZEqHU13GogU0DiZO7h6FPfaUseRD9HV+XWrWi3llkNdNxZYwpCG
CzH/UjQXrqveN+4hSmvs/zuLPlhY9yWtELv+I1n6jIPeAqjMDW0fNbr1HnUnfGDk5yZyYn3D1TNm
nLyTuhE2HY3+/3FfwsDvtDAsgUiQgqnW90hxnGaGgHi//xXIFFl1hHdFOF8nFzLESTZRhbm9UGXJ
BlRoPGTmu/MS6eiqtt1L/stETlKwHRSPPo/BSmCkeHbVnpK6sb3RHsmwzYRbV1NbWE42bw8su4Pb
+teJMLOKMporw3LLIRoztbrPFBhnpFztaLeBTZ7nwuWNfMr3imbxak63sG/RTXoa2rATcTCVkQyb
Z5Y8Gh3jJGx8wImMh7c+WMF6rLGChr4Hxdk7HRHcyqJsN7l0/MSW2WW1cZ/N4tQiQX0cMMRrHhuJ
XsLhDprgJl30ZRFIVtmRUbZ6xQ9d+Qp5/kpFSl56NgZliw44EWm23ce4kvJFpWZbQFONrEdUoboC
1hkyEtkbf7SNyGPZEw/mwwmLtWA6Q/MAkqJUBsb4r+SU6ET7A5oWAFSYfVIedAYZubUwJcqVqCEg
JTq0/VLrLH7PFqGTmi5j2Acq5+JBFUgUT9RE1JjqcM0/dn63kfIRsMu9DzDCW50TDYnGKSQn3cYW
58dU7XFhyvWr02NMJgZRYW3OB8aUx6Vl+91W/2lFE3uVdhUGPiDxitaBUlFqeN8/z7OYBxa+EQUE
7+gu2QzLOcyupeFuLLknLtvrKBeS5kMN9SyIfQ7Qo3BI187nBb7InPdWpGIi1rtp/s/nZDgkgcES
etAXA0eP7L04H9jp3F1meY5upb3xY943dgLZfYvdVo3Z+u7/SafjtQO5+ox9Pm/jebl27KTgXH3m
Qp0bcMWgnFCps0Nq+kWoXX2g2ZEmgaawKzvr+iMbU//01dfR2qOrETR8vluhF/GWWzzlQbEIMniD
xG9BvieGGuVL9L0+RNk0lgGNR1udoqZX10CGoy2fZbiu+HqrbQ9vxsid60yIGvtajhuJPt96sBn1
poLgIY7PQudXaS2m552mDRuHSBa8YN0/LC6ChoDrQlUySgcdbCbmlDrUUBFJ2tBplKeAVsKh/qF3
EGZjCpGn9erVwbEwWzvW2VAqy1l6+2iQwMSg8SKSMW+axfeqQOIKACmg2cXVeLUo0aP90wFG+s3G
CaOuGR3JH9Rs/XTNupoQR5I9/T//HDTaZ8wZmWP4RCRnFtTc8u7/H5aLnEyH44HepRbgKuyfb6Qw
d1N2ubS4MzfDmJJ86iOBJQSF+c7LZxqRKkGDbX0k1hRt0rzd3FOMZDcxd14K+DzuxM4sNT7gSUXh
DaZh1rn1R2wU3+Vt1h+GNO90kImcW//uOoW5s+YDcbwb0OhMxedDbNuNo/hEuYWE4nNrb3t2/RkW
HuGupIxK+jUd+bwZqql4RNgflVfI+cnE6YH4pJi/5SgqoBRqSc5j7hkWCYMG/ujRFiTWcxhq9Byg
w3AmHnmQWWDcruqHhTIavjPtpRdDCZLPX9D6tIFU5ZLFmxbkobcHM10ria2iUYChCZ+i3Ln9eOey
pUxDwFOWtzJwzGttZ+qbdEEsqiC0WrJ/IiwuKeHZQVW6fq5l68GfgrXUWW4lbQf8C4fqfPyHiAEr
1muEa0f/So+cx5zULZS1w0Y28XPolcVd8YOKBL3fMPNyhXhAiRPPI/elfoBS3W9z5E3dpY5f8xD5
2gUEnHY1N3CP3PfpjrOZMuwImIRl/1+JrvrZC1JzogRCJ1PscayZRQqq+1pAhUBgVt/vuHcOYsde
bui9eDAf+k5m3y8f4pCIwRoF+MFlU/CAYklt95f7+uf3SWmugzkNjxWOVisvrZf2QZqkNUbprmzL
IS+1lZFCvWEexWAy6v4bPDa2bNwqkkiOBY4U3IH2GSx38q/DvOVS/jROcpepGHeTTLfA/j/x0GHp
V3DFr9juoVM7oS/yTFczb5ZV/fG04xWUyRYm1HA3X9192poYU3B9/uXq9tD/sKJxHqqGjsa3Rb6/
UuZNb7/1kQsM25qadMW9+8x+Wweg71HK50upBRmk2ns/72z0yX38HQQ69zgrzud3sMcL2nPUfU/q
DlXM68b7MVzaWRmavueDVRIuawzII9uahr+1gaQPuQ3El0qitRzORlxFG9imKbrhrpoBo02ZCG40
74W/kU0Xg2davF1ejbG5626B9lJ0GNGyIkK/5y6fO4PO7s73MmfzrDZvWvmX+ewaJwB3ACt9zioN
KDQBtGdbwuP5e3UN1yxX9QSylMsMg2o9UyFtxO/z6zZJjddUbioSkwshrSdiPSj8lWlUOvK6Lv+J
Q1MFPt5uS2UtFu7xb6HUD2heJDyIR5l3kTKqNTw/q6/q4+K3rNMDkN35/9+Y2IcSBzNLNdRku3Qs
tU8gid/eXNTbbkBEquYtu/jKLOS7JKerBOctBHLL+IzN086Fm8djULYEgLE/dosBRn4YDhRYC6Oh
OyJwp79vohseS6aSdG0QBgV/FGogMicOkfF8NQpVucUO7LyC8AacghQ1bYR7g3NsvzA2PIL8E5Dh
WtS1gobzdEQfK5+Qfnh22x9EqcLQ3DqaTaDyJgzLDDl95B5qcVW3fsUXKYbakFKfaRjwa/loWlL4
tOADdULxyrJnAGWbj6AaNnxxZmrs21a6gAtTpqrjdk23i8sQAJzNaVojl7JTa7xpG/k2wng5/XOe
tqpB+UCxoLGC96l9nZGNZf9lTeqwydlKb7naoPqqy6a0Lv2e2jxnecyLr0aXwMHulf5HkScCP8QA
KgXtoyePyLC4t0tXNCWPgiTRfLRVn8atBQ/c82Q+uY+7GWBzn+sQf7jFpJ5FOZ3M/0uGYkJxmS0M
+eKnHPyXtjtm2oPYs7mB6R2wy26wFnIjrNa/C0eXcjU5KnY4R0+PWUz+sYCH4MTC0svECMkB5UGR
AoEZY2QRHswlJbvJoBJV7z3v5B+e2zLy30yPYHhx/+k6CmYuYRwisCkXzq5SNqEapEcNRbUa2KjQ
rDAcjPyzNcMJU8g0wsMSM8g89HHxL/8RVtPiUu6iqXhuefTXaxzfqAN4fzQXEJ4N9PnvdGeYApZa
35XtixUReGh7ozlMCp6Lq1/jALDE7MMlId1jqLnIY2VXSw/hlkOAKcB5RJ05AUSN+h4nYK43c2M5
gQnqYrP1z/YKQDtIM98QUdJcmrnSiLjwH7JnPdWUWdpClAhnuv4++1vWqsDEX457q/Xq3NHftS7V
TBNtOE2Q85x+WPGTjMetFfIuPnVaD+k9Z4S4UvjmuIsWOYcVpQ4Aj+kxQ3X7+74NYVX4yCrtdzpw
je4lW3DB/KrTLswm348HysOvKAblp3RTdWu836BOThTWMFz6wt4wY4nnBRioCniphiEGwRgDB6SI
Z54q7H0RKLV9wopfkWNGhOv0x8EDlyyS6on3QMA9vT1sgvHHz9minCrfNJhoa0YBG9dVtyZ9vGkc
8CdGtc5fcKuanax5Pf1QCxNIDOJIdkHifkmgc1JqtWfPQBslyTTrnH1QK6hg94YgmS7r4Q9KzYsS
vJC8jEO0JzyS0au6ml0FiNTU2hxLjrPJh0D7z1WGEcj/4Id2pVQlb4mo/JwiNbM1AXLYV8YFphIw
D68qfCZKvdxfM3rnjFAFJtJ4MYm0IkZTlZNk7WnQRyukBnT2pLiP2gNWZgAVZggs2EH7Oaw8+gzf
PcW1+LpAfWb49PZLZxg66vwLYM39IA6DjZKpvuWhTd94mycTEOyZ+GDIjBptSRayEumGMdjj5sJ3
gs3HarP3LB+TUdJoK6EA8zbaWPa3arRKnhk4MW+iq7EIMpu3JEZv59N0wnaeB9H4oZVe2jN0Esjc
nvSDVF0NYbdNpICVnR02ReMwi8S7b+BilQ35Tpf+yvEpMFyb+3Lgg/Zfayf4beyEyZ02a4GFGYRK
xdNyjgFQlOxPoqA98lYhOSKoxYKvhJQPFpaRDlqrMds+70R/CfMiRndxhX+BFm4i2oajBuHM4qUf
GOZexLlhkrLh/2L6I+6Yl/n8/CZ4ybJzLGBhZc5bIrItHGNxxKRFbOz8bNTOrzEYBrMTplDYQk8q
mfzqFKxuZI5j9DNrnpATfH9v5+i7+DgUopg8RZ7bCptnF0fOXohBvdLedOzJLAWTbsynJFpphSJJ
KSmWXVsAuoX9NAegFx6xBHDFZPaDN44T7STTFOBKzoEJ7nNvJ+b11d46aKSLFeUFnqCV049pb0aU
XCzxNKQgDCCzoXyzX+JwMPUwWSrXOLqUBKfyoF3DYJJPqZ2cfcHyVnN6OI3eijxkpe/PzJciJh4e
nH0RsI1oo1qE5qTj7PzuXA4RcULG6O5X7v3EGBjjSZ7OIkWc9w6VLg1b96VVA4EcWJt5C60vfrRR
D5ZZReVVYpPfXb1bhTg0kYofp4h7clPdvLaINFfRzjZjcGbdQicUGewjDan/mLgfgmKLwVHMwKTt
xzPqa2wF9yRKfUQ0KL7BMiV20MuWljWpYc4Zz+k/6Lc/6xc5OIeWw48ZwY1WjUeF1aK4CIuUQkrY
sdrIHhyQR64c/cqAlqw3BZKIwYPvU/1oYmvlBnBP3kfzSYDYmPda5+01pbuiIehNcWb94fn0kKQW
tk2I1vBHZbM3vtbxxd167b8wgDREBP4+o9zU320Lf7T0iepncozAbXfRzu/A0zTnEyUl5xedkp7G
SKI2Fu0MJu+aneQ7Z8OjQuCnpWQhowe5oJ61SDB776i4omhIw/nn07VcxlrNEIAnDSqly0GGIvsv
EyJ4rW8rLw4qjVs3ptOewnOkQVWnZf6esS/jSuaYNVv8v1c6GbiYUgv7yf4oaXotciAbqonxCHiX
PViFf2zRpIlPbSFxcCKOFTIssiHT4QygElneP8xIvkyC2RQ5mWxaCRaO4PdlkQc/Yepztvlacwm3
FRiL3/EJ+WdBWfs/fNgQRPqDpuqSxGFigL/lJzO2nmQa72RY7EbKCU2Mfpjd51Mo+LsIDOt7afhr
HbP+WELMdA58zx58LCY95/ps31BzrCUhC3MoQT2HpzGbg4hOVFJrSj5mrf5VdmgEuDlMdRmyxPkE
c+1YrJtnW4mG28aIB890Iz6vAwEyZ3Mgt8bE7Vejegx4mVGJz7Grt1RD7s+0/DIm4Xmx2mejV912
v3coeyEx9/8V1Bq/tejn8hnBVK4TJKpR61/kkLHDTLiScWS+TwzkirJc2KlnxPvyKk1eyEbOY3RO
iPYZ+LX3SGwIkTUQeeE3ioDiElfbxtsFF2dt7BwTTqUH8qNCo6ZBQqf+W/ZPpmUwVCT9FVaaVpCx
QAPQev3F9UHRSwbrLzWVUZviAHoRwdaFOjf366xV0oDWnrL+7AnJjPcl99pnVxY+FRtf34TtdYrJ
WE/r51ZeDt96ST/9rpJUA3hIZmB1BQ19Z818bJfo6LRqIVHzs3HvQB1WLkZCydBJ31W/Av59qk1+
b+hR17DwxADw4UCzdbokD6FODS3IxSUQUsURT0y7jnnlzV6pyUua5vb85uP5xoUZrScfpja6U6kM
fzC2L8nmFBgj5sKOd9iIDFRBBL3yxtmE0pctyL3jGyd0rApa+svhsr5kZQXwYDYNlAiSfailXise
508zp72iRwTPFGyiL5sLisX4HMVIjdTPFZ7Y3GElMt8YIWKFuyg/3NQ4/dlcxa+84KIjdIT8Pc8T
IQu8+gZ3269Ax9Z3EvFmWAQKGCf6OH6909nFyrHUAy4m/+m9f2PfqRD1OwhuZN3oIaxbC3KTtBzi
6dUWu2bAdxE6rKcDY/l1GQs69Gd2UPuUOd7fVOwNHdDoX/nazVT12Tro1Wg99lmWoARXJNjlQbLh
lwAZ6UmzIs2P0tYma1aOOLhKUI3E+76awwGg1ypJAYLxtdPEdHQf+NlqzY4sszQl8lIYZRUZKq8L
9RR4+q9fV/M/q82GdHigZ025L6/nLnkyzKb9HuP18x1w4iu7FZTFeRIWNkLHvSjo+Trj69t9Wa20
qNMvRaRiW7yBlOzjXH9SIR/ebo78V6dFkCPhid7/06hpe6s6eDdnA7UKXaP7hOAedTulYG8XElbz
1SPsRS+EA3HOZInNKOoedXVHRM6epz0POI5sRUKmpGR/oVt/jN4sVDQcYsmdZSTCN7zlKX2xQkEL
GU/FneTm0xJEQvcH8XT/kKB0oGizh/DecDarYUecer0HOTY6iatbEOtu6FE89jrCoAC+FlB3ujhF
2KJiEbgFUP4eiaEQalja44MTEcwnaBy3OOkW35I6CrdffSk2u52QQJk8EwG/YbbwqNtHsO0qR2nZ
y7Gb2FP4aIMghlotqlyEtnMxbYUjg+CcEvb5Kdr30zcEPfs0+6o0275GTqdTt2e1DJF/8x39tziM
wxmvkotjd8VIV4rRxDmuo9KM1YhVaOoPqmB/A96UaBWWmXVcG6acfpmymF+J/qBsJuVflBHTQpBe
tYWNXKtzWGAFztryKHfnYihfIFIPKKS9TZhs85lWGsfGBXvl3yhiU3Liq8eZ0gHl3NvGI84/MUCJ
7oreLw+2ERnqMa1757wjgwzrFjvOvFLXGGy4mqyx1tv3pYRe+gdOrYHHDtmoLf9Fk5l1T1jFVHwb
74ol929tUrpx4LEISpD+IJdSydXEVRxs4xWoY0Ll/Uh0DOui5dFH5LcDnAn2OvK7VKWd0/P83rpz
+b8uWucTBsK7MUA9NidypkNCaYOg0VObiknpDh2SI4CaaB/D6qB9LxxEVKn2C+yYLHo39Yf7m9dz
sdH6YUDf4hBsCUAE/S4nSFBdiKMn+LhPCwuUm178jQfcmvmEwXz/DjDEjCMOjs6v7Adu8QREv8wl
sGvZasFDEQ2/2WDHwm2a4objyqS5+GezXHugBpMIhA1ZgeotzERpikw7B8nrHswpcDIOihAggqn8
ENoP3zaR4mqO1MVn9QdGRctIzQF6BZAO+O+eT82+ac9+5ozU+extgLVJYFZTh8s3HhmnYGqsS3Il
rahs6Nhbolb3ZLmJrmPDFZ1rjAlYDoTVns//oMKVJIiwdEq0XddPHdFP/svoT8WNGn0EG9OqYtO5
IejdzHL5u/0Qgv3pBrm3ktaXFs+a0OJEtIdcDQZIgdJas0Do+1wyP9V0zNpOEkjkcxiao4xTGI3R
yXJ3g6ijF/8mY+WuzMzpYJAyLVm2usP3iSnc+wGmgagGNBxaFC6euiHqQqZc04M4cW6OXUQ3RcXk
OXFw3yF5Ul7eRBN4ypJGf2GOgPn5CGgPeKrR+MXK19z+RSaQKKGz8MlWxWOxvnB3nD3gkM20SjPH
uw1H3GnlR0fB3ddLFV0AzUtqBpKaBxGCzsX2a1xeU0vFO8fGqwkPDTJ0etBlSXL3BXhMkYGRghVH
FC02l5FzLDD4rh3KDT/0krxO0sd+FFFWUDEjxGy8eZ7kbNTFTLE96k+Vsa+J0skEVMPbnJqQim4Q
aCwVL8mZE2G4l7zURDoJ8jFsSEtJI7hVlSP+UkDk33av7le1dAKTdf0wpEx3O7s8pctyvZD+Ot8K
bBRXSlIeP0ZHaKDJa8IWxWzhSfDjIB+VBM8sE7vFO29V9xkse/iqmxZx6AjdtuojUP0vw1A33+JF
U/ItlAijK9SpLkxQHQFKvVkg6YffMUQR11tKXHFR+kfhUGJq6zsyI0RFTtt3f7zRFtk5yX5GIQ5N
UXSfRND9DVGb+O7ZxeXuvuekuXCe4LqfpYVsyOU3tHPPZ6l8uJ/uAGHr6uXsxWgnLEzz1T2XTvgq
ERPA5ffPBQ7TWE300Bu/ttCL1NTmg2mYDeYUOiv/vsNyZlLA2aTfRQMCKl+be+Ss2y6JUXE16LfT
fmpsjbErGIV5HdlH8TfYKRF5Oa7cuEvOk4wJAmqUHue/2JQW7SKZlph9WDCVu9x3xSt+oWlBHF04
4WCSrlZcdwQzpWd/hcbHkKlklwFrcx0kOdjgvbNvG79kiRLQWkkNuUPX2o4ZgyByAjDP07ZhIAbL
+SA3XDBYzmXVt6YIKV4YbrT4AjTMNg3xw72g/r6FRY5g/XTnT7IJv9AWSt+EVdGO+Ll+VxaM9Zqy
vnf6/3q8utjPCMTX1h3F7TaZ+7ChyoPJVvphcDvC58IKUHA/qY+t6nKFOezkf6RSpKJ7SgNWMLfM
htAbuzhtcSwefOporAZj17wu2Aq2qp75BLypt4N6xlPWgHtAF/dyxbCLAgfOiZ6SxivhQiafkFr7
m9lJRWFmO9ggufJdZdEKSmng6H2RlNQuXOH5ehCr0cQpnv6SfLoQ67NJ77U+GFnIQhDdN0JOVv4A
TxgjeiKiKG1n8fLT8918gy67cypVgqrWeDYmJ2x/ivBQsrBUkui7yhI5hv1SRdOL0HJHh2IqTrv+
bW9Qhkz2d9pM2lsOwFhAwmH+zjshEgYovyxjeKhXponoIkBQuGkIkh2l3YZIt4NbvkkLGtxIARI1
M2MyDN8FQtPT5F6zgyRDnuKz3LJIi5r/q3FYJ5nJdf5Xa3piECNOuSQkbYhazjNB+KCeeqlTr3iO
0d5uTF/HBodrfwyOECw5Kz0pKKBZMmsZM6vebTjOjNv2VcQb1pwmimAvQ5OlCeUGFjZtjF9s9Jp9
hBriQrOODzsgJAt3P6MSp/7tuQAtfrxd4GkMk5oq6hjIXml00UmZQJO6Fd939224eQYHfY9vNjNB
imPdBorMhkN5MPewcOAGJEAiS+dNP5L1fFvf4pkZ8aVUVC15ruopZuw9sLZOXdEniEpp1FRIkNaF
Oaq/jI5kPSHxS/NBcz9ouwkixP4uy6srZry16QQSXc7MQ/DsjfLqGcfGX/+AMNwGMgtfpseRfYse
UfgXiYkALdAttfFuSQjrf6EqorXK9qSI52QJiBAurHb1ZggrwLMVyruGG65tj8U+IK2zkJJ/MCwf
rpoR6d0RHoYfpuuf7iq+vT3Pt2F5ECKMKk30e/HlwPOvhBWB1VHVVqBXS75EGl8g7Vq5k0TOjnAl
aChMNuat0M7wsk7dLJpz57KVGVXX435U6CFYBC1TY1VMEECaathGybOLxj1Os1bfcBX+ih6zY0Wn
yiSBrkdv9s05v7HpGLVMewRC6zLD2vNiRZY1dAR2s89uQv6V4o4p/kjjpZzvUtvR9f1k0/79YbF6
739yNyJYSwPBRJ6gmqwcSdxWU/rRT9E4zaYxO1xGnqpwMbCI9JBU9E8Wz93zzYDoGFm2iEOJge/i
eo7JwYGTtEvrQTAW4vteaGwKejAXNno5o+A1RM/LubF6kUr93/53OdybGrwcXUvt5L5uRvqs6E7j
zyRraMFTA33pZnNIeqMRmLcvN9nuz4Hdt5bNYgIpqHe05t/pXFT91kQePMVeuYVITHZvYocqq6VO
EaBhfwc1Ev4+kT5HLxQkXGUowSRSU+J8WtXHadXsK9p5srX+qZ95aehQuZvhjQUliV9FzbtOZ/9z
4WlbAC2gksDXmoQtsCmDKe97MMqyZPfCDrRPhwPp/yP5wUOtZ1wk40Kfp2fJh5lbEJgfe1WohA8T
Gw68Ja3QBuFl/Wn0OyujhzcZey8aQypiB4hc+yIncB/BLnvavLksAwH4sjOU4GNL+Yw/Q7eD1ihS
zOeQxqMxrl9yr9OriTSgecun0icR4+QP68VvuWfnHh34kHOL0sMEqnL7oIG2qECGzbwd4qCDc6yI
VRAEdzmB+CAHt1b9pLAkDkHCseZw2zIbEWLxo1QCP/6OHlYBDj7SGGiBFGy13QOCgk/iijeV5ka3
fJVdQY9UK3asFfz7Kdour1E8cP4SricQ7mRKKiySkMUAk25Hnr6IpLm+Uzzw6ztrHgSMbdcCJ8wt
7q9LbQQu92P72tJjrx4F3qKBayzMdPvSnay7JvIyVPDQ/WQ4Fw4VkDktBD1wpFXvLiSrID9LyzOp
Ds/iuWHVhhmN4FC2EcpzK/QxL+53eEAX3CWUsLTFtqZYqMDdiigHLe6LMmYtRuwyXInInBWpIDon
vqifYqnhWElg2u7Ocd5bEfP4h2t+er7IC7xms3wMKN3/3oVWmez2HDLTdS984TKpigsQ6FJhP/xU
hx0U9GsJ+l5ljJxQKRk3OULzuucXU3F0ueoDRx2LsG0tkEYPGtuj7RQG/QwLDLqIt8VZ32xAiHXL
1P12TWZMM4Tu94+M7oxhYeFnrV7ruvZyVJ2M+v6cyRwstzjkhQcy7MSu1zEradqzwHR33mGBRVX1
97xRruGJfL8kUn9uVtMpp1ijmTqHk0IijOPtZxS2fCmEFF7dlUWGmGj5cwnm/fy43LUrQbyXS10y
G2FtNBcMMxxbGStJcKn1JBag77D1lAeXXXeiHTCSeuGFGzDZ8UmNKaMnkocFHALeS2ZhszLE8X9A
uzUgZKv0kAEKrQrtib6gY4SWbeahhw1f3wdC1sszQdG0g4M8FKHIwYbJErI8UIb4Cqnh8wMzmDdu
YlyKECTFBckn3hRfWGFMHrsm+bu1AGOJNdxBvBMDSfQbYBN1WgSYQKjxyGGr7Kdq+Gk7Kt7n6nKK
Vh/CuvqgkYgAR1pNsPV3Es4jSStVZjwiqhymsA37t24Zb+XdB/M0AIldqsGkUvJ/EzTSqe5qqFBF
n8jwcXsQKQE3gNWlgCa8IDiCgHFphC/HJxn32dTPblyJH5Sh1DINhLa3feQaxjKuGHEHAgte0S51
uU7Xt9K6zLBa5EoGTehfYkHEFkoF25GaZA44OCc7d1ERLc1psFMbKin9Azu54fqUBrwQUpOgezc5
I4YfyxhgvSLfo/hR4dAkgtuSF/C3H5WWqJgOGOsMtj72c2P48ay6bQJI/oc59KGMHDhy6XdPn0pO
XeT/cAis86SzJ8aGxVFsqhiUplk3SUfp45clU71LEKa6/X3hhaL+JAIyJ6DFAkBesD7LMoQyNE0l
3Dn2MwF6yltdN0y4ftKKoS1LftdJGJdHUHFbPocL+43tPQAas01RrZ3w4GRoqm8yaI7RkRJ6f3TR
dxHZjHfAuW86ECcr0phe88BERQ1701KvZTRLk92M/Gk25YAOyEJMnNDC59EWyc3IE1J4qcpctqF4
bRUBKp6TCcdlhBGUuRdHhZxub/0xTtNK7bNxy5QFc9nisojL9tZ0j8P5nWazni9ckUAA3XOy4r0/
YaLJUdG80b+8QitkTFBY9Wki2kmfndk08NnT0Bap1ktFDSQDAQGDR7Ml2c8Omse/sYqDdT/W7ctV
QAN8KoCVrz1V/E4aWDXoXpVAo2CwIpZR32UYN9CLs44nm9Ot1BFPDigLKLRxScQq78umoDwQ1R4g
k+iDoiG4loa7+jpe3bqymhMVK5X3ZFcH1rNqIja2dHYj2hA4/wy0jB2UMoFEpg/KQWqlA7T/vJAa
mmpaDJBLcVz219H4S7JhjbDF1wklapnN0x9eX5HCef0xutCCDUo5TmqYXXStDT52147GUJ1rhmZh
wzZxGJRMrxxGA1r+I71WdmLp5OdeOc6gWwBq3EpnN4s+UIFKVs8MhtHS8U2x7tsphSANulXPFqkI
sSIc0iMOv9JfGYhZ+IkC90XruPHMZsHjw5NJMMz5eSEcNXx2dBVV1151Q79KFyQkxi7o+6CetS/B
9D2dddI5bb/QNzDAjywpoCXixXYMhhTyjR3D79IkxXF2UFGusRGBqcL94roHEUGDbYYwuTmQijBp
Qjxw+wGMYmHYCXnauIyC58Fv/Xj0jN0yMSuRB492SICIfqP1gDU9fhzFz/Qp9qtml1mlaedjhgzq
eQEDl9iITCXckBm8GfASLSbzNL0UCyJTMmQYxlDOqcJH3/GT9CU1wOWvesrQePToR98kKDejeVfI
mVFkfUZGjSY+uQ0sN7Gobud2shTM33s0U/hUVjpv/Kf8R2gs+GZ5fI+KreSJvvtaDD1j8D46/I1n
Q7NY4iGedYWuVvtUCJzmd0OVM/vz8KXlrp9yhBQOu88pBTfo8i1V/XQhv/0VWbmX3s5ES/EvLFy/
+29RdNYxRjQgBlfy+ZqaOWwx62V+uTuWTmrDYNUujpkGg30Yf2Z/U/lh005c/J6St4YtDN7fKCYv
QDoYyWWWTtrhrIzeixS4UHI+SKxAsK041xkCem0DofddGoubBm2i5HXLxdA4YK4FzsG3HxQoMlD2
3pY6zuei5NKGcDtZpYgG2MAu2L/+EwUGX/U0FT0aW3+3beBhoY+URtBVx9tK3WgTIsD8C4gwUPfo
7IXFKKt1kHwtEtE38Eu8zqQdg1yKOVuZKutB8+5BeLDE2Q3jb1crfZGC2e376g7mL8qxXZesIkVj
OJjcrwar3s1AhySdojODV+/TjKQLafJ54ywbKXAp/RS6vViGvySghUOtJu4s0U4cwudiv8IZQGWw
fHb1yUPC74WI8IxITTROc2g+v4qaWddnHRAflVzzrUrInSZO6mIrrVftpmS9EyINw8ge/6BiO5sC
1lHfkPytfssjzLFeM3mIH8/eClkxDw+AYxJopdJt6uX+UcCbF+3OASTaYjZSGWSEXrEqEHNKQlbU
041KsGu4r04ikNb2tNp3Ia6t2aXDXY8BDdXw7rg0pwNClpmIkrNQjIrmeAFzb/mQBusercbsyZiY
H6gQFfgJpU9qfxovBfvzSfAG4KP1a4JWRnKNySQJq3d1NJzVNX+5LSv1pSpEJfklB9jzPrRK/skS
uM3EBMwfSmSsbzLPLwfEYrX9MnG8xrROfi/VDdBVBaZvDn+SNgzHQqOcNkmQIFRefw/j9KRBEwg4
VBp3ryUVvONVh5XajOyiNw801ZWGd7hICe3W5x+1P09uAXzWtdOFbwPwmPkQ1ViJ+gXCwHPVIOxD
Qpq/VU3YsFRdiVyo9kZh4L8jB9cNfWBy2xI0Nl4s/xKsOXt4lEwzU3cgOsz5RYqF+2j4LaariM7E
PvGYklReGMFK5XZ64EIkKG2xcWH7VveYjLmN3AOespfeUdsWYeq16kAn9mzcPwIJQbWvkmTG5lmq
EPwm1thEUFQGAZF9JGOdKXjsxFFaGItTyfhy5OBgVhOmYmqw4LthuEkey6bbcBccYNYiq5Xgphpq
mCgB4gHDH72d9qDDgeFsDk7EI63CNV3KzX992/IcATirjQKCgcees22SXV35tbpjaEtMHb+MB1Ep
Wpr90X9hPNmb0b3CbsaySbwhlH/CetgwtYYIpQNKZalOQ+cRZvAttAvTeVTCIA0iY76SiJJPWFEi
oCCNRw3R+IZJlzwhnIxo7vWu3L4JToVJ/oYoC1SJBy4rPd+iX4CsqdICsNBrgPFXkq3ZKxPHhvSR
VsLU4r7xUcGKIbAPPAYtoqJtG8J/QJXiRiQwz4m8NGcFEseGJKZhX0Dfg5saA3eT/XD1ebfBOtmP
Pi2Pdv4r7WHVBrzD7QA060kHE7P/++y9Mi/YBXJTs8GRVV4P6iPu3z2J2kdpUHBLjV/bene0bkex
x5wJCxnhTyMXiPvoceBYTPQNdOxH1z0CvJGhZ8eXMluGYCzUc041jaHiX9Kc+vYdOVF0p7z2SMgW
6+L8eI06Ge8WEse+00IVx2kP8U6cl4CQZ490fl3XkQf0AnHuRC2mwrglema08i9u2rFGmSAttZSM
DD3i8dLSyxgNXp9W1x5K1NGsvb5p4VS+vE9M/dQrCGTrXM0zK7eGcM6SR5yNBb0FMlqDDuNeihBE
ZF6LD64KPT+Xhs/9afIQ07gTbvBmCw0lm6XQx1dn6B2ks9t/BgDvlc5jhayGAFlzSGAYkQ4dL2Ms
yWGrXEsdUwGKnz8F7CaEZzScG/WGskGroTc9I5mALKPATtjRNvOOzMqwQ3dLB5UqHn+BLwTLUQgx
ZSQnvX73VHZKmTYATyexfQ41M0YpspqMN+H+SHZ+WoHeG5Ywe7dPMKc5D4HxEQvlSkHvaAg/TPid
bDuXxk5LwgFyIQ9nQ71pPhhS6PZIGl9SbzCCZl/kNhQ1imF6zooESDSo7xKtzomL8WbtcuaHpOO9
3KcIfSoeqKMb7ZafvzIIfz/me2AWeU8sXlmatMdLi9F6Bu2LvIQGmmHPUob1JsAnw8Ec2oZs95rN
zV3LNYwnyu1SAZxDeAq1aAYRtXQw9L8c3tPEeKWpu8dqRogzhBIgT2i6qLMRxWCNbcDz/eJAylkr
v3dX86Pa49Dk1k71Q0KarZnmOqsS+y2zZazZpoF8CGr+W4kG+yB+8sis5tocs40KrK77BzYU/OFK
RFx5tdblMCL2qCRnTb7JYeMw48sT6MmpRRm27hD5u6WrlntPMmwOV+qXE4ePeeL4cIpc1TwWN5TX
eFzRvFjAlSCDkQMKIbFgppuwIVxmHgtLTk8LHUsnp/21ljBG54prPKrwAUkBFwQ8o7Ah9c/sAVZg
SDIsPiYnrPYPDq/8psJan+/RM+OIHxQoypkFxaCZpb/pP0RpQjg+X1SrphDGjvzpkmMe3tWbS/Q2
l0M/i3uQ3KTnapmNUFCy97agEdRYZHpBKl83cSXaWVAGGVwAEgfm6gkImZbGzKawzA/E/3XLyio8
GNwymCVdwqIAPXfPX6Q1M4VPZMpcHDii9RVa1yXStuss3ieGzzx4c8NlMCwNV38GAzd/NpPfHJgk
PzGw2QlbgRSfRRLa9XxAjFEhyYISutelajoxOMuYAnKJwIK3TGTXW7+zBp49JMGUdAG+NKcqGwwO
QBsrDbw0Rr4xzrYXzrZY31Xu1a4geAAG6LvvqJSabNBQ3coFBrrPt1hdGynO5Tkv0W+0tG8RNi8Q
FmsO1Fz8s+aYdQ7XzSty2WahO1ZcYOhZF6PW/crOGC7m6OAMazWwQTq5MsNxiGCZiMXB+C+uUhM1
ilOXqkxK+CEsZAm1Idw657fU4GnAtTlv39Knzk61pYi/jkU88SiOgwRA1DFRa7I9QkhoC4lGTagB
JI55fMp544Wb0+N4Un4y3Bz6ZIsF/toHQPcIdjHwybPECXO1+6avjAVMBrxYbcVLDFu/SFYYZf1K
BU+UnWR8kBvj5278cA+vXs0FZQHc2Kew1M2ua6/1++zxjPxHMytkq2a9FlgsPQIL6h3tgB7ZBPpS
clWwvthYIfNw1WZP7SMhxyqlVeMh2cMT2R24zIk8B6Mb2A51zQyj5PmPvSxYrPyOwWOPvauEu9Ku
3+AGMrYTZ/Bdt1d2x3bVWF8d+U6+Vim7c3Y8uenBKXRyv7xfVpSnhjOml2ReDVhdQWgz3dU6KUPa
3yLnG40+VOdFUNSg7Ggxi9JBEHvWPRKZ7UljHKlcaqYNNM7YKy7LhooU6S2F4ybbxH+RKGMCYvAd
0jgE34SOGPkpG7q35A7/gJp3iYck4NMZkN/1uYa+VHOYkuxrYjvW0uirOUFVlSuX/DAXBl4AEUi+
rWyyENXcbEaZ2pakeQYmIkG8/D1SRahTbEgMgNIRGHvo9J6woL99KURdkG/YM4O1/J0YCy0mJyfG
4xN1sX7A4DttPEwxcNsEXurvJ4goupNNjA5ld5J5j2THobx76lASXiRebi6kCS1yfFpRs6kKpZt+
tNWph8OThOiEjMVX+RK7RPJKXf/s23/bswq9ngcNUO9Ge7P3gk45WPT0YGIyH4CtYFjHZQGxvD2i
z4VBiunxNpXSrCw10ZS4V2akf0cHJIWmuozYrHDX+BtxDNxeXSdzj1g8C2DND4Z3IqrxiAJJmfcz
uqtzojpweB8VUFSAsn7tdWE00/7tUJ9TFoZhyeu2ObUCOORO4Tai1bt7TvzdCLGZrZOEdV4J0UlM
x7C3eRcOA0RcyCuBls8SQrmytCclYnXsYXqVlDAnM4hsDILWCG0kxglskKTWszGUR3THbdhq6yOS
aTC5wjeujMpjR0/wy2UEdZMysHm/m9epSJoVMWMBeENCbt0dgN942JGZsRoowQ03YhHxPAohN0g0
BBbOJr4aSuWw1EkHofs6KkNTv6JclgDSqkqc1+dOkDb59TXya6sD9wWeWmu/BmZ7pNp8gU0fkji6
JVk9x5OuvS2oWTscTcOnX22bgshAFoN10Gfh2Z4v0L31Tl9DM8zEd1bmhhkmCf3Y/k4JpiMVp82v
W2TQhXF6hJGKZIzHkjiMycJdMCP2187MmaoLlJjw5YJiT/uCne8N/DXrfcsTn6PU/1aCMRPgvmXn
wYMHoo+H/P+00cp/3e8f99B5U+qNkPTU9Yzt7u+wjfdD5WW16vQl9uO0HoZ1MeHThRXOPpq+JSeh
dVaXRcXStWBRs6Vbao2lleUBopaOksBfypxLElmazAZTSVLCfzY/9sG77o0yHtfLbUiTOdwdJLla
ZUvW/WlSdv+kMAaavLsdqG4K3IFijE9ZkGbSdqAm436vLlcLBPCZB2vbvvyUhjU0gMjqHAzZSz82
oV7F9QtxMcdBmNeve26Is+cqI6o2cRxQiXedJD7YOG3w/YUP+No2uBUO69Ukk7qSNi05ymZGYm+4
nP9EG14n/PP22c5rf9+Z0JxpmZNI0NNrBCOO8LPZjhr4NQcRrd7gcZFO3JHvddjOCWmjLCW6CcfA
MqPIXl3N2H7LbdZH5Z1A8Wv358THnLQ5G9IRAru2Mv0AvDsk4cvp2AFKazF+zxKZN3tHacfLP/nG
ScHma3cIvEyVc7sIgotqxuTVqYQtnfBTuSJ822lAjX36YnVsH9xOd+IW82RC8gumEEdA2xlzFQ8I
BUS0REv7KQMM2SFhS7MpZ60xS/3eM3fzDegLHUKY8bWmDtsFej1edByn86/oqqDSytRfxVHNiw/8
GLGRyhjNOqFjWmZz9PVAKwik6/elt0Qdmv5zcuU2zaUZl+BV8Z77rQUxEumDxddWSJJhaWQf+ieG
10SPfwdknkC7IF+tARSpt7i5vz3phpR9ASyE8dn1gRbKJet7/Nyi7M2F9RfQMKKB0SD/K1/iv8OS
PIjn9uJtbJfvuXKyC0TAcsvzB30eiKdSRgtpBcy+yb8dFGBM/KJO1K78KwN3k0lVoWInneVqPH98
xxV4Jgyu4CLqP0qgSZjCyN4p0U2HDBkq0BoEtKOV8kelRM+BOgWrRBPVk0NEg4snPzcK04TaBxCo
gPHsHVvUvYanrydZG/d1DnJcGWKZkxbM9fnBqrmBWMjAPSgHJ3MdMMWYWniBh5mOcp1VRvq7BNrx
AyVydYtpzNP6k8gjA8AT7OsalKPAsNu4BCLZAsI02QvUwWQSDPcOGuVvb0m/+SbVlk5r3rwNbOGp
6yB+vdFOKLBpUWCMeW84Sm0DR4XMnyZEzYFP37oDQAjAeKxVD6T/t5rl1AMBusTWXV8qH0Ixk0XE
tEWXJQGouKmEtDKElTuCwtNFSNSYwBsAKZdztgMgVDs+QxJ+23DkTtAWeCgz2q9WUHYB2QrvbF75
RsJGp15od6IQwJercbdks6wLMx38lnlC8gNyuuUfEP82fP5iGmBOexFufs5Q2hcrjR3Jki9hV1M3
roSAhqOAkV36501FwSUna34JmA9eJuP5mJeynBh07BliwcvS1YTj8KvhUMvXfV8xQ461cTKjcswY
P5LnCROXCjfL/Vejy05mIQVjAX+sYgAnA7XRl446zHRZ8fLCiHOkcjSZAb0nTsuR9H/ExZRsg8/b
gcgep9yQzQqOcwYS4SZmjwdTXAePxeSh4HpCc9g+D/y/MAgn8gaeKw+00yRR3gyuKvHkPmZj/dvY
hlAZjDF5PfrvkcKGBOrfoyb95SQ7iWKQQQAd/CaDiSJ67edMe4O9nLbkHOEji3rJh1kzYGncQ8lH
3eQQ0v4gak51RJ5wpprKESD0W1OPS/kUYPYcLxDqStyQE3FXaOKTN0c7XKuAB6Kp8dyan5VvQd+a
dv+O40hmN21BdcRhEaACzXkpgALD9lpjghRF+yAQD2d2Z5WGVO+M+gbqirzpQNGBMR+gxWwbE7wD
Wl1MJ3uqQ+jHu+eSZEJdJ2TWx/xCCtdebyNvCm0qJoyozYQGdIzlkxRqZZQ3ZwLM4eSEMFOZDuDJ
iR8DL0YXDH0NXOlBl8R31JIujhCmkFGz65D0xzEfl4ckjvGhL7pGvwSWOADLXC6/0ewqiadhbjdN
TFu7egXSqb8tKleLONMvjrtVoKfjsTabf3LjMYpAXQ0/iJwcSRRefLjvRHWzb+Tothj2OITwsX79
FY+4tVHu0uIiAiqH/9B44XuovMnEfUO33pQZGQ4fW/j84//Vv+NWBYsFSmC/ZTIcddt1s+45l2Mu
trrEaRvADhNADpwOZfqiJ5QKuHgouGaVD3nyLlZMFMgP4i+xJMQ8VdkYrvMOGVkYDQrUEvRjRx+T
VrtZ2KPqinqIOV9sHBgK5tGs2u3qKIAUfvo3TxHIMBriFPMLrLNaH1sCzMUTPQAnXHIKge9uwK7e
cVOovQkE6cpRyy4WBCGE85sSIjlYY0165NNdAorR7kn7uzP5I77/kU8N7F41I9D6CWpF2zKU3+pw
eb/d8nh3Ha2NcfP20YJxAIZR1eitAztIFEK6DkVWOqUGVLhD+uYF4T3OjJ+T1NEytGO/GxhfGBhC
4fE0xoZQVtjmlSBhdppL0bCFBJ8m8fbGzVaQZGRH+VnQwvT3v2kVX8Vb34iWZtJWD4TK65nybbut
3SsnN0xSfLO08OiW1utCYadPeBQgdMKKET5FDrsvvl9OfNfenQtAPk74HQJYgXK6mVQBDtSBsZNk
kVOekwYxx2PdUT+/ey6997J7YXZA18+JPUTLRvG3MWYGS5+NN2chCIBqapdtQFnXaxsQ/S1MFzv3
2EOpCa27KtSOXN2U64w4v7993w0q+Mm2ZDm9Xp3Q4XmKQwUfT9OFYMV9d76kQqERTTwKa5HJ+nl2
uo3Xo2DXAWi8DvWCY2c1XmE+tPRsC9xabHFQUeRM8lYgZIaXO4O4bsfvSUqVIqA3iVAvkOFRXeSz
bYZVfBm0iTMe3X3mUpIvSY6GPDwspLlpG3QpVChpkiA2pXMMdtaSbGxLFSCyrus0VnkJTI0fhkHh
i0s0jHuaOb6aFo/feg72nyUo+FsXqNCTLa7SSeYno5i/Ti5hGe+deG2nbYqo1wS8AUybE6nHmd4Y
i4jirvGBB/S5BXivZZsuPYJFWmJ3Z0M7dPeydLE9qJkQ5OLtHkqkoQw4uxjTCfJqIzdbgIdRfTuu
7fh4+ExCqGeNIwF9NZYgI2FJQNIiYVnlo4yqXFYqHprDfgY1r7NeWd/7Lewgllh30qZXwnNNB1fC
SYi35itQSwDDCueDkBZaX3xyYGLJeK6/f/DRRPE2rtswdHqw+Zl7MYxhi0nuSjlJ81Rc2MHEDyzQ
nLbFwY2+wO1bWoRWGfU0uiPgRHyPRpHkQi43EtGIUB56Ohc1PldXvrAM+fFtqUaZ2GFXWSA4usmI
gtIeCeHazFnIkz8WyCE4Jtu/Jx8RuOTzTxdbhTe40/+JS4XtEiBwS5WNNU9J2yIU0E6D01YHoo65
Zrd3R2OumMxfOVmUfmEH9IR7O8McbnPxzv9xs0FjCl28KlxZbsweL6do3sgFwP9JfyYFJbIl6w1h
pHcwAI6PrT4kUTQ7JpB2ijaFeAIQJ8DDPePh5Sk4xReSMaQ3N0NJ4+XyJTTg8Gf9uHMmEwQ/9x6A
rgatIv01Ig69ROjLapn/KIDE0gVJI7YxsQ+ZfSIPJCjPM6OUQJy58cduf5BpamKb/tFUMLd30yTl
3A8SSmdys2jxoddWH3+500GXkMWH/XjIn7cw7D474DGbAHLsdWkwEYkmAdamMaqZN5fh4wBXN59J
CrQUn6ebM31hNBvF2ZGOVOE4bCHClcGdZHOXQ7YSjpERq+qDg74WmAMhLkZKxwvVMQx0Tnn9Q389
jdDU9gGoYMho9Oc7RLKzmMbEkiLM6nkxV1L0Kvq2U0MF7JfC0fm250qg2+Rhoj54GWtLgcGdPANo
8lLk7R6X2PfMn+GdmW8FZRNAnGc6MZAUwbIbr5gusPFkGh1eBaA5O0klzk6cA2EORt2q7DWh9E3l
3P+FvTGFkCzYbscXsZ60u6rJujqAEOwjU2+FJkQ8i6UMpuatMnpAQUB4+QUzxeVn+84yWpBpFpcJ
Oco+hOG/xNFGgCSPxTVSu9BRgZV2f8Zcmvpj/foCnqydRD/zmfEGG1sJcL7FEr3J3d0sdy+0qOmx
ppsnjV2GCbYRBJIwtEgSdB2AKwGAXO17aHrcGfYEIA16V3RX1QlYksrkkcpoE+jxo9hZSBnK7hcv
9Q0uSaJ9AJGBVriwyNab7DxBuiwL+wJ5v2otAhlnFAgtQkNczdBK0zLedPFi3TJAPmCDLQyKblEs
HWIrwTMhWqxC8cD4k7UQwZs7uHySzo41MNxv7E9AOO5Y1+BjSF/X/08wJQ467LCbSr/XNgRKB/wo
9lWxiEKnNQXGrzfPNA3tWeRMEl711jWsY0aF5oEokppNXmQsUjWzAzcCMQCdlA7zka/A7qIQgMfa
LrWKzNPQ5FALzYUlq1rzK013DeKNUe3fGRpdldTr0T5Y7OfXIlvi8DQCfCH6PExKoKox723qFMcD
0nj9pIh2fv4kikd4rZY7ahRGedn+djXvuPKqXzub2K5vZgkWVS1pyl4QmkqJvGggabDJY7w0P9Yp
DZEHlYw/027cHFiCmBNApt2J5xGmcZXfDWDt9cEwT3rGFmALKZahti+u/g0za/NpR4E7sxTe/EGe
aCCQ+fXNFyyd3RACH7pmalS2mIqXMy+lotH0nKgX5V3HkMtWUp0rmNIaJWiALH35VpJd0UddkFC/
7fvf4HAp6xPfvCiYJcseyYe+oWDiPe5PSWwThhV3+x1Ohm25zL64jpTOuEV8M2MBhzXhAt9NB/Ge
JtC2PzUhYUF+EcBcDuo3zWmWnFbw7Ht3lImFpTLzVSgB4TVDnxV0F/Q3rRrcUWP3MEmf/kln6w/h
AXZ/JbtbRHP7Wyc3QR3uCjgVB98WN5H/ByBE922MM3MfVSjDOO1zZBjBy4Cx+neaEzWhe3SfYNhp
HSDHLVGjWRgcnfkDc6okkllpV4Om6YbjFOlJeS3wqW4L6vDrnx/Q3VafkyumW29XZRK7V0dxlnYB
TEq1iXtti2U/JTMYeaXfNXohbgD+8QeX/OGfQD2ldPGWF2qkOMBJYd0EIAdCtKCoC/dV0wpPC6kv
szksi3fwSBE/zo9Qx2cOLaKnJKw0tIu00+a/aaSrcSeCTvkjiNuhigTCrFEF91wwDgNruPYi3AAA
2aC6cFKUu6NsBuU424cfFV0Trmd85AtAXipfdnJVstScPrP5JZ9x9sOe4/v2Swrln/rTdhGoTGrd
dUUwEjNQoLZ2FpiskVZsrzSklRKkUnRAVuNlZwF/0c4kS2gIcqtOPIL1zLt2xu7dcKAU5sdz05fG
v3CtgNhEvf+C5zEpFwsln8Pm4ngh92yqNxDFOlFuVQxEbU7RjSC+xJoe+Ay7T5JG160CvHco6eYR
NVIs5HaoFqYTmSDy+gtfgeuwzR+gLP1B7zY1ltltXx6N/nqfZZN+f3are3vg56fKlKPLP13n/GjP
rV2fTq2uuZKHRbSRNTnfA1fHx+QEfFCVqlAFEJWAM3hwK7x2j4qlnel5KK/vhY4UsdlPYqqoZ6an
qPUvGaUhVrtQJjYZFek+g3mfUpRl9Lk+Bb6fR4NfdG0CP8Qx/Ou6+gUWTo9vV5cpOSaDSGL66FxV
kaL/bMcrAXK6f6RAlomQu3RabZdvpGLlVWUwzXvQ14j/AyPw5Uu4FvW+yod+DTy10WDTQEMr7L2Q
Ql+IFRKDzoaBnXE89fe/BzneWE5+hpsxkoyko4wt/WcXD38lRoDUXXkrFGaIjicDK3kEqQpnW+xR
CniXqOznHv1OxyvEFQuNT0eP5rb0Qbq2AnGdEXWdT62yhT20vCEUS3MjvlIH2wyfx/haSZgDOfgX
7SZDajMkzUuTJQGUZ5skoJL0nEeqXQE49CGynDUkmaM01SYtJWlRQCDkxtUHsNm0EZVvwLwbJTAm
ufm8FQYXoU5cX989LBG23MJrVdMXfh/4saOIvtT14HEWNQptCkYTPlIgNY0Y28xZJGUOAIcnBA0I
hBXFktbYf4UgqxihNVhCCdbxyOafFOM41cgeCieY6wlgU2gkJ1ZZlDXnvW1F4zGy7SDna/lOSQY6
ADby9lYy0S02WhP/kqKTuQK6N/ZPcRp2P1Z3PFDkndPktZZf4dECv8QhIZ+4WpDF0KKaMUP4uV4E
Bv33CrRgdG33kMJ5lfWYt3JGZxHJfHcJmpl0l8KKRNIZka2bhJFf3DBoQWTABg5Vusw2RC/4qopX
ougPraMeIuPHW59S/2hqKeAjiRu9GrTiLeOKHCJdeMHn5LdJayfQOWYqXM1rElGtJZBuHNgbYsB+
6blpnd5YXE2pSCysS9lUQFWpuwKJV/i3qSYkTMcbKMmZrwiEiQF7IahwZVcI+WUib10c0AAToxlC
M1kTMjSHn87T+gUwcPSmjKB55BXiQc/t7e91EfZQf7CjHCJxE3X0z64AQoxkSfQ59Yj07hQtjW71
1tA2+9Ox9uCELarcTIpIk/rzCL/e/J+vOGjUuCYSZ8KxF6Pi6iCgnqHKBFABveKS8REdHdVgAJEq
wSRqn3lRhwW8i5FR1pKj6qS51BQjQwuKuGJeyifjB0FjRzq+SlXU5frNWSbfXqUWrhx1Ez8HbL79
xEhUENMOCIQq9WrGxdcM/wddu7IVLUd6LMkQeEKMxvxFREIKr7f0ZtHy4bzmVlFQMjDJKK95pB8k
ac+9Ba3busnuCTC/k/H5c26OWrkEpbOUAJ6NW5g3jBPp/WqWCgdTeONozjnErY+f+g5T960WgiUX
2NThezwH/wCmvAVIkegMFaStRvPNi3y5IQ76CTVuhkmyaryQiyqmF0FAmVre7YG1YVKCx34lBjed
Hu+hRYsrSbPsbeUHxKj5rE49DBIEQprv9JZxBg8RwHXArAMqrV1TOnhyeAgVxYay145UcSPLy9CL
uCtZDR+jMBGRlHFLQMAwF4nrbnHSItX1XXz6Ie+SL96Zc7pXOaAFAxd3H0dl/feRqnPaegizoiA8
FnjzAunRrMYCHMd8hWTtYksYXbZg0W6eTNXuTUuuuv8nc0t+A22FU/AII+sg8cTU4nlhzx9SRjxG
IjAt0L7bbt8e8WgbyanZLPtOeuqToAt0fDyXvR0tMtCxuJPqMyQuq3Q/DyXM+T76GmZYzWYhfcdX
+u76FTM1wgMZSmQsW35OZ7Oplj/vYsGrmD83GtglVsCCLguOVE8eX/0V0RyTbLiwAuYM+JkptKyM
yieedO/M/vYbzTboqR9qVoIzUbj3mzE057ricX1rhwXnHd2g9xST3jzZzIQEKDYLlp2Kobckkmad
PeJst6iKAell6WNMxXT+DqIaeClhDVhcgdoDnQ6iRw+hwBrkGjN2LFH/D9S3FzWAIl3ZWj84oK0r
GArDrF3Aan7v0VkSxfSf1TpaRMq/AuGFCIY/S829t0MnveZQHcOxsEf3in14Kt/MLrXoy2F7eHUz
vNWoh68DhbppN2ZIrEx9K2OBRrsmhLYsoQcfpstoy8yI5mABEZGZy/tn1j8cb+0zBa9wIa6NZH2p
x4i/2I9B3oCH5pzbez3fAxNlGLuq0xunqkqxGHTyqoRM/2itIuElhK9zaLrXKWV/ZEVUK7al4u8u
sin31ENwlU2pxJOG1aUVucHMKVruFCtjN9t+14IkLklx01nvjqSQtb8SGdGGlAranm7fQyJCx/Ry
FYWoQ7Vc2lziCBR2RQDc+0fFskpaK9Pp0Y6Kmxkkw0emiYN1HptcdQEkCScHxcVXyb2UY5nIsobP
Iad0xMTpXww38CoVBdMMk53mDnMuVce1R3fZOILoDuY7t4IbxF/yI93eq7gXOtzP9zNqeqPlwOtD
c59BVKdKYAUQOOcecwQNGHlGdrIrK5aSj1MEJHgdRsnyQBM6zTRtzLlX0WpnTVihR0KCtVt3eUFW
YfXmV3i0ZRJznF5LV3Gw/TWjbiz5JW41SszHBB1wniSVIzLj2FQkenRwwaQuv3oo0rJm4FR0VOjE
Om0BQsDP4qm2+6VP2gR1jdsvfYv6YpfN+N/aFYFZb/HwRNhX28fR6OK6s5MkcMtE0DZLy89hGAm6
7ycb9HcXDaORrsd1Pdoag6Mc/0UmHtj65JkyWOO4Jc3FFsRCoDHJMCW0TW7SVrP/NIVE9G8l+i1O
LLa0T2q81NhMUG1pDBKIqeD6mbGqTaJkgd3xe4+dHBKALTVj4+TT9sAC2VdGPXSFP3pfobpl43yu
GJDc4rZiPE7bma/vFuRcZ47FO9NAj3FkX6YbLsn+pJtGsCY/uWWAeZ1OYKHYrUqiWX/tsYwtzmOj
ANkLyJgSvhn885VQNxRZf8uuOfj0kEjEI7QcRtwyFZx9fNFUuNmpRmUbUuHfb5aok4cu7SYvac6I
s5Kj8zsl5NTMlOG3xdHKpLvTfhdcT40Bp0QlnU/kPWIASkVFET0Bm92kzl06f+DkP5N7wHvct3qS
hZAxME6PQWwRgcvd5F8Njol6ihKXvShweO9M0PVB3WZIv3MJIMIKJSt6bFA02ZIjYXfP3k0al8rX
IxtErh7tcuHpW1yPdZBnAJuWTlB5BjJykg3slyNpCKTZFmobJmSWEsl9vyyZFOGNieB5F658tHfP
rKzcjTHKWAZxrorJDMqDZNKhaX4sqHWfSLmEVF5QMdGgFEgdcGBIbP5g4x65xp/0gFN5OCFjbd0Q
IInLa79O1zwIgL7nX/lDzqcYfQu3NedS0YZ5cDlEHPZyunmclYAS/wUmBV7xUeXixBm0iTCxV1I1
CM3UE0CS/Hp/dLVcQj3Lt85qIfnd4OEN3lCb/FUOyPYIF6GqO6y6wYOae/f/vml4G/SMJCoFaGWC
Pxj0/txpzif9nwCmQkmQOkGOYy4OYyv8Y6lQkRK3JF7p+mSM5XuVcdkgZuvSvkpLPUylvtLD2kpw
wf/uQmtYslqv8jhLulx97lSokO07UGVsok0/fO7rRLZe8WR/36uhrs4Y4vvN+YKwcYIuOpgz1V6H
ZwgtXkajzwv6pp7/yhZcyva5tSAqonWdxwECk7D/kRuBq5+HOgYTaKg+CW8e5kDlTrcAThKimWQv
18rftPEM8oyWNVI/9+183k4byVSgdeKtukNgVo1hnnVJCa6Jg5Z0ASAapZWZI8NK8UKBpuA6pTTX
LdmxoU5Fde8yZaYDlEITL22Y+mOcyW3V+yNJpr1BHWN6yak5tL5wjGa3/U1Z+5PyHQbO4LHSwS37
+lz4zy65rNC0ZuDJdYKv7SelmNf1qXtPuRQRyLa6Ck/12BSrYdsl+f4FAJdXTKCgpkSnaDBlznhf
VwYp1DbFFYHHDQOSHjZYm+d9Xie3wyfYHCfEiOjPid/akXf7MNjD0kAoYBBkPYAiuqVIY+U7IgW1
UiZRcONSZ9BmwsoBh2PTkY02Go9E3koY701aq7yIpMf6DhfGnXm5LSByKWwQqangZ5XGhVGVYXom
F/Q3x8c3gPDsYET5ZvHsKlAREYxbRZGLQQ1kq38iQoULX5Tb/+iJCet/6yqfQdGFDooq/O5f6Y5R
ivd7OoVPrmeXJJtMNvG47A9wdjo6U96rEClTSxAg2Sx7hek4nEgYLCczpTiyPkrDVucnyGEzHpyK
lyTTlLLjlA3JOKr1Srkx6iN+7oFwgBPiy8CK6z9Y1TBjJ0zF9t7dFvHBH5kRV66moSyeR5iOMhsw
mT8bhfMO2dsgCB/Nc86Du1HOrRHUIndldzlpOLAvtZ3xYPqNYGa6xN1O72OqL+KqD0hKmjYmL2nN
aOp/7iIs5runcr9cTchgDtvX0q9zXsla1mX1FzrA+mTybLoPUX8xuILC9lK9VkqjUlsFpNRpdSUs
uQkZrzfEluX/4j+1nCHVWgyNn4yklkAI07wJtdR0ixl9Yptt7zHLJIrSpgQqgUFKzoxny6iBfEgF
JIVfsab4ULzyY+zwgmtEmxoSX5thIpcVDq5f13gSYlGf4cZzSF3U0YYEt7vjDgWKA6vQwMGh31/w
p01q5My5z8fq/55xuTGxoRG2Lza/ekz5hXfT9gfSk/vAURkhID7NoDkOYoOTT4iLnD9PIKNqmd6T
kBQW1gFr3sBNbQFQLg8dnmL23k2WfG1qXPioG6Vb8Sr+ckHYJIRGC4Lbz9wLwtG89wqv49ETewis
3oUsSdnGE+5+X+CkijM1X/rt01nPxYAeAxPRHQIVSFxBr6Inwe3EqwtRVtEy/vbGuveNrcjnl6w3
yoUZoVLVYE61t1ShdWl+OymL7edOKOB/J2XnHJgUquXrTDepAS+HloHNwJlvRDXXJtDM+wwZFlTw
CPj58ev2l15aLdSQpdl+Clb2cRpm6cbcmoom/IbyaU1ciqvil0Gnvk2BkuYIhEzP6opO0oAOfUoG
e34nfV6mS1z2N1dZIjWgUcmyEedYWcR3adzK4a+9NwHN0fkN9DqSe4YICK48DJySS+At23PYeybn
QM5epsY/1IZMLDOmQYdODU0KPPZmH8ALwversFlSqYczWgmJTdlggkvgBX0XhEclvdCCUOEeAG4F
tsTZHIrjJj7ZAOI78WTYWA3M9yIFIf1T41BU0ysSej+1PPMdAdvJlNMCodgV5Wbp6yI1qoETM9u2
a1AbS8D2w7YijDwkBV0DV79rHgFAiIYJSOM9qPjCvD3BEGMQqZcoadwn+OzYybO1G+HRnLraW7Pb
33qzdJzwCShQoRTinpMHiUVucNJvkpECBZEbMRnHzGeJuCuCEGtrOizHFQdgBVBZMkW1Kl1YVdLR
UJHP/EKY2qTRFf89WMv8Hsb9QXC69uCGWxGsndiH+gpiG5HH8j1AJeeekaT9XlAoQKG+embhFVsS
OwEWxNB/n9sa3aj2gqZrez1rwgE9V6hrRWC+owGFsLCsKYbAHHjubBwEY9t9bR+06DlTI22Xs/L+
wWYfMomNQaeiJRb5uSgn7ThbxuLWbsvhHXRiKxYKWy21cyXwTxF/+DmLksr+a7rc19atu6bw4Eiu
7EBOMcvnA+M1IZX1uzSCHLYARpWmC1BKuTIZLjAbbUsknKenr+sGdouN9t6hR94uf73osPVPPKvU
chRxpy6conmdLwsphz7ThzKPNyoe77rwpEr+33g+KBgw/TWIhYklcOKHrMiJVXQkNONQZdgWVqaM
Ydom+KI5D6nkq/f2jg93tNPEFOS6mx1XHNieIaywsSI25eazXKKf8sRjjgadmbOju3FoN5fbvgQQ
m6gGCRo/FQXGiDiPtL8StrcO4ishfHY5Xe4RVmb+4hxn8Hli+cRI1dxqiiR/qEWQsMMt745vhjFo
Dt0v7u0xJ9CChGygRUzzgZw/yP5jxSJXaltYcDfBg+xeEr8uHztOqX241RqDSDrDqONiJo7IwBvA
38l5rgO4ANiwF3eA/YsyQFiojCi0MKXN2l9wSMnkU+rFgeEpkDRk5zpxnUa8km3WzGbMZbGk1mWz
qfrzIYOOIENcWPvjUmeptx4bcx8faZ1hUPQU85ZfM1itLrUw9yjEJOWyYKJsEWVkAiG0/jAPMyaI
7lw9hI/I/sXra26mvE1NcCzIaCS0/+1iU8d9jqph7bMhtO7bACjmlE6BQdNrvLnLNWCyTKeXBHP4
ZbP5AeYCfO+46fvAud74UW4fPnv+Up2Tm1/Ex/tZ0+nB+FhYiCsr8AG+Q0myx8F8FjiCLcGn0i/Z
XeFyDmj0F+QczDG7G2tkcPLI1s5EvaQJ/NBs2LIdh9Nq7uJictjxye0kRe8byEQquOQTOGZH+In3
TjHPENW4RfRDEA9xFzTEAuZJkuJ8irz6yKg7mknYjr0r5/C32npKEIROMb1ugUmhKECVWK3w5K+y
GuA5zc5dJ9WttPA41kjeM9fcaw+gE008WHveUHLU4T3x7Om8tA47ATileap17Y/2oV8J2UleoEyg
RCjIrWGKDBnNy+joi9q0a6DLAQGqvHJdZS+YF3Cua7+cAwtoXcpeDSde8znzhmvOjPaE9Dng2KlX
TFc7TzFKOo5bRpAxraJZoWP6cKiTuOQYcIxNWX5P5kuB28sguAC2VVr4XAmQCAF+KRmqZ5AMI+/t
ndT/hslKZ0/0sLNyzYhpNnqU/GmysuxGwT/ROiup8MbZamgiGFQMfUEg5sM5/0pX/cFUaixOPBB9
D1zVde8btDQK4CdVvoGHmm4yX7sRSiJpWcYH0HibZl5CCnPjIF7a4B52n6nC/BNlt4Y6UGWPvhrg
kgqquzupQ1WHcom7BZfviHxMZoPN04CAEbaoBtyv34zgxkZYWyuQ70POKvufeSLCCnwXvw1DY87i
totbQoSyNrp4Ffue/HnjlO479I/Ok9q4xLOjcmKliIinUQDcqXlWTwi4eJQFnGX0df0KFA+ENouR
76+0lylYEMmR1FHdiAiTbyNlcTn+zEwOS/4XLmuBpmRdIe/Q0EztxX05suUVDYmcVCd0szJBrqWa
KLjpSalyfQ6U9stPRjqundnyRJ1bur+blxxLggUQarqHBd+zFm/Xf4okHP3w/t16/+uk5cmRhPpp
kQq4AhGG4RGbNFaylgxtuW+p5wg02Ob8WAI0ufPNxDtDUnf1i20swGaXh0n0FgI+aOi7YgtQCL4S
OyBdSMDMJwtXvEey8WDw22uVBY94c2Ik0vf1/mwmnXga0BkkDxir2pkkTtCooAJR65WEYrU3o4GN
RsxjXPN+01rGtQzUzh9J+j1MmR9xaTi3AyfOLOP0hERbgKKHwbz+/5PyzmRHQpfK23Ji/l5Esav7
L/8mhD54DRjifnzSn4i81uSEhOAT5mm5yRxVLu8zCE7KOcwckq8NltangLZnN8tdEXiM74OwPG7c
7JozRudeGej26ioqHCo5VilWUNxiQgjY9prHAENo1hsLT1U1/V/uA/5m4jjdkTPwmw3CM6dDNCP0
5o7+bLSMVqkorQEr/1HeOF6bF59caJcbn/xUo0Y0F2MApzBy4BWmbQTuQrDxhsyP/ulM0i4Bl07s
GtRKAMeIoCNGT0lpFo0fSociXFqlJHdSJOWS2FhVVwUhU/EcBt4ormkpzyVj3T++Dy0zppjohZ3A
p3vjLX1AApgGjDPi3lQkamOETSoEH35x2rdVlJIB9dm9iUcZkW42PE36NU9ac4GEvxqZTkgmiqs9
V8iJzRm7DGpc7MXcTEkqjss9WJZwwkO97b+B0rLKDIRrsnNEeO/s2kcuoNSgtnK/s0DJSPziCllV
p9203g2ReX35D42zo0iAF59PJPtAByAoudIuegcMmzvMaRnX24t9S6JZ1R9XfsKR98Op91waWm3f
xyCNNsD4N9OUBq8yCInttt4NCsHoTgFDkKpUDMJAoiVtOskcUaJ4MU9itjuG8P10KVs697s4ZxBO
Al8ernIbYcle2IKo+VhgttZxhaA5e1KB8+8QO0f4WygDKNMZBaGCgAgSlf5xJpPLRDYPE6Rn95Jx
nePQVqiBLdUqk0b/th2LAVI/37dAgctjX+5kBcT7y5TQaniwIo9KNwaIFl3SG6JyFEqVvjn9mLsv
fYuDesKcqTxSOw+kBve/DgI0PXXz0vVdvw4aVIC6FkuFTH/GT/bCDUHobLpvKAX6qChPtQkTd6B8
L2fLxwSJXiS0DW3UbECsnnPBsMC8QNI46/qD9GrJZMi6MnrjeRRuokSIHQh5QenGpRZsxYg3OCUC
Sw8meXX/B2BVTIm68vC/JQ4wq9V+6AloS8WAeXApFsAFK1C8jP1NLQxkKVNruCZzyD6Izek5tLx5
AnDX0U/WIzh7UU0jtom//sTnQ2whzi5pul8qnhbVdHGm3OGO1ibK4ZgRry0z+XcIjT/WE8yhDvGe
v7vgtEnWYB6mPhTtfrey/CtLc/RAnSZFtIiIajKa0xsMR0whCEWAjWZrpKeKjl2cj+wNFGjnCYxe
hLhzDKqedOmTSieagE3V0BJPRvtDM9Bai2rQsW68MUl+YBgjyA2wLNxhTEkRGadfEn3bjX08DYxH
za9vO09AysTCuvJYWWLc+TQIH40Yq0WThTS/ume4vGT2a5haIWu1HGYYiORdLdXf+jKBPNdRcVRG
RGwKvaCHiWocpj5eHVjsKu8BeFcNUFUbV8cUvRNAGLbOG6F8BENLTDklQwYiO3MzkPPsG8EajIsy
kNAU8UKIxbNe1HPOA4xyTi5n/74MpV4cdRYtDjjjvb9a3+yRXCTTU070pAFcX2ujkMGaqhdMrYA5
6kHYy5CQTYOaSoLhbX0oG9P9v3xWtrc3VuG1k0kBOG5H+Xn22Emv70xxGbuVc8sHoeNWoruQVwxc
oMbwiREZBRP6Svs62Sxauso4UovUpkrUe3bgSgbXzt3Ny+tcCJafWrCxtiXK0vY5TA6LPo9hjLuL
te8otSIp1OcIHMtcO5d8vz58mkpy0fK2NvP9zujYl7b5V4jAy/a08X0DNSuaeRC46DCXHKLJD1yP
vyfu1P2pcVfvMe/l16wTncS1PL45eRHGXndUyGjfa6rV1/X6EKsDYl6sJRaGpah+UW1xO91Oay/k
tEXuCgVybkR+GHCqNZpI82kKl3b1La37xBuK75RHga3rLTCk6aZzSMcUsLm97oP3IM4oFru70Oxe
WkljB725dCOJyGZz7xjalxApbFQ74qUGJzfxuI8yo+Z4KXyuMzNi9arUQ8R8D6zoE8GTmYa/fLxe
G69qQP3oW1VsSHldO5+/VRZPRytGgVkXL8kHoN6em7P6eMeY5zlilRxdRDnEWeXUhlfjHqXvEpdJ
22bTTeeqQCIyeykknGFGwVqqUQY7uLF7Gn1dcIke+vfJMbryqU3vHKIckVrEWCjVSfeQ1KelcAih
Jy7sEXpf2H3B+/DdFrZXO40FUtkQ5yxXLgPwfehi3TWRT7mKcoj63ES0ur9aFmPg2BWNIzQZxbBR
Jku+A89ZfXGUwIzZQOQjxa4O0PDzcmlEzPIcQ1Kpu0BnbHacMowRygIFiSmz2+ijzmVyT1ot3Owz
vkf3Wju2KsIXBBHq6dadBjWm96rxPFpPcVyIicDS+PBZY/qIYmrGJ6BYCsMKO0vaTxsuwYuO1yCl
6jygpxXe/z0d27BP0y6WEvso2NXiu6zz3eDipXIxEqzLinF1RIvu28ilNkt916cpXKHhmCOYJQKi
sZ08Z+wzqATGST5Ojg0n57qfg4uHRDm2kzUAC8HKxGhjxYmRxoHWRBxpUOWOwh0u/IsrCl2ptP/I
8Ff36ksAfirCmmf/GjzScfMPJ2lddGwcEJDTl4wNLsD8PPPezNJOmeqWQVn6mOBrwI3bfKyEqoVK
O1P9f06gBk5d5xoMVVvTckOsoEFC1NY9ILtRZL0Jhn4JOugoOABw5rqyVsai3i8kbTVqdnPx+pnu
WbYS5s/xKMiXuY407lUGkFugnbTdM8hjWkKIDGUBZYU4FbCrjQM8I+IKsQNtIX9dQRuJaVslpdMV
/CMTKnNPwEvg6u8bww3gt7C/j9/tuutVvLAmN3CK+tQ7Dsy4a9Z1B9U5ZikKIPuGqqV861P70a92
33cuHQuugT12677ngTiVvqjEAeU4/0dJrM/baLoBTrDZDSNFMdcGg9SqOpAaMBXmpDkJ4PQACUhB
nOuzIkqPQ0JHMBBPh/RpvSp22f9TX/KEMrixBU6aVRM+H7JucExJkndLo/YlLIe7Fb/6sVDfIW2m
9eQvwHnEKMKHDanne4evhr8bT7/v1Wt2NI9KKg5fD+9AsGIFws5AMOfA60AhUaUwZ2NEKRZt7PLw
wJY8L42E/AKXXXe+3XOyIUcLP8yWKuy4TkVr1B2Y/azNujmbFJktLqJPYe1jhpyJ3h7GVeNV3pKg
wxChssn4AHFdcK+J6Euol5UhZhGlRL8FSTvt0oucBLgjrpPJ3+w/iLAswsRE+Zjx+fho1IeUcYUs
tSubD9TV/sex96XhtAenq9AFiMXSwjuk0WVwy8nMknaXraSBmqWCbfxWrtgZYkAEC8fwMk9VPhmG
/rg9mbRXIJVRl+33KGwetm6gc0LNqP47Y4OpOzGqesJ/F4b6Y6Rp4L8QVH5OG4Rl4l3hnpOeW65M
3PT3vUbCSN176BJeMZlvp7VikqZUrvqUm4SsbVfo6VHbfysghJLHCI0wEFN1fs8Zr60GGYYOy+hT
pqamw4Nhp66Uw4XqoqkFf3ShA64bIs8lzW2Q0Q/LcscvW5GF3ZIGNBibhFziBLg1qLOGwQGL2SbG
MePgXbHCe6cfIXuomQ4r6H1UQN3krnOefurAGgoStsG5HncDS6GCoI639avGhK/q7M+xcbW0NQMe
gRYmN1MavSGTRY4OEIJu0k66v1Yrl3uFakDWa5kOYgt4xa6VBEC40xQclPHOQSl+sQq6nlR4DsLF
lg+ySMyU+qMe9aAv2wxMVrvn+L8+/TgD3EhyiEXMnu80wzSSWhidsgxy/BuWFmR3CsKfjzptiBw7
PBpJ/RYHx63FcvoaZlG0HCDBzrRU28X5bGlQcTTtfrIVMMMzcipsbPBEy+ItCmUtWPOcKNA1RskT
we9LkWufNwlRYt8VHQ1F1xnemugRU8yW5gt+jqXtzSFtmsUGfq6COwRKzaZoH1/5ZoIEESZ9siFI
+1J0IocfIG3Dz21y59uJnIYf1EBHKLSZ9CFyXAggoM6bYXFOfEeh/j/01dDKLzy+qoqdoOqiO4No
JPGsviV92DXx4YLd5dY+23UdPX5RYtgQKrgkoUlqEl2k7ZEnj8gFeBQaElUpWbKCmh0HmyEFlsZI
/o6m8dATn90332LEh/67DiL33Aloc3VaHBmp0Xq12ZlMB2n2+TxFM2zGuyleYV0ff112EHVS4Ekv
kKchgDJUVgy1agJgYf9U1k5oXI+wR1t8BeJRIWb6g0IiEm0XQBQulTwaQUzTiVQ4cVkqv5qHU64N
nbajmG1+f5jNlgEpDyr4+ZdV1hMedWNjIH+4T/fOl62eIErn5WmFGISKxLMI3wrRuTj+nhE39ANJ
ED0cCgaIHX2+g7xvuoX97cQ0ax97zQ3k+hID0ZUcjhA3lMP33qd/KvjJbk5L2BceIQIvTZObRTwh
xGRwkWlquMmfmY5aDLk1blgAR9V6zLUsP1+V/a44A4UP+WNXpzG+L3QQ92qJZOVDb+p3qO4welXL
rG1nTy3ZDU/Nle7LIJaupA04RfTTp9MSZGWMSnELlH/xx03mpv74MruvZjWdZgqglUdJMUwzLVAi
zrZJ6xF8r0pocmpEMEk4zkBfAzdBLkKkboZmqLOMnwhXRgLnbGjIzTPII/AN9hKzkT70fhZwr7K4
2kCWiB5hnIbC33TN0grQwE43asN2PJc68t7/8EoWuqc/sIEIx7h9MmZGobbLl7GLCqaIZ4Ck2v79
OQGyiOVQFGSfDn7OnvcbF8tBXD8aGw05hcX0CFOy4qLt6o1/aLOsOVvGcVDk+6sQWmwz2uOzQBaI
F0DkV6j8yNkHOWBpQcHePLmfv75wqibJmFupPcPTwgFDG/jiUqg/HsQb4/ivI3zo/LiIRjydWiSd
yiH7DkW/HL0cciAVh6+j1w4hBAHhvi451wbTMOIXK4eX/KsOty9nQkHBsHAIoxdI1opTS173ZfgY
CyjTGjHInsKDF41FQDysTIqjpZ7TrtcdOMyr1rPLI9lCkocALvx+R+/d14iCK4Xg7TUJisCC+68a
4CXl1NhQfVh7c4pFe2pNHGg98k32bfvZ80XuqgBNE8e1AlV1m1ziOjvJgEr10LaUueULoJw6rO4x
OqouhQMzbezFLs07Bn0mGaRyIUhBfuqmINxoYvjndQmwRxdorcvZ0cY4+Tal62vLD5bw/aw5J9yg
pI/duv5w9y5bEgS/FpJMFKc0PMdZxltMIkw7l0qXKTj13RqtPS0t72z76itcvTaHzxrM4IcDQNu8
dOxNsErbEzcyC/JG5dmIrb4HgFVf9sTaIVNPDBmQaqESJKcDPR39om5k47Q/6b3uN7qwsrpaZE63
yHlGz3NAgGoNgLLTFv67Cq+elBlHk2ET9c7D1imMpSgtm78Of25Kp9dWrvRXaAy9KtW3ZvhzT07k
YvkxgX/lbw1Z/ksG8/dhmSw8Q5G+Q4GYBJIZljB5HxZ6kB0O8mIu7l4KVKX85r8ezP4tzicnjjGJ
Qg74x820veu/Vg2F3IixoAZ4Fz3dQX4EGMCdrt4bR9A8rcoVX4pXm6IFob/xv9nuzoHycxjspIVn
mGRmcTjfw5ultIGPDN7PJv5oGc1Y2SdBnojk0T0AMZKP5AqG6W8lCxs8DTZxaY+egAmG2YzoIJ5z
BmzhpoKzhzKqOFb5j5qYovPYFZkDsRaYvWTl0L3VpcMVc9eqOthudLDw649e8AqsygiCmUWoRgTt
itV1qnhRSOVdfK15Wx3b5rRw/zgWH/YphbNp9uoilff5R/xncdnOv1/M8w+9bZB2njqLFZx0jJqy
dvv0lx3QTAYCWWNMaJiME0mXz1MsMmkbwL8JKGpSxyn3l48VfM8aQRFkRHcLACnaf5AkQC/SDmlk
Hu2HJVUUHs4OGlVPm6aTmOpThAoqgB8T9D96x0r7KHUoypJgMO/etQSyjkMIs4AnIRL/OAh5VkA/
QTz4Esrf4pWK/zRFySfP89oUDHl74vX4sdvFq0rDKkk9LjfhpGip/wBdEYTwxfd22VZw7HKZMC6u
5H7X1AdRchzrZ3mbNOcJtNcYfYICDaj0KXCJIX68MSXuvEgQrmvudUTTD4jFlBzQrw/tJaRVfVb2
X0L4O6ztU5kiHmUR/Gdf/pINvV1Qz5jPB7b34qLLWRviGTXwEQ2vQ2sBoRcNsPoNa0KRWK2tiLr5
BUjonXwc2var/irN/vBKwY26Q9VvEg+7aoOARqVBs+ad9Dn1vuGAakNMQ9YWhdpzcnTL5pJkTc2M
AG1eFEF8CIVgC9GvvTZ1PY6b8YDWvriNdEf2u3XwQMFf4IZRbTgE7JPACuCICcXwm/15+WXPr0B4
YajcBRTxUq8AvnE9H1bqXL5elmvBdwvNfLcY/MurO19n2tEkhWLiaXnYS5Y9U210unDLtl2zlvmu
Sd7qKSzY/0J7v9mJP+Y8nq6Dd/HfNVDGUSJ+UBGvvtMIVx8yN4ayqpxMwdNBNSnDk1uDMy3jzfbS
l0o7NUNo6KkdquPsUewDpE6xrO4ismZGe4SLceCQfj0xVhiTc+YRInZ+CGTB1sGRWND90zq+th/k
qyBZD0BB82i/7yaaxWiL85UsDZbZcfU6JVsYRrKz2mjlQ+a4KH3vUFjGQoGr51cTw0NRJeDUDBWz
7/1bu15Hm8flMsufS0uN49eGL6ycTssHbE6QsMLuA1Vla/DPmtB9U+no5637oFN6k9y1BCJABAyD
nHKtBb7zXMJ0SLlEiqXJqxbFm0qF/twLZFack6iYiruwEO/6gFskWdB0JRevAIazGC5eEOUUFked
A527mP33c1Sqnnw/bx2b1qKkHJkB2FTUB3Knf4eEfeltwQ/8CzRALMsBvqsJ9Xil+eUlje2EjhfD
fCufRPnmmthoo/FzxIdDxQgwPkUEe/Oar55Ye1oOxQ8ztYlVr+BfWL9GC1s9VOr4qs7knL6vTy+I
p8ftWmTKf1h7+2Xy+OlQftd8WsMv/Y+vG12UCT+MxTQ85PXMC97Ak2TnSaFmJIwoiLANgARz5akE
5SuGU+Q7vXaD9Tl5Ju/i34QqMAxvU5peAen/UTnwO6X3z2hW7O7ztvKJK4PDOp2Z1TjLezL3IjWg
iYPtQXKn2a5aCzQdqjBV737CnYEBRJAAxArq4XxH1wQAW6YW7Zy02bnX9yo8f++paAq+mh9Kt56S
/zDwlIEkqdsw6LT2EpSbGQL436sNKKzc15FnQaU8glwt9TnJ8oDwGR95lLMnzawqBZNHU3Z+gQ1i
gWVoITBuxJh9K1Uo0uV9TD+t74+AcBBMVA89JI08eU+BU6AJZ0m6C9rjsHLesetoSZrtZDYUckb8
HHF/8yxlm44UGHaJ4H55ZwW9uzzgQMUx4AiJl2roUZY/zKEueVYfs7/W5NvOQ9aImjs3lw2ZyeGM
Yg912fLSIc8hu6V1uF7NtikUCwa5K940KlXGtBNLvf7/UlFyTY/s9lHkuNVKn038QSJwmW0L+CrN
laf5dPtwR06u0OAgiNS5aSv0WeWkxxfUwes+6p5X0FjjL/yen2Tg7CiYggv25pNoIPrDn/9bWgEo
VwqcqHosjtwc44vuNE2H3ksFmq4GXEpr1zMC/7oengP+8SVqzz424V6WlXy1mqBeZLMmjQ9MsiTM
K+ryIKlnn4gdZLnHt5ms7yPjE8rUGUCW0pgT0gkqxxYcB3wvGdE7n5N1UC+DOL8a18sSOS+sw6Je
gKmwtDr50YVl3iOg9/Wcp8pBDew52XSXtliTeGvZqpPyVnS1noFboy4FrG/aSWbNIKZ9LzVGdK5S
AYEdgWE7MHmgqT82B/XvcCh1YhTquULEEP28nrr9FhbZNteIMPoAM03eK7pfb1Qmww4kzWzBkPZg
DwZmCjddZNPuF2ksoKD4L673QXlmecLIvQT2C5s8+dxoS+re8hpy3OwnVOOyzXbTW0C12sLFoQyy
BIPaK2D8UAiTCXxs9bpCujuWdjk3lnEnTs6C7t7xKEI7YSObG0Xw6UM0g1BxTIyUmbn6vC8chEas
IgZcQG5/qG9r2bte1pG21bAUJr0+ybcv7U+i2h1GzoCe6suosnyYrgFMxtGZFbUHglotQ1A0Fl6V
6Cx+eD90FQ9JQMKu8uKlguWxaj/HMgUcr1PiDgSpyl7qNvtIqnCI9aHZF4zdolLgFzHv7JWiRNw5
FY2Ib/X5rAmAedxE8/oFn0FoGANqcfEwOFOKo1nHGlgLDL4fFEjaBWRY78BJmeDvHu9GhuCkdinH
WM+eXmQd3wxKiEtR62wtUtS98eowM/6DL0fYA8sxsVraYw5LgcZE7Elw1snTSjzVRJmZHEhXaJMD
iWDWW462T4OHXEe/ck6S3uRtIBoSzN+UsMzG0SGiGqDhMUNK6bcTZNHD9LOCME1Y9LxYYHnT+iLA
k9J632HX3i6+VpQ/uYxWWE9Uvgrmz26IjhihczXA6yTEpb5+CpiS2kdYuVWrDZrVbr7COvv0oNCU
cQ7zid+7hEO/Dy0bjLhQNwHKefBNaLVxz4i59BkQ6xaXqmEBVJbTKbi4c3eo4NxqS386EiZjKP9j
lmCTRBLYopPYwlazPpqfCtF1hoX1y/tBk6Jsj/vI/zES3Qg/sV4brAurQ+XYhxhA2aXc1pSIcXDp
7KnKG9C4tWiEkWrz3mf4lZI1+nb7eQch5THHwweDBE7XkSY01GSwcxcmEoxPLbf2H9NNa1ku/kiq
8cI+CaU1qYNVrrdhghOidyhrLnfX3MPmlM/DFGvmyOBFIE2RgTq2f1n+KxnkmQPklmEpL3kDu8CS
UH5nGdD3K2fcNAvjQONI34gXOe0Xn09d5JQ9rbIxEY/jJ9PPIn+gwmEUS1cxd16jxGsC33HmoENY
tMbA+PTiUVj3w7Imf6mSRL4wWFScsDavitpcehH8D28yz6oq3+aFc7c/15Mxpf0RLZV4EWoVk4MC
wOCPE2yatd87SuiZeKin8euoqhyBk6wQ+5X5nQ+sislTtoKiQQUrN9Ab7FZDkjTsfS/ejQloIpbL
ZhlcUj7kqgYdM6RimfSuVPxwfOfqIQzQ8LPXGKDFMkdB/4R1nEkV8dfqxbCdIzu/PdVnKrRqUeug
1rSbCGp1EbAoimeZzZGNu2T70yci+b8Dmt477p5ghzNHkllq3HYXubH0eKU036ij1ay1g9Ixf6Ce
2PkYFjms3eKE9wY7ilnFgU3dsNOV4qqPQauI0ZzSP1XSRzlEyGRQZU2wHiZeqxlmVefvtYJi5ou4
N8s01BUwvTeMjC0Pxdw4Ke+wzvK+pyzcvC2vNpzPgJxCdU5dv9yedIZ6cvJAb5K8YoQo3n3oS9ud
tFsPlaT3JBRKGgPS/Fk+VVuWpz53iHfgimtjp7hg8T5IJ7InuQAQHQrWlku7HMSRBNIphJG590cB
ToO79P2io4TRWFTEPGkAJm+PA80DXrsCPZBsUla6CW7XhnzYboKeeRkrewk9Ekuv2zG/xcYd58Ux
zMcMFqyuf1/1k3KRu9azJSTr91HLdozst0J9Fkyjiq42m5ZDLrzAfW4Wk/o3uGRexgpU5wQb6XPa
ErvW3GSpiFlPDqA2xfhzm62VAB/3uF97T4ujd2plsZ+cgFhWuitATeUzc9GMhi09X12d1rZSS97n
5yuBXenDsvDhXlbmanSL//LPfy/+/i/sz3PNbOKXkNeBdcCKNxIZ8woI0MQow7aclryZU0/ifLL2
CGfSKBR52dcI0tTiR5plrR6m6QuCpVW/dh8O8BNoa5zcX/5o4LVsPpn0IdQkHVjrOipolRB+OcwC
xvlhmhho9ZgFil76gFWfcbB7aGS+FQpnE+kiv2u7Aw2hVwkHcFD2jbx3nxkg7hAFoRKaJOvPZwQr
G0Qi+GEuV2hPOP01ssm5C1sEtvp/ts6J9RpnWtxSz/ndP50MYQwhW73jkPX5+Rd1Ttib6+81SLjt
b99L3sDxCu4z43CxnStGBxMRB7BPmNDd0CpiCMErFl8jSrpI2u1l/e8r9AaDcDZDeMxk9bXMelLp
hhC1E00bcdK3ASESu6ibDmHpkHcQ3tG1pKxZL64wS5na1DEb5mV0Mr8GnHlp2fkoA5Qc58DwkAdR
+j14sKZnV7gocFUgyMZ5Xzrcj3Kdy8aqJd4L8DIpc/CzojYV1qEMotqv3uKadPZnOTzEvLvev3m+
98tSRIk7/WgUuaQTswACHBrIeoJVjhKs9dtYl0OZ4q5WumxmokdbCNXHh4Dm+PiDwVaYkpdv6HXK
SQxnMyVz6xMSCx8zhu+oYAuGz5mkGPn0peH6H/wYon3lMff75i2I8cpYmzT/c0wH+2cksf/vOiQi
esfyKTmGBgxpoufgVUkcmiSPSQEIVnay3BnFPjWFJiOPxheyv+WSAj28HbHq7+8xRHh+SWd4HVSb
UUMS3atUrTkdZ4nE54X4SepNUR9oZKgRcELPRGga+8o1Nm5OxjFv+iz8TQFUBnmCuP41Jz/ji9WT
iSEO6UGxquLTX7CD6IETDoZZZsrVA8vTGig3JIR5YR6Auf4mHjOFyWRpHuglRVtRmgi+jwBmGHkh
7Xi3Df3OzmYNGB2Cdy0OZkq6jbhyaWhrUsAO4x1wNNmx4+5LQ0Uervve/iORmDqpDAi8ECsr1d0A
C4KsX/Gb9W6w1dvytxzRzkD7jOrb5cT/MP6fI4q1NzQsg7eMv2jUnxzSOwNNO1XjCAb5fkYQVTP4
P6GEh9fYaSzc1yCIGyfZGqFM6Hg5eZpT5ZfB08P3h//S+Sn534tlFSdp7oseTV3W4iW+q0+0L+zf
891o++DPjxH40fkNxg2FlrjJP18VKSJYJgUY+OjaXG+AWxa19d73FiBD2Kci5dXBGcekgJ+M9Jlu
1wtHsrM7Aidj+PPoMA/nZsoE0rjNcT27qk9AGPcT/wt/5pLHf65xPekA+gF+rVTXzonMz+AnfW4Z
8u1RQznWg0xPvg9TMHEgpb1djyG8gY+g+rKCAdexwc0jZW7ulXZzYw0m6tfZ8BLVmwm2kFeU/Ohc
TEYnSuUOHVnZWnv0zTg3NZyqAU/ZJ0211wYo+BpId5f8gxDweaCFLZXRgIQ+B1hDski/uslRzq6G
CE1AidjrGyqLqORQF5Ho50LaLQWAjMfLUEdGlJGszGlP8cVDF5e+xNP71/6UOy/gyVmRDQd55yHC
lxAOnJuQSWmrkJEwWDkpQgBkepC7YgqCVnySxVb7K+w+PEMAmaTRtIDutrO/xsP1G05CctTYLQcS
4hzTjEUaf+KyR6x3Mz9OTEy93G3dnYANhcqGp+vMFLLfSnI9VByuWhVGIEKIrxcCv72VicMfu+vq
H15kdtcZpfA7usb2KWIjD2G6a+f0+R47jfo25ea6+XiuABmFJidJPK8LIV1y+euIDmZ/huDFELVj
jAwmzdkUQZWpu+rgLyvRfCTcRgCu5rvKAQ9rzSH1X+0jbkwh6SU5kFC4Ud1gJCk8juNl2y/DitAe
mCQ215g9S6F82VbH0rhR+8pf6LzO7hpug5tccJ0/zLBspISmljGR/j500yx7EsywNLY4BzW0rQSF
FFCPXZoEhZilbFfEjcxtG+jhnLLwtKSDdtmLm/da4+PuceyNaeKHYWh0PLZsfD9qF9TiYd1AMrwi
Jj01DtPLQlwt9EGBxBJVlrLGWLtE9833rdo5VflDF996YkeJm94W1TnysyVVAG7InKLuD4X0VP9E
ZIjIBixmTdjhFs6Df+4pVJ8jKGejOoohabOrot7XqQhbOsHUqwE4cFXrO8OW3yBvKunvlYssMduq
Shg+/r9Q/cGzN4pcpMdRsNzVbqoFBQPPPZRl6mEFr1NDZmhzhCn1t4Mo6RjXEx6vOhHl3nT1npoP
61Gh5DHU2wW4jUlk0az4bZeMR8sdMQLG+DEiPtLodwBnZpDG+Lc262YsEVtAVqgotG8So3LP/BQy
8Rm+yUqEqnHcqoF9upSbZIJLPGFtDMvlpwvKAroGRsBAbmp3oGi+0Zn+YEia5wc8vzi8ZAtRJ0Iu
hglqNARQ0myKKg3xJ4CidvWGJlOwaAvVLAqqZ05IZsMw8yS4RWaY7l7li/H4KbimM5W6kpeX3kkp
jjzi0RM1CFKRMc5NBHL//+je3lc8pKl5mOP2p7J/v1eUoieB3/3Ep9qA7zJwA8u6V4KKUzdqrDse
IsnHTk0JblWe43lHDrSyF8qcIbgaNHmsqsACT9hAsosXDchWNS554u01ouYHsnlJQ7j+mS/nfCEk
K7uilf6rcktjJABxg9Dnw6n/10uS7ddiPAJxnlXavXSzyLqGjfdp9utAfVJmL5ZjfpmIO0ycY+YQ
+9NV+CM63dqMQkCuBszCdb+ckpuIy7K+XIRFZuuyu05lCToh1ZqLsuYrPIf1K0rZ2G2ZEuqYSMD8
Z+06e1/TBw3Z0gF/yMJzePGM1SYJXfDciYotBOF9haisHsnG7ukl8BQgWnUIIWGBO5cPr9gQIXIU
M4C/2SaMHgAc09sjd0pKEDMlo78MdO4TOgIux6BQ2p0p6yazohg+D5hhbwmbTmztBB3ZwWpMDljL
s+hG3k5FT5wjmueLtjSx+vDKiibGDpVYip69c8WGss+KP/IZIiW5IG1EB4/vSLepuVifMW6vc8qB
jSGK7PdHMy8oHmheyz6tn5DXUo0FI0PRllGA/ACc4fJl0GPsvMduLCPKjlahCqUA/iqGs2dkkKmY
zLqt1Pw4rePOmo5tXY1ysaR+nVcrqhMdIXMfdz5AYGc2DJ9H7ObnOupfpZh6cOw8SvU6+rx8zhRB
eB9jy8bMNB7Yhb5ZIVRgSN4RFl0bW90JoGm4zLfLXKGoJvfPoT2tjK5tOdmKmb08lyK5vJCqpPrW
ZYc73XMkB9t+PN1XdrhAkWt6l6JWZnLAxkZMK3htuzqz2lmmgFBwLTb2a+YsUfdtmfJSEufd6Vxm
j/25SKVJUV51yKDXAdf6XTSeGyRiEudBx+SO2JvBZKZOkWYi9OajrKP32WHM/aZ6oPWLO8WZplZf
yefP1HzZkzd4TioCTNGxkNTryu1RYQy06ZLVC5c6753XY/ZZIoqm1e7kchWBVyIL4pKbBlFUylz3
gxDeqTGDBM6K5EvBYH6X0Z0xOxA0Niars2EpwzBwhtWerItJaAKUCHR/T7kUAux7m3W8m+GeLG0a
ySiCjfC/DP1HGasRHGBo1EdeIWYpxjR3z5OHeClXB0sZzsETgEYChCAZcXVLoB8qv8oEPRE/lv38
4Y6aqx/7r2bk1HoqzONjqaJIe57J3m5Zb0mao0/2oEXS2OcUJYhU2cxs48Nmq9fSHu08R0yKq1lz
0SXMc1iRLEdj9HijBCAL0YoYcc+0tTO9Pprnw1zN5uy2uUOo80RZksRSSiVYH54tncV+7MYjM37X
OwhrirD+FEVH4Nlud9E2qiY7XX++/KcXBiMHT5UyPSNNT8lsV5SY5VS0kQeI15UK1EGsW8BqgPw5
HXTdhHVoq8BsvUI05A8m/f7ez1n8dgYehNCKaGXUQfMgQsX3Sobj/vhg7B0ANKCgKn+tqnkKFBLH
J+UJ6KrY00u4HaSpZzpm/ZuTCHuKoaO6BHwG5sKeVm0xluG3UUp57gqsABe6xfhFIJB9CYdo6FUF
UAp3NAvPuapvb0vjW39jaYUHGo41scgOidcliy1fRz4sOrNp1GLFf4IwO7qzfa3Ze6WmHE46yfhR
ltzPodqnFMY2IeDYmsKae85lH12CQQ/mVFoIyqjwFXksJijDfj+SC21N3xvdiIQ+NrxFzRtjLyv1
G+cONYzp9NOtxVnWUV5o6AfkDjpZMZSPJr+RQKREUUjU+0T/If8YVBtEmbi+wEDufGKog1VEkoK5
2+nIonIzWM9MfVql4VzFbu/7c4xzZydDjrih4FISl2Ny1oQO99z45sRw+HMDXInxLHuywXXP/XEN
mu9ktUWNHBjU/6asxYar/HEKb6P0ZC1Ee4h+dyjiD6qgi41ttwc3w8QboQFDWh7xEYLAD5C78PsF
kRcv8J4exZKve9o9+uP5RaOCjCHMMQdtXrqYGrBjQGz1wN5iEEnAQihKUOZpyGbJEqfGMAHqY318
fIFFHHA1UIH4Sl5YZYMrHETSsqhTyBKytKJETzH++iNP721LlJJ6eaFFKJ+Z3Jif6MeujUugl3U0
4TCj4gvzUOe9h4N0dyWJK25oWZUEy4UnHNgKNCIi+6GLA3xZKA/SHH+ESfJ3eA6Nc5MODtXK6FTi
jIJawN5kS+qIj443NB5TB0wx0DDxJwBQK3YsiIkqkX2YJPlzXZbh+mITQMj3pWwOEzsisoCHEu2Y
6XrMPvp58u3hbYKxkAZ1ajSjnBszJciym55nEWuLm9/DUwycVNmZ02EvV2WdXBHx7hlIhtiANywE
Lc4+KeaqOCneFlCih0TfbcZika58GUIC/p8m3f7XBNtgoupIx+6t+cn3PvJLDbVCa5WQbYWLtlj5
vpN6cHNoBxjaWqEXyyNMZ3277+y7CsxhMlJ4eS+sk1QS+4AQ3n8z0xcW3L6wovKSXD/fkNFuozgo
XO+2KOoDDLkgE7QuYnBjAw5pABCIEZmFj4favZaGJUQ6h58tYJOSUn2CKo3VzjVu3w6la7jdbdQn
WtvpyX8oQgT16ehivgGU6RD9Hct2U7NuE5K0QolTNN8VL9SMZEzH/iOqVNRab6CzQPQqeFWyppJQ
Z8G8IrsNORL1d4pBl8BYTJDo3Iagu8WwMczqsw318wTOyGFwDNyj4Ufkr6qkzKB3jMBhLwW6Y1OX
O1SyfxOsBx5vCoUIREpoX0K8fpxo/wANiFqTOVHO5AP8jznulyjx4v9Uto1GEpnEEBQOVjjAuyvv
H6062fElKJ7iV+eWROlIwj0ROdxDVilpHcMpZh5bmuN3hJj49i2EghWWXuDq9RBe0Qi+xC4qgcHt
tLMISHufV4bXoxu0+xnIKB9ny/6Yo9uaQaXahax9Fv4ZpM0SAiRdluJvGCQ3letIYqB0Fs1rSiGA
SE9JCqDo+VYX6KimxdIiL+J7od7J0eXuJaS0Rw82enZ1WcwO7Gouzv+2x1wP0plBrj1zrFuNOMlL
EUlbsGKNC3QFIjYH0I3x0btemmkDhr8qrmKL3FNamKmLsXnqDXSno1Kym9tqMnmAaxUF0rOfo4DP
cys+b83wxLiBNvwnboYOVL2Hxe9FbfLcgLUwsW0MVe0kkGThZs70BviJTw6HKMWWUxyoD3WyF6qU
zj/L8cuikTp7OXhelClOFAhwUJQd0M3a08oa70a4ZG/sBRX3PXT+t2XAqekVPXIphJG9RxwfiFXT
WKoNzctbS/UqKDEvp32l6JBwDttNNXHBdlLLXP5GSJfc3WhxSjhI46rkCmOjnNwe2lDN7NFISjho
USyoToC3HH1XMwinmGhfpYk9r0zvgA6TgplK6QYfizSdptykC5akL03rBc3tHv/9acYpDNz68QM6
EALbuSqNQcrF9OoOEnQAEgTUQYbM9cPWaYTgTk3GG5qDxT7LPOjY7naPg0ek6GJHP4yvpnFcrR/h
xKKnwpLHkm1aWV/gJAhIcqR5+9Dghb/TX0QTkNDQ11sSptRZJ01rYVoLEz57tTfocE1c0KPztJH4
+aL2WwjrxTfhw/5gDmHwUKMNprfnrKTWENisNJvoybMVkr2x8DGKyTwcfEdPZkPxeeLLyBouSpRL
pvag8mldAX4uVFloejiaiTzoxboDSPIh7VpHiEoWUnuMZIYtEpmStmB/b7Hl09E0o5KdT8QwSG2K
tPH6BpUl0B1qyeWNolWL1CWz8mVEO7GEL4Enmb2vsBOhjhI3Hj9rx+VG9nk7quoBwjucgd1glf8F
d1nmct2RLeR3XL6PyRarGkhf9azDxRPGStt+AmihJAHEK2aI2mWa9iLP2oVd+1xcN4b/NRsqE/f9
T2why610NzDiHBs2+9VbvJap6GzhKvre6YGenb91VZu9Kyxq009rqao37L0qlsQ4GMtDif+YpAZe
FDCZCWr/3tG29epCOymjmyyz2yzttjo6SCWkMkInlirEnc3jp68sERZGVsJv0RZt6+THbgc6r5PP
djZ1VtAQDhKmTUsL6/lqhVlcJF80clFdakh3p02BmFO141mL6YCYyG0evvCwRquOBTWSC3DDhnTS
olrrDYSa3IJebgyjz2nFlVUk6D7a8KGs5aTwe5ycTYKB451b5gF0fKWscNYP+uszl2rLVfNTfSyB
blyuUiS7o2fgG8Vf8r0RCX6TgZR75ufE22iYjhoRr+hGhDfSf8ncR5fkd7I5rxmxPaeHbSHAQqNq
DT8Y+9ag6cWOOvBsq8V0/GqqsxSbvGFqr2nPRcMUPw34O986aMY5xFoRDkOR/9Mjb+ZoKdiESWgH
04ntX0l3SZhE5e9c14PXeTAEnLFNd6JqJZJzdGQUz/HXpW66FeN/5MwOnXaTkwgZuYPQWRDFoR0c
5B50ZYv7OluCaSKwGmyW7gFmE1T0d/7E8fejXz+K2ryOG+WsJdGP4dctq2aHyOGUnqgi/pk4xj7y
JHYmZK5hL8xwcq3RjyfJB4g161U+unsdvfbboCxOPVHpvyfODSblTv4tbdK2noMqbfLfPp6Lg8a3
G1Szclf7Fjpv5n1G/IUbH4xsKlilXOPNfsY+vHuArfWqosqVtTCyXrSNZCvU9a6SeiRYZ8KqTJub
r+Yu9ZitV5y/uiBg0VNi2qGraE7sQhHFLD5WA3K6Y/y/p+cbfJHLv5TsLueLZ5LJcNTeTj/ElMDK
YI+0MNxCBfDLvaqj0JPpLpaNLuMAkyME1bh0svsEXswMBTT8plOlAOmn/DYH4IqzDj3VuSxrDERw
hymmbdqrwP8BgcnqeXJHkvKVS4Cm5kjytnSJIeD9weYUWC2uCLp/rRnpfZOHcqolhWsKXp3dOrCK
6e8yaszsBjOk9pAncdCBu3ETSnwD6gp0ERR/v153H603UYmS8eAZZo0evHdppAOSPw1VYiQwF9ov
p4oSo+iXPOg9bSJVUdqU8gY2Hp/H6YVugsrSkTwa5vZDha0qhh2C2ZyT5N2PsaH9glsjfYY4mh4O
6odfXGtqypj1314YKkRspsOI2h2I2kkf8hGLh3gukJDssWfQMDic62+e269nZoL0NyUZdSp9/Vqp
Te8DAQVMbGcPFzIA5GNE5WPVgUC8kWNDky0jmCf3FkTTUC5My+z+I8xO57TOoNjcINdYA5GCswuz
zlLeCgGLVUHf6YMu4CaJU6oP1IuO3JTPISec90uQc7LBFKCoU3oyZ0482RGOPyzARCQwT1SB6iQa
ZXoCYX+vnYcUxKckkToCwfLDCUiW3Cg8hQU53/tPmY3CM2Jtx5uEKNX5CiAUpE/lCEPZlbdaGHV6
ngvLNNhng3XT+YhNvUzjN5FK2ZuBJU+4dm4x225UigB/SZVCvhc6xmqAsF0O5U+imgX0wCXtYCyT
DNGy+QA1sBuiHQz0f2poYwUxantiNd6anD+WcEE0rVNMPfwxPLaXo/dHGUlBmIFUIfJtnaHBNdVZ
GLgN8rNLtcvbZkDJXTcwLRMHjonCceHxrDeMRWgO0S9lyzVZlxRbvFJKEUbHfyzPLGMgwZyV1B98
+n5qqLtvCG2ItpRwYPv8WHMTHjR0JfDO1WSzCaj0ymI6wXy3ytDpFmfyb24hrgkGcSVG6kXpBlp5
z+lVQaJmJthkuO7OR+euQR7KPwhrwPOHJoMOwJHpdtJPIWYSUpAf6Qv0vSzg3fX2Q5JNJ5ZH3dRX
3ObpkMP8CdSw6UMHz6LGuYiTY4svaQJIfLU2rUkkcfFTtUrEM3doZeHpXgUtPXRymobE/LPQdZHa
nxqir3B/jPBqx3139e9xIDASPgGSJJ6Z94T4y3jMKht5WjbmcgnnBzKY3Uqb+0l/gqI5EqduzCUO
8ISesxuUEyMwj/msBgkOGcugsappN0C6t9vYfPcEEMcqRTj3QSi448DdZTWtN1TlVQFbS4MWzlcr
NyueHlXCYu9Jzt+D7B+0ZS2hzmoN0cJAjEAE1R9C5a1A2BT7fFdo+ROxd5rKj4nKHTm/fCOT67Vm
CsgzgDzzpaY+q8GkztLLVb/Y08qQwWwblKrQLrEGaLGPmbDpGLIxl3JvKj2ynxfyMI1h2w5OpeA6
i9psFiQfJ83eiuBtC4cUkmhL4vhRLylBIj8Y5ffscQcPiLL3YHIbhKfif1Ra6gWDraQCynPQYzQV
+4qEE0+7cv9Q9jjX/QiQ6mwwypN+8Z4tnO3scv8oykZZXli07u1H4p22mYDrhXv4sDtx9u5tqmsR
irNwv3fDg9T53e7NP0n8Aib70VE3b+9+1ThX91m8G27xHIP//Qe0yCe2g8gqqqjcyt6ntQnkRrNW
fQmP/pyHUNCi8Ay7lp4AxthgSiKoFHIPBvPRwHsOW/p5/mqWgfO7+NFq1aw6FYs9MjbFFx6KbQtQ
0Sx1Yv8KQcw8AosSp4IbyWZJVH6DDYWMxnPWtMbMy6Qi2Up9kYgnOtI65I/p5Vm+lzyuFqvwOtoJ
+whzsxKPDy1Gc8P3b+CB4FlFf2yY2OPNpvbYFBNQwmQDGWkx1bX4mKAuNkipytBolnj/u21rfnBf
sLyuIou38QJzgmougp0nWH0/Uj9NRcrKEEMhw8rWlrgenbWrEambjXLODku6EbtaqbFqXqgEKnct
zjsV3WkXw44Er6alWoxyj9ObYUT8N8E3RbnNfDeMGbILgPXfaA0tNKEZSuaOVGrlsgkMfP7YVIIn
f9AskWEvzW7FS4aplOE3Zd8rhGw1B0s4IO+R1w6LqssEo7JHWRqhpRhAQk9EjUgO+YJfgLLQc2bg
NjJ0YNLRnaQ3uRw76VjIMH5LyrtysNzOKbE+1AoGZgzHARKt7aO1GSWmOkYLo6fqYorfkcsHXgwD
pCr7rBD9Z2G4HMdcwoOdWo9O1rglKzlSpbP8MDIe2HiD00bqQl3XELQj0pZrrZ/Y0+lTnhZ7WFIB
ht8d2961ZNaQSc6Dtr9wa4KCM7oUSPuOn59d2N7bA+3/7QicLE3ntNH+fPMeGotLcOej1VQiLAYL
Ar07JQSzwSVqnlFvVWtC7NrItCfp2DKZHAeNOfNx5hJ7EI9gDWxW4YLJ68uprF4GHRJIDezoz1PA
qmHhjoMlNJJY44ZbvOc4PxS9w1NTF7WfMlN5/+0S6CeJ7ZKogXBX9l/VnDxd2WXyNBa9vYlnb/I+
CWGa3tFw3x7EbN/u6quSv0bzW/sImAZtPJawy9XySfyKTpr/YnE1j1PqExnTP/DbhzMzProqiZBS
04tGUvmNnlriCZ0ZL/YEteCihvcKps0OEe7dn55cbI57JqZJSE0GEC6F8LoJWHG/6tRmaaq+3MZc
Yyg+PjA7aUr4KgzCWZ/5jylZoaZ1Yjtq+6LVWLKZ9T9D6iIud5qpHeoTP5Blwh9bbnf9axAQB8ge
aXaTrIo5Kp5c6gZQpHtFogLiRgosbwy9l2rLZIkq4i7j+7dTA3QlPTf96g+iUzQoHKtdVNkATdlo
Ad9V4WYJuxpP9dOBPGY3xHr0RdKWhXTa08PJ3hHRPUDxeH9Mdl+DKIuJ5suX+rybxyW4ogIrHLXu
mRallmR2Lxl4RylH3ZPaDBvVfBbQMpLL60k0OO8DfQ15HgAbFOVor1t6yZF7EkXznbb34plgsLbl
49P/WsUqOWPS6QrLFkrmGNPOACnoApUMuhmgCjW+rmMPBWItZ3jjtK8Ky+NBig8dDd5eerrC2G8S
4FCYIMvrgvAsjflB2CBiiwRh3kyrGjWJo0GHEy/yAh7xchDcK/HYIGl1fQyz6DhvZZno24nBe9WR
7IOPs5fDjXSzt39q5CkJYA1erEaBtqibZwsZtqzuSypTGTtnEx2fihaGzb1vl5zHCmtqFONtgwey
gFsXO8vec9eDi1MYqkDDeOyKs1PUPxbTLITwk2ZYr/qct5B1l2Jg+E9mLa36Q490I5cmMpf2upjN
lQhZ4en6u6tV/pfUUmxeEFYEps9fCaH2LptI/ZfkHqy7hK8adAdojgmzCGVtNwWepjghwptQJpnt
5/I2WpzN+DBfMiDPtizRyYaqdR1eDjjiGQaKyce+CgGVErVCfsbe2BXnGd7inBs3qyohLjHSnyuZ
1INjHdz2PjJBjBR8ESAgWY9AIIWKpilhjM7SNSiFuOYFhmdThqNaV6WdmuNhjhhW0PNSszbM8+Ec
NWgXRE8hPQfdtgiLxknoYgupnCgXhn6h6H8qI7AD8HAuX4Mdu0wBLkVXWOgtYlDWBIypFnDaa8AH
EcB6erbiDIp8LI8qSyiHaXWsk8b5xvpMPznXSEaW8tS3fXxP3bdqYhMz7n1+v7PiJ4CQbYUjgoHs
6n2XnrLOZeC7NYhCW4Gd8v6Vut4xzbIMeJ3taRDWO6h61zg0aBAt/EJh1iKFu8+9agHmhxKf8Xp5
qzClwLuZFMNaLOQMhY24siQyeMmlXlvlFlacbfW0IP6+bCTSzoYwnEMmQplhGtaZALsFTjNQutz6
Q5XGHL1f6cdTAdsLdI4/npxH6rIBAS/6jBElNykes9xQIBqZeOq3Q4R3H/oBGSARtQ9JvdqlrPHu
Yw3tWluYNMB3rLUoisWCLIUvfo+rL3V6Jf/6YMa83fRQx4wUru/hpEXYVSSwfu8+zEWSiN+d23Rn
YCDNQidbRGjClH9QPRqWmj4oF8hdmeHD5l+Cab8PL6kHoqLmDJXgV72RgPp9VkEhaxq9+DuNpBNA
f68FZYKksnzcjeQzwymD5NYyGyRw1ChSHzGRxwr8E1dojVp8waiXPL87N9a9KwkHlyxL2gxdcFi8
oKoszU9FgcDe59XILw6EzYgfuqqqSEtRWAkDKKmwSAozln/HSzfsFxiRordMUGEFwjBzQyh6EQyS
m9h56uWCa9zRV2c6OzLj8IWzqPEkecLgJv2/gRDy92JA77hwVgt6b4LUku75HUM7xywYKU5/sVIo
8Cr+igAw5hO3mEZBxQghovNQA0E1EElJOwOOlyLixXW8MfxGdfpiYtwbrBP0gXf5Yk4uYilK/8XP
wDr9LHy61d5FlAyfb5Uz35kNMXiAALJCyjgURzqRRQLsIS5/LS0yrq5pFe7y+dCgPe+FT1yzXGQG
MLyzYLgkM6APl18PX3FSNqlBI4qzYC7onBwH2eTpIyzuh/4sqmdKG696lUN95p5MwCE1/bzRaHiK
OSY/7fIZ81Uulz2hY8ll8D1lp4t4MFP00zU+bYzT6ex70gJdWZo/a6XliV3YcSrqrUTbmll+hpZF
aYJhm+xP6IsZtzD/kw8TA4CVvJpDDW21RUP7ykzaReBBABPCSiSpMOCmI0ASJQuj8cDwoRd2slXR
S3/a23+UyupmS/BfM2h1vGtWzt78bprLQXHYrxJ9CZu/+upCqwWZ5GA+TkmAbwfmfHJWIEmA2/SO
y48z2ivNPHmIQNMhGAiqJBCDstkH+Yh98RzZidjlbKu7SZSTWFSNa9sCClHzT9dylZ4j2jWttOf9
tqUeavfgSogODNZNoE7D/DLOWHj26+f1F2jHYvLinOITwKX/MSt8gntXg5F62brNNKODyd/7EbtJ
Cj8XaoZujAyCjCZ/m7g5FJz8s37i8F1qB0XvIMjesorbetjcUJGcTVa/dvsoclM8+F3oA88Crq0X
tyL+a2T/DqdGfiqE2M/+VdJIH8Tt72nXbIC3jvr3ohFsqOUGlpJmf/mg8WE0xgjSDs4LmztvVrUn
XcMI14Crk1yTW5RfbK5C5Gtj0hByCqu1/D1Ko6LCXm7XhDJKemwJqxiskWiaIE3cyk0xTY0sva2+
rzh4jgaHhxqywhZJ5Q5ycUacRryZIddTlwTVHC4hXuJm7fIeLIqqg/GvpPsBRnAWlcPraDRsuRV3
JgS3PA9nSc6JQGo9XYOKF+rwKgy6EJdcz9S0TzUBsB1fCuSw+fCJQ8HE3B4myrYRyE4S/5CptvVp
vxaticz0uY/9Hn3S5XhkAM6f0L05w8XUfb8UPO4HnxWnbREl0W8zvCwhGjsMQX2Dqu8czXOq/P3q
Ob8X/9o1H+f06F0Vw9aO8n8FTB8kbIreC6GVr9o9jKFFmb9WLXMzHqMBhs3kVj5kSUGG5zXeM7G+
/a7DpoDLqzvp2FGZycjYysyJCtNi2Dy/d6T6HIwiAtOEbPFGYBiywmcrRVn6skChUAPYxRKvivqM
fbFlc4IxHqTa5bfbf7w6W1jEslA3DE39Sz2fF1DrLOFPr/eMLJpBkGwlZOaoRsOdgeGzzx/QgwiU
/fRNJZVy+a8MCevB+gdmZ82PtWA32sQyjDvZ+lsc+2d2oJVRgMOqALtv5KNMkeVwMnvtNQdU7j7q
RrH3Xo059Y2FQym6Go04XZNygyh4GfUs25awmLjl6NpOKZfYRKILUO3SqBei1yRIScvB/33GVpW4
+DEEbxKUHau5vIBQehLISCQXvvKcch/A52BoKUZNkj8LFG9UshgSq7V3d9ZVN3eZaDoQHK/fd+CN
LNeajLtcWHrb43HO2kLW5MPS5SZnr1mjv3JQ8teSLSxJfv9atlYrwGm2BCaro7GtOGz2UnZ5lkMa
7PujzwrjVDcI5Es2H9LGBzZHNwJ6Yq1Y1+fAdPLvcHelf6jiAQvtuFYurYUES3E1y2v+hiPykttV
4kZzDwUX7l4M3XkSPj4zhN0p0jPbSrZSjw6GJcxJ4QjS8s7QtoNdDvMrG9fxBg5/r8xT3PEyz6R3
N1RehgmfSSLjDbKfuZXTEbvPL2q69ZQpSkN2SFvh+wOmEsnuyKsWy6ZCUcwq83X13VtIl+pPa+lF
+hXuUbWUme2r0RzMDxTd42B8twY8RUVWfVzj+1TPXrB89VQF26uQDz4VOak+cDLw4NIISglfgmux
psxL0gP65w8lSNKkI4UTI5Gp9l9Mcr2fqyCQ0hjyy2JyDh2VyJdqMJr2duaIgGEEKpYasOPxZsyg
8Gqi6aNC2yfqctz5U6WdougwoAu/7UzQy36HTovzaWcB9kvrDz7gHRVuvVmg+gAeA1Zz3qvTZiai
dPHi6O7CEi7cURnXBnJKGA/0SKmoLwxVx3cnIZGgxy0xes9CQmEvyyepHnJznwzPUHDEnVmNwH44
P7ygFYg8DiKD+Av/Snp0JLUKn7l+gxAQ0AAc49hTA7C/E85bOAMeMTDU1PwR0mDVOnfOH8Uek2pE
YWvoNtBvQIGYC40BDJG3nWpMf5cLnVlkaR5yKpqNC+9c2DneSXLTlzhUCejtLpf7t1VGDHrYx7GI
MrWmxXuC9yFJysh0PSf+vC/yzqAzQT9/f8GqgJlyktahaTzbPEQHbVe+hbQoCsa9U6v0c15jlbID
oXcz7r+jtchX7EaRrbg+3/SwG/pRJwb02KQuav2q1syOR9L8IgFGhuC+n+KCuexBUUCGrZw6Nj22
3TwnRdxd/pRsnBlFVvxCuDXbmaEJzFXwQ+JXCbsiBVi0XRWK397Ng/otMFwnzLLrtZbojoHSgqOf
nE91EsP31C+CzZ4p0LVtB6AbbPbvgy6L9t/B8XCpWjShmhCGK3tzSUJdU/A7wzwraD6pnDt2xfjf
Y5T9izwYQ32PmnsXik17Ea0m4RVubYf6yEQ1W13jRhlEc6xGZfVr0Frwjh27hnTWH31Bm9/HdYXP
MvvV149HVD8TBnJAxApCw315dV8PY93hTmvNx5HzRHrQba1Q+WWesWG0dJTMGBIjMj4N7nR7BlBU
i67jY1k9KAp+Mvzfgw/eR5RvI7KjPcvqanYhNOIHRWV5i3zCmkMGqnngTxylVHZhu3V9BylgHcG/
OrRQssJuiQpWh2QBYSEldD90xdFvqAr/8rhIQ+YnfTR+ed0iPiKvVAKBXYHxcmRVmdPM5UOBQ3Mk
V1PZ84VggJuOMJmzDsQotgg76hbb7/iltW5tvMW8Jf5C8g2fjFXCFv5klYcKR1FCCIoBODWg0OaB
wRkuI8Vt/HhkvvOmcekF/oBmtC5ndtHNYVvQ0a4DHlQoLth/SDKaEO4tJhR6qLc5v7+AY5Lw9e3w
qtRWrjTjkGOCKXZqWWi9XFBUrifSOUCE6ISEiuSpuEaDJh4PSyjoJvdau7Zei5XgZiMR6Nu4tRpp
pKKQo7TwZCRioU1qs3SfkN/DVbwa3fJyFJtgtZtU5bXqU3CSs33khp0mQaizrH4sWDd7sEAk7GQo
2D/nRj6kmFnpB6jma4u45bG0zGsZw2lVoQXVi5vOW/L0EfFlfFPaq74UzICog6yHyzT73fm5qFvT
Sueoijzdq73WRNx60riM/Ikpkr/Q5zxiNGizvtKyTWC4y/zxBWcXH1qlOJ+gKmkNHkR/eI3CAfVf
TtimidRxVPQ7F59P3BeTBEdf81dHo4GyGDjH6UtTwhpQgt0yQAPJZnvrgFQZAvuCAUHbssfGIusW
tGjzyNRfJJ58o1yYKJcWzS8Xi0ZoAp5mBZZL1LpgxzQZbFBHkN0fvcezglAYmnAPpXY+VfDrwAuh
SF6hTlvDjYoQawE4WOqmH0LGwYhrPGil3zPgsIth7/aHdN35sLxU+zxDhjCaWsqRUtDphMR47vtL
5s8uvdWRIGpszfqftBCPlXUe2+wO1fIaEORVu+0llZ0l6DFHR+TLbiau/QlBo1MsH2l+spiug/aP
HqM2H1OdJ868Mfq97NKD4a+yj4pVxyZYAtXrht3iYE6dpFSEwGJc3PKV/DJeUGGnv1j+ahpc/rkt
yac9ToiGeK60kyiikZ0/WLBucKHeyBBqvbO8+KAsPvPR3Y+RFWLhlqPc8wDREaoSQ6jOEA+JzXJk
9IKFx521nkHW1afEnbas9A9T5rzbkB6pTF9608qFbPaFBZIqo1TsoJ4JhzupLfpS2UxK4oWU8S6+
gTI6BblP8f+N9JgMECzgFsR5iL4BJdHjOXyiuJK8EP8VHXFqKhl2KbWOUXlmC+wapbdsFGouSXVQ
3c1vyLQQzQMfUJ6U2qIhN6Vh26DSXX0Mw2udRKW+AKU2azvKsndt6CO95gTI3e5VsrhoiquFXKp8
YK7/KYYQQOvSupCbgg36w+FsxIdQoMMpgJHT1LaPS4H3/RpCEF82iS7LjvBc3FoWLUv/QNqkpsJZ
2U1Y4Kz23B0xKtqyy0KmsyQlAWqHDaced9DJz3khckYXDLJOgFxc5YXYc50XBsvP9H2NnWn560mE
FuA4RXok3ss6OeOIO9qNwiqGMlN8YchVkzXMxioaxZmuKAWXfPGbqlEk6Ma2dyK68FIoK5yoOnhw
vsYBzpQtwzKgZpP49O7g3k6/3/rPuRB4trbfsg+KmVzF20n0mNCuPMiU1M52bkElG984/JT6mMSH
eIOvZBW3FJQ/XCxmMBWzo/aajlGUuzJClu3Yn85ofMWo/pGKdLcpmAsWqSXWYAMbEKBUVvH++KVg
js7t4GqzyWZF7kYNu7Wuwh4jQLuYe71Kpu5eHOdEll20T96x5q59gr1Y5Ghbni8GiPhYJwCBq5/6
Cmt8vPjSzyHQjTBkUy5jm5n7Gmzj02BOAgd877C8wwFudep7/qOCpfxYPgKJi4IuKvqxIFdOKyKs
kGYkqG/OyZFtOqdsipkC1rdRtkxV+JeBNo7rLNoWVTQxtHEMLUA4VMJsfelvXjyps9rbLC5ahSLM
GbUaAItEpV5wExIC5bE5s0k4zmwtMVFefwJ391brE8IsFCypNV5Vq8Vy/vOgCA8MzJPPrBr5aTjl
ZeOZUCmgKKVtw5AL1DqxXa3BUSKNzqjzNN3QINjUyoTZNlCHc4w4bZnxV0pz2DEYjrrZzJPMSJEp
qvtOHV8um/yz5Ie9zIWh/cKTaZUxj+luwealDr205qhK5PCt/shd/rZNjGl0vYU3SYYc7c0lTnjm
GoRwn+znfm/o7YEhMjFHHnmzG5R6ejqMThVY8SAF9od3LziibMEvSGSIUaontIMoEPqygvmW4bJa
Kw57mxoJ9DrQmh9QsFS8sRa3uBtdBIedFBTqT1z8+6xnCW/hpxY4lVE+NOML16lmIeIsAgywKzxX
ZwnDtHjkzrNHFcvGdNVTPlBsMF2vc2d+O4irbdGFY2gB+xP5jCUezsQYu417/q6UXbYtnSR9IZVu
kLjT88BsRlxocz/kAWA/YU71IVc5a4o5Ba0QyGI0wBoo2owUpEGru1eYsIdOlhmCZNKPLpVaHq6j
TLDtDZW0TVWCbBPB72ppDsXyv2uViymNcF60bcqC2ls9WT0WIfh+/i86wFSUdmqbnoXyhkJJ9a3m
CpPgC5rCj3AZnB0HDEzw/LyzrEZDdBPtTuAqCFSrMZ9MEye5M+blfCqy2s8m1VyYBMagXqo5i6qT
ZtYY9GNuRc6kORT6ZyG3Fss7qIEDT9XaSBFq2yDtDxcVLvmV1iTtj6p3pO4rENO0ozWYzTuad/fV
ZbTHVfkau0d80ls7fnsHue8whJCLENf7jKCtbrIO0UGw6jAcw6UVeRQfx1l1wslMssDAYIEaB5U6
NnVL4eoEqOeF3oW9x/EO2NxssOokzxHxg0g3fN1aTkKYHnKWLfM0caO2YHSbf5CiNWJTXDKRvuKX
9Rwznw+/ias3zkyGY6vABlHCmLveojmqM6Qc4zx4edM3ZqpbhlToUjLoXBLGonyrTnibB0QUfiga
d1HZPfrvfoSNdhGN54dcSZmrCMgFt2TYjf3xPy2dd33oUtLwfd1LVcU+L2+5dVYB927/wW3MCDjL
YPMqvpbm7m630XhTz+gIB05Wt1M+EWR/8QHCbDBFs5WBWad3SU0lTJ4G4/LmPiaeWhhGozpR3/Sa
ujIHzK+1wK+gmXaps3PAFp6JioQYX1ZyEhOxBv4Knz7uz+O+AD5assYB7Dpus1up3o30Eq6I+2dQ
IXrtf/UTdyq1ddbJYyKH3L6TYpgnk7TeU2rXKs4G/t42B6IBmfImeshDAH46VpXsjn0xsU1y4lnC
xf0i9beIVko4nVuVs625STJvsSKHOVP3szha16clSyiR0hO2sY7rTPTLoH9Ab18O5LbCRyV0tUkv
s1l+F1phUONqQl0sO441Twx+j2XCd2A0oojf8bi05lXE/qb6WfmDfDHK7LGY0JVv3smGc/T299qQ
WdsQc2Mm6bUTw2yu6yewcDA4+CDeCAoDzYQbY1jnK3xZl6wI6lP8XcZSmGImRGsXP5XGZ02v5csg
7bGI1Qa+gfFmBqANZI1Hw0RNXiIOVdnmtuNt904P2LIy3PISKU5R4J/AgQzX0FGFfqcsDeM22FVD
6zVceIXDR4K8Kw55QjM3nOUXGy4ZvtzTePl/aL49ae9z3e6gdHTwDGkuq2pO/qrst3t/NM17Ae4x
xNNJUTqAzhQPfSAuZU5j3cixjCyfeaxjdLS5g4Eo8lBxi2MKlbqRt/SmBwSWXP/sLuW5mvNarJb2
eAohEKN1aj3cia/0HZoTqkWNq5J/DQqxldsizlJs+N1andiYVqii5Q55cbkE7Ne8I0rvpfmK1pws
0otgTWWx9jboiJh9+nKWaOknNgbN4FnOfXXT4butGnWerPP2GCHvNH++p68s3x74ihMeSVF9WB/t
PytJ8X9Yj0i7QDvf1w3fOYe/JOnisqo7dQNDou+wB2NIhRDErnsLBjFBZOrWnaDYHG14QWWXRksQ
CpLCwiONkow+W3E4kktrgh+q9g2FQjaTpHQWNKxe+17BqM7AGgOhe9uoITdv7H5kwaiAd7QGTNA6
Qf1m8EVtiG4e6/f3nNDMQ8iJdkMdfa+Q9slNTuZSAWzNDE/PCvst3NjqnMJSm3B3vizglX+e1Tav
LPPzdyf4jPQ8PFO8tMoxvXbbMiYF1dX0Ao+5P58sx5oS0YGUo+FTeLZ86bnTABYm4Io4lGYDUGEp
eSoA9W2NwRRgMC2AM96f8Kxk18hUE3TnLsgHL1qlym0UZex0bRGBcFq0x8VSbhaMrd8BG0YoA8y5
IPbvZ6Ds8Lgs0mmkoxDZ5FCt/VX3R0aUNDQVuyqJlV3jKMfK6q3Nfcz5nxoGM0w1UI0o0DJ9dDP9
hteTTqei5MF10V3peG9Lx6kHhrz0tllDC+okUCCP2kBi3sEmELzuyeoRf+Px5rKa798D7OrsSedX
y7OpakMhDOSGxtY2uSm1w0NzseyXo2mKdNb5Pw5T5NtYnxwFcTO0ZfnRieUYbbVe3KdlCtUOa2ZA
cRqzOyMa/uQj0C5u/H5XZiyN6Jl8pvxLaK3DX5OqxPYwy5PPoCRFnkEMCfTcDqiK6LKJvO/GHKDK
2AGBBeTPWTKbfFGunmqIF5XcHCHUVF0SRLKGZ5YXQfn/BHv7ETJ/xjEVHZPOf72JynAGe6HXiCl+
JYF5GeY85bieFhi5cCrVXKVaT89MQN8871FO4dy/EcWUkXxzmweP7Z6F2LfqmoJFeTyhY6kva/7m
KqtglR4Hs97farUO9G6UyaDxquPv6zyAvUsCpOp2VR/kRP9hpV71SjOSPte7OuRNIpNV7JQdJb5f
BQ03X4hN+xYHPbuac/SPyAoAuQV+P4l1VJeYFjC+/rOM3hqTqFXmoBx4/6S7qwz2uFsKLe7aRXEi
Bs9seBuirHtNg9spbXQC0o7CIubBGfZEYPk1+m6eMTTXfZ61YXzxx9cE4ELvuOShUg6TX8NCshEb
0PcgNzigwSXI2XgTJ3tCKLjIoMWRQuBRTYkgo0hQPVkQaKma/yJFfi6jwDmoG/4/tK6elwjKqsw+
cNmdTvDz2OpbBu7jwQlqy9DvjVCbbPXBpuS2qY3g0kCpjHp2l3oEfbVQLVxVVfvN3BywbpEr9ugu
EeLHOFWYrykb7FtArc3jVyBcBBsMkEzAkItps9aC4xcjaOBND1zuv9Fi5C+ONy8R6khKZ6IjfyqU
lXhZ/uwQZrarHkUVVEHvb3KMyS9IIG3Jbv/sNk8K42xGal3rL+VA/NBHDWvo12L69v95dDeqEJzy
Wc24uraez5o25GxdtQcLIXQMPBKyOk0wvctycnCKWcu/WYOKA8TLCtjxs4+BW5wElgemFBSjWzNV
R+wmn6bUAFbNk+vNC73NieSZTO58i4kdsvCTkznWGOOsgBFv9aQY+mimRF9HliTW7DcnZ8HB/pIi
n1ShhbIoHqrBrfmdQAaHTYTHrGUX9S82GPqf6Kx8c4rXkKNqTBTAEcfSct7AEpJaD1SvANBuUTbv
EPu0DPWwLK3AZz6slQy/zO7tsJeEIadbZfq/eIKF3sJJzPgrTVnB3AoFVLoDR/k/vX0GsqNQ8bVW
VOFRfYwtvmMc8Ic7SQrARt2nQ2vOLUcMSmjNgFUz/O09QUXbmUUxPpXB850sNGDEmNr3YErcqimu
igw7wiMmWtggx3qmf01sr7CdBf54nDg3mXMJAiz7KUrH6Y7KCi+tC0ndXqN+AGwZNlGIhrkayXM8
xW1lGL71cmHMJO6MG3jIXUJSDdu/OV1nLqUpbcKA4s7U0Pa94oQSWAOZQyMfT4/8EQ5HdeiGIBta
EMouWN51pnOc9s45mLVhTZue76CIBeX0rsVBc5zLMQWvbsCm4dcakQfR/bDCwhHKQwI9Coq9dXwd
dhfBo1ED0qOknhaffD0Yse0CGxA+TZeWhnE8vztF4eS6eeqvUrw3UCtFYXikOgKs/Fu9Oh5SccKu
O7IU4xcdGKc+1fuH9oUpmbiLRmEXVKjI+sJrRDi+UvveSn30gPRraY7hsmIOZtQxoJBVj385nf4K
iWjSrIRVUcl3DQTNp1ZA4TKcJWpN7d/XB9Z9KgIOxDIYZH/uIlCjM5RYydv86Gh40kA457HXMbYh
oTDCj6Nvlbdxy4U/nTX/haqkbKRPc/g2mhd9NmKrRtE/wQpQAb7216nktoiH4XayFvles5ngDoUC
fA4dWjyOCZWvqxaoYnDEMLfUFJHwEJeFTHJVn1Rtqfd1AdfY/Y9TkxfNRRT17Ea5+KGT2+uRBi2M
xN9y7oci//9iZDcd+ny8xppoNGIl+mQqNRxHUpT76q4l/6FTqNu2hDPVuyHKns9yScX58EA5WYfo
0LElmIVCKH51KzEYPjJ2cBblBhSjKBM1sKTHALCcJJ18D3OdApPGxFka9bwkhjDhZhddP0wM7AU1
uSz2tEQmVDuV9V168RORgTtqr+gFLZLMbiwJLxcdJRoMSepWbmUDPJ7Oqk+0o5oIMmca7Ri9aYc8
kCIXdo7YZxGSgSCiMdlx622QVeNm/Kvw9VUSvsvtCjvO9oFJq+A1OF4YJtppgyFX4ulpF0IHy4Ti
cFTDQeNEjlaCPsmM0pCIPoJN7wlJ1jIICqI9TuOwxiPFa7Bv85VG3zokneR1LN7ci06js272MOGo
Eeno6/PYX4atz/MLECXAn/iqKmkgFUKhxs7DuXWNoM29wyGjYxvdCLy3n4JDnTKEVQYTEKQegCt0
kXhhRu0JvSDb/mHqMD6Oh5P4s0sTftwihtXD24BcpxzdmEfJPR4ngdgJbzbemiELZduV+D/lWW0O
ZjFhnT2oI0DnZUEuhepx7GvYxJorBBuiNq7u8WmNDm52CdQ5Qh2nwiyb2TidmhUnY9kZ3vrP2VNi
YqbcH+oPLxFqAeeGQBvilqWFisNnN33KImRCsSKx7CG7k1v67vsxjscAQIYLKostafUnjartZgAF
Rm5nFYLo0nbh3B/lo9UF1c5pS/ibVpnH2GWN1tdj95tK8AwD1ycPyelkIEkKVJEZlRFiBAjQTjdw
mYBlpg9IS9iTH8e3W3kYAbwysUvpqnxkN71/FpTh0zDCpaUC79rRpeKQcUMysqfpgMXBu9I5kbf+
hHrQjWtE6cXUGtGiT72QeH2fKEwP00nrsdY+mwfTM5VKQDMkgPns/Nfstbpc1omcd3UAY379d74w
Rl+tLJjcgcnoPCRtQ7YSiyI21K6cADmh5MGLYUGS9QkR4BjLX6l8y/v1KOMOT5QsXXigaJ8ZB4VS
f5pWzk5FdVUxPp0qHb699j+/bbRKyGF5uKrl9XDDIZnJczUJkB6FC7LT/1F2l8c2tRFC+ZT/VQR4
oTTJ8Fzzc4chlyRhBjWfhwVuB1ftlL7KnVxEFgtGyZHCTlWj8ZmHHcRogoCv7lxgPGu/t3PDjY+G
fXmar3C+V0rOTfjbfQPHsFJ7U89nTEbvDvMA51CwWvlumRH7+X0txUGa3qajIemrlSepqh5EWLkP
SF1awnTXTdaB8XZ9z5mg9iv0/sZ4JczzfvAZyyNEN9M1aOujnVs7YdKXwH7Hz59+5oXPxXKsTzOg
+4fH8neNN/fIxsa/QhMD3KIJnxKgWI7UpABHtLa6FhYSxKSj7Ze5BXAGrRmZJ9TBr2DeH/jzLG2F
4K9i1Nm3EbFjOHOvWiuOV25kDUJJMnQ14dGR5jO7pDgE48EAE/bKdZPw3xD6hAR7VrYUBDabj6Yt
WOXwJa5OariqzfbuU02gmQiiPcWo7eTbpziGgWSmnhQ/XCTQ3rBgPd1Z/e0EVVFk5mknZMGdQYce
9vt0EqEybUeReeL5KMnDYqM1LEpGRHRV0ZJa/Nmz9BFx/+YZ384EOTKEOBa8CrWkjou0b6uIoh0x
6U4rElu6k0P4CNqDQ0649EB6RviujS9qF3j5+4p+bkuhDnCjNLrEdGiEhpDZALZDyVDEuIIuEMbE
r4Ry+QBcz4wwDiYbyR9o15W71i476sGD2udwwlmFbHqL9i/u39ecZjjWNuaWRUV511hqXbVew8eI
qJHiRAnyKWh5KfJRUZtpBTN2j2yQ14nzimK3XL8ySSvE51Cz9q4B2JCooatJ+IPk+opo6ftCeYVc
Za74d86gYr2xISjlGHVHALOmANOKZk84RPXiB3BPz4KuhH+GbLQBdKuC3oO0RhUNaGb8arznExqz
BvLoKwqRKL7t5P7BREdvoyvrYfFc7hDpdFKhu95R3wo97aOTNkEhwnIO18LaPPch1GmVJJR0gFbu
5uqHbQ4u7WSmCy6mChsxUgD5SekVD9F8oDGc12EXaJbf8NTIS+iikcj93CSm4VJpzyOcaumUOgk+
FYXu1CMSymdp36uouiuHiHlVNQRsKTRhBl3FRSPimTGelchpTUynNArTWKCj2ERKBFhKWDEOrDrO
OVxj9SDce098hbbbmrE7f6ByExtxZ0o+JcMZ/w1MitOp9+cKEI97NGHcv14ydey2Msvu3sLs/0Mi
K7s3mWfLr549HuWZVjlloeNx4cLp7nM8qCrcxYWynMAPJaJBqNgQSlIBYC+F9hXIPqv7m5YgYkwi
PycIknJfh3w5jDcH9JS4STQS2bJjenGBsvVuABOoM556+0aFEiTQYj2TaJUoVaKWIROGf76OHvVS
ZXk0cPkl9df3q09crjfmuIxC6JmZD6hRm1kJ62bb5rUYCK3h+BkMVz4an4CgwAXoI9y3U8QYZyr4
4Ak9Yqi18SpIrcn3Gdo8zZJiBcOJV2Pe075TcJ5HsNh1o+nLwt1j4/2/xdNrNUmkys/0Fy7pB27z
g3cb/vxWTmpD9YgHquVXaSA0/LX4KHeAm7Aw75JPBFDaOphn5aegapjw1309cvtHPeSM2hU3zWgV
SxNnRZglXvmLaCb3AhzUpi/oclRgpm84ZrQWZUioLHfimd0PD5uYoPsTz4Aqe5z/wfCSCRTDKLO1
/sX2hJO4dwIhWRAxqNrgkXAxwkQXyoT/dgSXmQgaPR4CS8i0f+8e/OgGLiQyk+8PcoSx8s5wylmk
Lfu8W/buxncGLq05lS6ZJZbyeAqhP6cGMWEAurBgX/xgmAveW7CsLwUZLu17EqHqc7KG/5vIqJU0
68gTjPdK6wEvftJpCwx5ymK70wMZCGCFd8IcYqxUjgxHyAcF+y/DJzEwraKm8dAUP/7GMTZxuS++
PkNC062z3Zt6V+0HfC1AsZS2O9mqTt4aBd93C/YrnIsexZdwf/MpY5x7+g6zMTaVbKMMKc0rf6kI
f5pEjHu+GqJC6qh3qeISQb7NSpgWiNqn53455KdESJUwVpC7maKHFU7ZhOq4fgu6ZucAG808QZtL
hp3IU9D6HDidircmLf0b26OVYKCRoFYoLrL1AIs6AyVq0RAh1m8G930E9Dj8+RGF3hJjYHxm4+a/
mKB2DwkZR3S3j+FtTuNosGQn/dkGt0r0oMxA38j7HddDVi1nW6g/jTQIrMn7cjN1KB55wk7G4B31
xmHH8gLdUprb6uiyG461rb92Iw9Bi4y0icGlqcBC+8bS/QTuq5J/djbyKVOrGjTtBjM/ZM1ig23E
8rDCOzX7lXd6to6Kxky9NKZX+5GoZ1LWsRVLfcd/wqJN5x3TO4anNaitb5lXw0RRll0sp1Wk/rK5
sFOlqKf9kuooWNkQzLVnbd0yjPnuSijSOYvirLd2hy8IE6MpFst+E3hpljryJIs/lwBaOwo29KYv
+jxZtAWb78mKh5y4mRfb8AhCTBM5ZP2/JiZ1z9SjDlybqihnrHUvayFhGQCYYiKo+EBjM6SuNbpI
drtTXzQM/kaEHgKjM9hK8rUzp2R2V9kcSg/HJ4SvbC9yRAAwz/vRffD0sbsOpzaVXCQzsTncPOse
1bn4MbotJYui2QGNuHJQjiImH4WciVOIQumIviZWjsiGhsYFaf1gHVTPbKNrHLsnV7sZs02J+Tj0
Q1A2jfHxXJVqs35r2SAs4tK7YXgFEk1errdFTdmxuoZTW/RYY5GD99ceGg/rdUzsslY6mmQoYYZd
e4qOOQklWwLrks29nH+yJqou2xqL1YA2J8TWJHSMLslsvHXlI8km40SBwiYBJlLfRgb7MhDriPpb
ge8Wb5T5Ye+SuVLt80sws/mukmnEt5tuDLra0BFbicrU6RzbeZ10Fye27zuZzKhP27TyNrOgnoA0
pPd7sOAdHBzkLx2aNNlaof6MgXd2hwhqvKC3FFhrj+ZqvqvR9rWiacT4gdZOM+qT2t8e+dqpYgY7
fZ/F7UlvkCIhATG4LFYvUZyF65CRb4bFr4hqWynZAMTDEPSyx3l4Nlu6exHlbtkXefuzZ4ihjjZY
xoCYABrpihNhZvM7eEOGjOwsqNIKboUEb/p9O2v5+uYK4G2QKST91m+1XpkI9wSt8Z5NUGZxnlUf
3SW36J1gnVA/INtnOaOu6qvCO4TkOTZxiEwsxJGWUpG+2CW5Vdqv4AEvHlQRWBVKCfpX5n2PMJv+
qGwV8Horq467Ok72CnA90Pf51pzN2WkSljZkBI4UCXpNNL/6+QUpEcpEHylBK+VOPUQ/OZugiqpG
pNlFIIH5A1jWe5zKPAm3L2xIslToFT+OXoocXFqShLT6gtwGuoPEWpDMDPOQnoGCWAaXmUnPssqe
iZy9q8bpsm4K4bHD/4ex0fQtdLmgepXXOPH2pQTPjPOECufPFJnnjC4Z6Jwtp7dxE40XhO1yzPQa
tGVtD0jcDP2fnBByE1rXd1i8UUJO6led2NCVTUrAKy/gR+0xBUU7T72yTQhoj2Dyrynniatjj5+F
qvur2FRPSeP0xKD9YV1Cfov+hPKYMKFadaTXI9EQpNf3qYuILmo+YcJ8Yg5h3oduge8Vemg85KRX
y417XxwcnXKWPjUatdJ9iKP4f5HRhtOneDSizKxs8cdSEzE6tauenyQQPr7E655FkokgFLXYnWdC
4lLXdQVL1bM41aARLZ8WBgQ82XzsrD+1yZ+tTi02IeYc1vvTME7hcGCKF0GLrO61vGD6V1e7fquT
5Ux7bk1IPIe0olOzRVIaGnuhuFELsK/zuQsryOMzZRnWH+WtvoXHy7hlWStOAewMhVXWboc0h9XJ
2hNokDAT2QxpuRMtxeWJ0q8VKs0FBcnphtYQQ5M0sgAvj9gf2Bvn1ill5PVPKmNAEJfgezG1nMV6
l7roInvdUAxCLmFh4SatdzzJkfNZdFGlEAxKLan61or5sgLA/swR+IwgoEyMnfdJrS1BSEERtAT7
Ubq7OEVENOBq5q+P1OwSGuvmItYsK4XcnJp3XjnMZ1wRk7Q1bBej3rx1kh5C8a7q38R1YAvH/QMJ
ObowESQJcuCAFd7VoXkkPqdiPHCUt2vE2GlZ6wYeCJ7rIH6oz/c74horthVTD0JFTrz9LOVIkRor
v302m3SsYTdmtwXXvSNLpuFxsuSVKmnLfGb9ICYfl+2ePCqWN36y5f7xM3QprOFNSeoo46Ad3HsY
+vUGhhuDOPrgAKQsFjRlThIjRjLW2Vhes/MD3WjO/B3xi6okThdFjhNWKzwNjX3jFyrOWUgthM3X
IwqWrSdClLaA8Y8qNcLZ5j2Ds9vQcdVQX1htEJWxUcVH9URD5e3vRCny4T2Jod4b/ch3i3BxC7+R
d4glcTBGTE0M/bZLxqeqNZfdELRu1gRcMYW3Rao0HF0uaRkOZDxnroULI7mF6yRhEdecNPakQdDw
rRCqFrgnwIUVm6/pr8OLFQfE2ICcz9N8NtKhX4RkKWgV6gllMmhxcNygYoMl52gSEHMV9a+B2ebd
7qUUWdTk3kyepMUyNysC8YsUVZiMbXIgQAyqIB1BQbW3dQPXMJAtVrseGFZCw876lpps/VAoQx6C
SKHdcH0pUtrN5qYNz+J61mbuJz9F3AwjVRmaVblEWKBJ2z3O/OMtIo3IA0a8Iu2PM4Mr7ilzA7tF
0qIHVIcYrRd8NnYo9MTKIfSuEZM0E2VrPSLoaOpvUyLhYn7XDyOgv2pv4/1Eb8HUdVxN/ymNXLXa
KStC/zYX8Zi8Jcq98ZQgijMCRet1Crq66T76/T/nlk6HYFTDsop1M4KxCTWDijWO2sRU3NEqMKdV
06UWEiuYn9ORrYsDXaAROGBQMZjRIhlbbCfrkThw0U3Ei9ljGJse6EK3+DfGahfY9cnVXCAC2dEQ
diO2hf/T/2PqvkERBj0nRj2hy3YJ1gvoyg0ymP+ce4PAcIdwvONkQSfBHGYZ2c/BCHO9l9H4RfO0
oRb8nu0OaoPb6zvlPOP6HJpGpHJIdaTc2T9M9tg9k1yhkS906oKFrM7X41kLjC81h4FpUPknG9jW
h9opDFExoZAE+QLO62bNFSu5DdLR689wmuknTeJwKSDqZKNZ950L5tt6v25t+nmJglWqP2DTpaVy
8f2xPTe5s+cqO+PHcMwg5VETReBY2B8fuNmZG8rXcLBsiURGArV0bJApqpf8G8b3+tmB6sTyprTB
g/AbFwZEKeBUPcQxCkoatfiEHIVE64XX+LsgW2WwUtxPhAL7VuaLdJQFBWjeNnlR2fjxA0gePih1
irjQl1US/Ldqp1DMwP29dzfIQW+4O8zC2Eo06v4bXzC8P+dXKQqYzLGrsj5hy1+GXU80DvQEv7k2
qXPbfxjNy0CYmfk5tFr8urWZgOeK1HlwpGZpHf+brFstiWvv7mJzMRF7LWA4m67BYAZLsbhLljKU
ruz7rKoVjy0IGlCZ4nE7Pe0STRKNeXz4E8WDG4sappmEtiYmc5JcV5WVqV1jP3dnJaRxjMZCCbXg
sh2v9MpXznh16Dh2AUwvD06HRmqzHzttNsADQq7V1/idFE2jiS2swP4ADLVeZInfu4XGNxq3BMv3
we9pytEHss2zsO4Jxlh+K0vdAi94lQQFwpLJxjzhyuoLtEudk7avDsxbM4AXl9D6zI4rESTHi3Xf
RIqDdSKiDttS/Cbl9zwOJ6PiYUu3ow6v7CsaBNfWcsW/QrI0Z3EvrERrqi2p1j09DbadGesXEq6f
eTGufGxRVriDPUo6tq6UPA6jKJHUzPOlnL+kgVwh+NmL1HryQhbYsmiLahK0nAiEPFglpSV+QQo4
8TBlziuvv8vxd+nOFzO5oqZmzYR+/TXahFd2h//Tdf/pAHPJELgRVCWc4iP8fSY77TkO8hRmfBTx
3bKmfz2NfEwgWDYDQmeEc2S3GRrri+DG7NLrRZTvXrZthej7uQrCH91s30Gdzz/uVt2ZausqMWbX
foBiSuAaTCCacGYq86X9dj9l8VfvKxJxzO+CQZ3NUS2CZNhZxqGA4XeOLskzbS1/IpCupky3SyvI
+0GV8CIMZgGebe13DrNFg3xHE8f8/vwU/B5I+tgtwePvmcN68Juw01QIVExVvNhZynzy8XOO9LqF
oECDyJOuwO8YrIN8TeE23C+GCRVBMpJoVc/1x5diBMlDn2SmDPFWDQsaUlIn18Ugjpv6AS9vXPEw
TwC54QOohhgvYCfXYGc8fpHjQK3mGoYBuDvhKy2/cf2fy7Rdnvf3sqvMIwhIojEAHTwW5errWsg9
qxc0kYoZlszdQRTBwM02sj5utzRzEt/P1qG7xxGTfqDuSdAvF3sil7xCHPSm6lce+p2ZabZ4n5wo
bN73j1dWMd+nlJm9HQM4oiDP/l7Em4G5z22jpFxXiy9IBO1jRecVsLZ4eZlUXpSsTtiqaD5TP+UJ
F3qY01lZpV9hN6kbHDztkGUcwwFb4T7wOIugJVxBKZ7nJIAZb9U2Mbvo3PVdZKI4nkwPBfzclGrk
ocXTMFL5bYZtU9pgPxkNq8V4do418uXzaQWij3sVFweI5bDzPtj0cXVTJ2SgwscstO61BLlHlxBU
nnk6WuZjrYj7egrWoffDsxpdvzqZB1DEKL7pwCOFdS5Dgv4VZOv9a449us/qMwa/hyhWCjthsxwl
2DMIvrRlT4d6hhwSRpbMPv7mxdTUXmWX1VDzVNMAmvq9FMXEOIFkmYMewz3moGupopyCRnrSC8Ma
tU1lh7S7J7hBqWybQIacHoBFaZG7vhVZ8ypQHY9JGqMHMgV5ayg+8qj/5ux0gfLYam9vF0IT8ve7
SnCzZ5S0zfWUxyMw6I0/8DHhtwbA8QZZl5/oCgt/YQdIipGKD9jdvpbc+cYADX8khOaaqi6ZjU7H
iMiGH9uZ06hYCVSDBpGui5F13k/epY+VXo9shvjg1qSmcxrYc8ZUJMsoleAGGrnMsyMVJWxXHlRn
AYbv2UJmIkt6p8lsEBkWP3r7CH8U4SdkPM0eTPOBNt7lqP9QARRAHsNr4EA7bdVybHv41QDSf3PG
lxi3AwB4HBRdsS2FpgQmo/DQ+ghwA+zp4teazSOzFwoSDX/ArViq1adys6BkwhQX4CZa7CniEdsF
TfhP5YYLpfJgWOoLAP+iQ8CINRsT4l7uBax41+ytkcgTwbmP23UAgF3DiSNX9nhKFiKa9qP02Gqm
jj/CEDaP2RLOuPoVoEvtHgJ2xtecXRhncTWDI+LJFRwE98KyFgIu4RJrlr2RYSXpGLlP4foCIW8l
6P3/MBW3epQEzF9tssfDV9PUEgsTgdhk50Wf7Gswm2G5vkxsK+PovLAsW8kCYoijQMnCYeQwAss0
rW+aQevSnKLiWE78ZzkvxX1a2bOhUxtXCuSrHMwtkuXSSaGX6Qh98XZTOoKvSiauf24r7MbQno5Q
K0n1hlRxZ5Ul8zobmv6n6W2W1PFwi9C9fLhOS73uWlwJ2wcn5F1QnPm88/76yxgMxqdwZETgH9xR
2BaiwresHf2euLbsD4xH8eNp+zWaWJGJY6nsOW9Gl/j7GmfGM0KuBv8nBmIkTKp8AWvKoZeONM65
IpoBXEKBg8lh7CIfwuc/3rNBgQKrECWsL7d98CgexZkclU5b1VqWO91G75gJFqBHSm36ZBQAXju5
oYd3fDeP6raPl30DpLHJVB/KPe9p3FqedHlkwWPcItSCXDY7g59sYUq9qbi9On3iVYI+yo9fXo6W
nfoFm4yt1yj5o2Mk2lR4leHaavbUvDQ+VdSm84JT1XWiPwcab1pDgmgAbkemkZBrG8AoZ7iBGqXI
GAfIqBDj8iU7syeEyFK5Q2W4PT4uYkklGc9qnYcIZwMHa9qLXUAROXYafkvXcvlO/vgYJwRoEjO0
xHehn3knm/vQyFLSf5HUrx8gjV1gsEFckc3gW0m7wHfzh0ntOGhZGBTvIeZ0IYH569PgIz7G4k4r
qwyfJADD16cTm3bbtC4KRBDWM21Cze03fqYvhkPKmJnk5jUdc9mAYCkc1+hewCkYhD7rkjpUXR8p
MHAESCUK9f7b3w6rajvWnISr+qxU/AXU8S6wwLdyBIY73yTVsDX0zIARzjv+XsybcRHjSrrhlYkX
kK9EPBBVGWJaNYQiKsuAKZ0roYTbRHp4iH/j7SJkLcaU9mVr+kh6S/pk85l9UuXBNsoe8v+f1BEn
Jn9CFxfSuy+a4X669itdohpMRb0dajRTX7kq9QviefN3DewF4R+BwsxC+DRbqrdvkxhg+Xn/pLaZ
sFpAUmek5ZCqEOy+95Fl3EjRuMQtHbFBUV2HTYhp9tYkj+L4jW/1jv03KAN25YxXWJbHamnWMdBq
j4xCuBr5xdMehhXDuVVE0dEzM8fZkCLDxvNTyBcnOI+HUk6f5+jSePaJOSxuESpNKziIPYkLLjA2
zlutZA6l8SumNiAWQ/Pmhou2sGNCMvJIMgRd62GA95/kmBM3TeNSA7hAcBW4KO6kBYnXfrlhF78t
nnVYpO6AuPFG4Rrid/buxDST//vmwDFhTpnNyqSlcz2dxZbTxHKfDsROusQRXh+TF6U7JyaOFNL4
py+emYh6BDJUZiy7o/5b4N3Mmq3yE4CVyoXorRDsY7SdvSJjnqeNCIazZACGfExs7AfmSJHGZVNv
dd6lQ9GCOno25Srg20nTd9qwelYQlVempFbpkQ9ETpX8Cx7J9VkMMKWBXgx9fO7gQzt3VwjdQoTR
OEwBmzvUYs/pNBCEivEYO9/Q6ztnDwfMf6iBEKKKTsqBEaStTvMCzgSW4Zko97QcJUjdWS+9ztyN
NwKbPUBkvvf2mL4hiiOHo8EGaTmncGrwAvaelhfLaaqNmDGcMjy0+gJFxVCbqLVMa5Ulk0ap6/I8
ivUCNyhpIfl78wGd8/kFLpV7/486dQw/AQy3hr9I4yTqunMeQkfX+IHXZ2Z3VjicdzdH/YgYiFlz
YPamucSM6/ofyVYREgIYSNuk0QDd24/j4ysvonEGtptjT+dn8zgdLsY9eoHtUZ0+ZZ+z7Z49MCVV
N8T3olP6WGHpQN/1UTXiCGomEXYooptz72Ys4+JTQkJTUrJsW2LA25e2qs6XtDI5ujYuVD1MVTF0
V/UbN3NQ6cTRuIwzCbBlYa0D6jlijNrPl/LBmVlUW7Gx+HBXhX/IXBIeMMgiHfBsP6LfFgryjlV0
WVEQ1gbDKgpzsawNenH06Ctq7qCLnT6PVBtCOwZ8VyDSCqUAMx4KYCyYFAhmg6+LS1yGrjB3cSQE
RSYFTvyErsuxC7DYn0etBbIx2R54vwuTNKoRb9Gn7v1csBaLSSxmuyIvuEK8q3EC5q8F+pYRXfNm
f3K7mb+W06P4VmTfSmgMsBrtvtE+HhVlKidtYT5SinfqL+PAbcnpyybq0NUA8ERCRUntKc0c4BNX
vD2PKW5MRygHcrDs1M4vtwxJ+MYL4iVxySPYKlqB9jPWD39vQmtJHnqgAavqB/RCTmMkM1TQvheK
ILIV6GKb2HS9rk7UGdX3+xiUspS7ZIa/vw5cfnuQZQgS07PB9M5q9b3K0N1/TMl4zs+v98/S0L+a
Lgt013PM8NbbJgcpy3zPfmepOOIF4baRqVhTL9Y90NBpy3rGFFgAQRPkr+tj+hGpIdtSwBvEcmNi
6KU0KtJ4piP1tWGKun01R66RDv3rfpyZLyFfk4JGSRjaOG2XpuSFGRKpvN91+vQndU1EKL/it05P
+/90+i4YFhKuTmOAE5qsP3B4lEjFLSKufp82v/Z6ddxaZT5Ee7Mv5FySP164FpoPJWvg97AfkpMd
lPZlhRAktjZqPnk1yY9kIUp66GNSXhMcRI5i8lkV39+aMP+KJKZoPHKC/4ZmU/CxxqDWFEtHcR0J
+5EimK6OlnKps+8ldAGrcJdA7UzWk8pwtFCqg0zCQ3Fg5RuuW4f5z6Gxd5Y316ob+iFvzoNdlJ2B
nposkOEj2uDPxbgct9c4MvuUl+jnEhFfcs/Fqx9KWQd3ljj27SgMdlhsQ7I0VT/QAF9bR9qqKLis
jOKOOCdBO8luvwWNIVZ89ag7oGfWJXcY/pKyVbfRB7ogdod+5+rU3v93vmetDOotRr1g9WwY2Gwp
J7CM+ipc68I4vr9UmfxQ0i/zDXbb417PAw/KQJClYO2vINRMalSGoMMhsECGdMFHs4UP618kfzLK
wnUBZQQzBdDhynE9Uazt5XskcqgtmwT4hXgGJc+XN/BjLXyzKmbjFkgSjRCU1BpKfSnwC6ycZ9Mq
tLN/UAPwg/pVPcRh+wvUqaN0+nZMa7+U40eOB3Uds/Fe3vHvnb/dM/p3Kdx6gYS9hH6yeoxWcIIw
yL0EHZNAEn0iGwwu4ALxUrBSRR23ShZRtAjiwBExvxtgZkCi7R2A6KHwSqrp7Q9S0iKR73Kv11eY
jITlWxC3tLK5Iec5PiHD8X9z5Hv00zwyCDkLlMv0j/ZKsCTnLvZFo9gb9jDgKUCqUo37SH1y9y8O
gLGs2nt9RWwXh8x4V3AZCYqNEZyE7iNlDH2cn8k0zscZ8YIvuj7krJcmGbpxU5ABv3H910q4a2LE
To0c8NUBpC7brlkvVSIx8hGls9VB6hupksW8xoDJZHHadmjN8ct5AYMWloJ8cw+xnQ7NEPSx0Gl4
wmCFYv9Ybmx70liA5FHrre4j7CC008cbKVX4tjCx0Xv1tGsKa7OszZJofsjr6uTq6+L/2mf7QFHm
xmw6z9RSy0rKdbckI5xXv1prn8HlPyiNJ27//T8mosE59sS9Ud6j85UfO4RsWZesU6lcZxUPJWNp
fAhYAPJ6ZnKEl6vhJvrOm/GoqmeBxftsknv2TzNtl4DxI6NWxMEeuMLhMpuwbldhkRR3NI4KCwS2
2ua3UFiLaY4HyYNbHQkku2OVkmQETBXUjx+XUaLgmqXfhtEXf8SSTWW/dCO0Cvxj9DaLPxi8u/n3
Oo4CrS2KwdDMJ3vrWkPE/AGGL6hza6/g6b73Pwr8XfzlFIi8cgCAZkht3ijEFH4n8C7uX+NNp8Oy
JbuFJ24QmJP3HMsOCartwMII5hMa6NT6zG376CxJ/oScOzdhthqqaJQW7reyo66KpMliw6f2Rqzc
wD5rsRJnacKMBKBOJboNJ34uPo9xPFbgulCJMxXprFUh/iEloO8sgcvNUBXLi/gwWYIq1tXBHrIo
TZB1wpriOCmQwj46ZojluHtVbPX8wMXB6q5E+saDCrdxhtX0wfVIG2rQ/Qi8XLgfi259gsT6NRqe
zVjuAAhpW6w5Uw3/DspsFiw1/4zKPybczCt6diqCWDaVwYn4rhTIzgAizXWCD0hNQbas8WdeMxcN
9sTyRdRMtfKI7hRnpK0dmJenhBSkTcSqoUuOd/UTvQhClYc/acnh/PMf0edsRiMYA1Bpj9yYMXZG
XtOJiXKN1CIwhVIUEhvzcu3LmnMZnpZL25SAyDFGBxw1x8LWEvo4zERbfbJ3vMsbGMq7fkkGi+Ge
szgcR8AvGry/mHNouiHVES++6KD4LiRy0Q68LNi4fNHklaR0QW5XUQrE/2FIY/aCaMRnpz256PqO
Jr3oOTGZQdunFf3+OUFy7gVAvmws/8xloTeVsrC+DcCMJulFp2/fQwaR4nK4nmtp8HL+3g2m+ozc
neWjEqG/46wpk6oQPBSJnBix6YodURDoTuaAnsCEb0OnerNI5PPOlWtSP0Kr/PXbXsrsgwygsFv0
PczWJ2oye648uvaTYvJZYAVCKfSBU3piNGz6DfMYbUeHbjR2EwkFOviEZNf3u+IftM8t9ZEZpmTP
/9w46x/dUuLGPo9Kq6PCd1ovY5fGSyr+0M52Wjv3PpEuRU7g7xe06lX+epRDmTh70Ci1VKQQh7vj
gpT7w+A7BJOvYEzWbtKmH4mEFnPPQYrJmMr8wzXS4ixnd3ioXV1QyBcly2DwHIWEazQ/5AD4U2db
IJerFynFfR/TjJoxL1s7CQOaguJXa6J7GcuS7yeCE3MdrFmJ4Cqp4z/5V85vIUvD0/o/0xu20dmx
K+o0CoQhzp2sEl5G70KFLTnd2mXA+95LRaMK96OqdXBaKxu/VXXe983weGYz/NJ2nbbqL//6fMAq
37cBPuOZPVo32if1qQe+HKN6oCnJl6dBX4Z0CCPvaYw8ALcq/MtkEcm4jc04cnn2Es9CX3P/p20d
ADV/jR7+rAbb0w5YUJXqy21p9a5XUmZn752YELoDt695anGb18+r4VFdE1FE2po1OtVwyb6I4ahX
o9CiErAx+rURzua/DCd/pyURuRk9t7vpzJ3OGsRKG4VWZNjQ/QWQPH0VLoQQLUKe2Q8kqjJ8eA0m
DxSoFQTLIbEYbllytaDC0Mb3SM+cAB00xlq+ZhxDinONog3A/miAxkgvLaXaI3RXr3msKeNkF48M
Qi6/sK2NwX+ZBveMdovbm3PUo80GA0iSuVQ6mW+QkNxYT7urF3yB6HYaylcEdN2pWMoGOGcp9vsU
ta2mpY+8eVyu7U5Sqv91mBNapQJwFZ0GvSuFPTTO3Wj2uIextcRlGftiVgpQEfMRNBBRsQomTRX0
KEh7ASt6BudwczbeguGeGZ6yY+51IXPRZdbx1hTVf1WKkpN4PRMn0MFWUYSev0Kb2PZjhlUcMzYd
ax9ze1wYEbqQ6HnhvkmomwZlYz+blPRhfMxQQgZRELsSra6R0r7G/qZ7RCCxc1FohZaP5vaR1uH7
odhGe6bwmbCfWWRZdMo0UyV2nKsDad78bDgQa88QZusnwhG03hjkHmEMNGDKuExTvHhnim2LvudU
Xb0WkevXKzRAZN7lVGnSihy1zeI3wW/l2vRNag6zIxX930RkRKQtujVxxpoGWztBYO5j7A2xIgCk
+Nyualq56LnAkiNW4brz68VzM32J4pfdNx/2BhgGaD/I2iX17uPbPxxkf02ZZvjCw1EWgIeEsEe7
B3wjxqJGwuohfPVyB6A7FwbwBKchb7NXKgW0SrB02O5IGqnKthK+aXcGUZXC5e0IhELMYefRFxcY
KpvIdWPlhnbDGd0o6Uoc/NTmV8LhdHJsrefRR3HjAPa5sU7PdUInfIIQbnWpcpD+Zjx4Zj14toZ8
IzAxAk5aLapZady53MeT9q5Y4Rm2cwdLk0i8IH7FuU/tjyYcQ4doVZPTlQWm+q24DaLUh5n41e8f
Raa0oe3V4kCrcAdzTYb3j8GYCa1C8AQyh+ydRl/qcwdmqr/n07rZfjX6OPFC4CjhnO2Z47CX5EEW
AwpTdiBMCMy9M1o4XrnJngNvn1t148kw1nqB9jDWxaApUWfyRlo9vqsIxMpkilva0xxDK3pk+cmk
gjj+lPKd7Q9V5BhS31YVRL3uWR/uH8+Z6vzNSm9wBrXPcM31W1BqbNQaTszxK6CVQVnvorp0G86h
sPJz5aobD0dXlxkcJErYBzbqY1BUsXtfjZSmtxW/3ZuCGrflRt09b3/Bojfrm/gyaZa1YngUqqLO
2xEAKyTzupr79QorKf6OSsDIa5PXtamxZ7W0bKyFFPNeUnVVxVsQtDOHUmN/kXO8DmYtjzpwzpaK
w+r62zvU2KSJ7ZrIm3+oBQabk81RJxHGsf9fFcQnrFBWOTzmGnmZB2NvoX6oo+R58AfZcCp+Z54Y
gMVEKGPAkCTJsdvAnGB4VzgsHMvSpjsL6mwtIAfEKGV/c/gIcSOL0REhBjyeu71IJzCVlVsjTF7x
PjeMrdtedkgaVci+H1ze/ux/Ef/9Zu4nfQ4ocqg9Bp7VAR1ooDRwTGpi7rNdCht83uxvbqoHkvqS
nBXWvRIAVDfQ+A/jE5NGOOQ/IPptvVQJqwmz8X1JSph59d/PE2mJsRk2AzW9Z5UelwHDWLiNHnkY
salR5uoeCFnTlR8xTpaw5va0AOZhL6IhfQbITcX+P78RMlhoFKCremy5DiVWh8clfAHXrioAicQL
gV340lUG4hPOaI3jyn07UUxZ1+H3hcQwG2MyVbbwDmHbqyCHUxUVqFgNRj/vQhnhNBDCn5iFgNjX
9QyRigLscYpN1alX8aU2ViTut+BIX23CY+BgE0KbmrNKK3qExbElFidzJJrEaJ7g0TAl/7okZZVh
JlJxmn56usgyowhJdZu26lnV8hq3A/7SUAeO39rCb9Xb7hIzO37TjmbXQyW5RLm0J+/1yKMKYkab
dNBw+MmhEtJuHEVO8DJSYBaMwzjqmsHVvbEigGAJecwaSd9J2/q9TeHWD2sW1EnyqyFFRaHGvKwh
71g0z/IjlC670Y0Wi8B6bkXRGOGA3Uo3500h3ebw3wfgOut9DKixW2L5pBk7CbpgTM8oPkdNWoBj
NdC7XVxvMxw/CJ50pl71YPKoaUr5rTgr0UvuWq+7KwowB5yPIWzvy+CtPJ+mXXU5S1C4GqxnPxjQ
jH4sl7hpQ38YNjo5UT+Hmee01eLuAxQs8rFL3vmkNVT7joi2X15PDb4nlJE4gSB/1QkWNqmM/9JY
IS+BlnkDqOBbRfd3yLpvwLnPUO16a8MGsPDr0q4pRtg8/zbcWQvwxEVzQgdR27AWZCdIZHAXhSoz
RNlEYRewutpKMnyAki4nbqWgeDY/PRvB4fzLUcZlVZkhizL38WbhnZX37SfJ2D4xqwh0wr8ilAhh
78oRPWW95bpRNhooJN/QxwWbPzLeAodQQvTMdeJ3h3TWNdE5oY43gikFcrrp7Ri2AUpUzQKciy9/
ImjBAtZJlREO4UXCSD4i2gt4tT84PdOC04SQBptVnCNYa8nkaWM2rURHAJyM0i54YtsDKLiscMjm
Zb3kfVXnBlFCK0vYsjC3Af/txcaqi/VWshuMr4oM4fM4uocwaIFjrMW2BDgvR1jVRPDudEJlhj8C
2Q/A0fEfRBBzGVisD0lCBm/yaMrt+GQzKwILqLDCDZfygZwWPeDQQvvOv5zFKG4LeuyvJICufqBy
wJ27dAa6e1L7izBLl3aF0NX0GfqpLD2v5IAP/niBxI8lHD1V1q0Cut132VRzoQjcTuBuMGWRFqZS
xvL6gahUnC0PEtGa+rVqf4GAQghnFHbL5JyfzxUYHErxta+snmpC0sXLEjwuScaEFPfpcLJw03C0
e+u5HRyvWwjGpY27vxW9VxWHmH98ZI2GkjEYJBWuoMMiFLIB9eXtxjy42cGRp9/qWYzoaSsKoR9W
NZ2zKwzRL7Ua2Pma+ekwxYpsiRjegUYjF6GRhHLYtRrRJCa0JdB9sBYcHi4gzDuH10N6wMgZB53k
nLeXM6lAi65xbQ7AeKqViA0WsHhHLzZQ0jX1QOlAFgiurmadVcKHMvviBYJy47Zw6JrppP8ljuEr
fg9bkqdRSRucUFHIqeawc3KzfTHazdsepHY375b2uxuPIJ2xCPTxtNQdL8BeWRXfTn7CZQgtLEll
u3wHQ9O0tipben9n3w0/Lv5YV/rWQP+SHYZ2n/Pha8fs35iiom9yzsIrfRimGrefddJ2tcRcTeLn
53G5Ck0m4L9EfWK+VuQ3F8R1y91EwUfTfGFvfhFf0raVaIgs5hpyoMt2PLFXk7cf6agsO4EfjvIn
84cHumSDTXtoj5pyM9QL/ciC1OU6vavHqpHVCCTaXVvJy7s9DtzqVBVuzka9Lj5FVlnkdIG3jGCu
WIbln9ttGwyXjNkZXefItBNlOEvbCYHOCMegtar5EGgDhyt+5eCxgMBgXaB3ayCvDy6UTXt9YN2i
HXhmxBmZvfgtOTgUUL6BdhnGF2cV6yUOWB3+Go24yn5d6tURePP7nd65LBRD1vWIu94V4CWJJbK5
51FYpkid17U487tSW9fQSdnjuQ/cLHVSiN1CYI7uoDGE7a2DDfnvBD3fAWuaHzEJFXB8xma8UXWn
hA+bUNBM4gfwTP9nU+L2nf6YEhFoBV2Sqp9vJjhsd9yw+MEvKN9G6Pkh1zzHw78S4tmS6L+/L5zf
sqfWGMhVZajhVr59Be2ZqvJPJ6o+9yTVdfshVHyTnpTbfiyPdvRws96R5/x152gmbtY0bvun05wl
J5AI15xBu2pMq323vGGDlb+QxXEGsDuWUI6OONxv9Jxpd9EMAse577OtBDxNy2AqaJRau4LWJpTG
xobd9u/PCaRdqiBJ7jo2Jz9ook4/Sg1Snxw7m01pp9Wg8Hvhjb/Hn3TZxuOlp2x8pui/prxsyPp2
1vpr5C0YxxzFwbs25UdIHVvxwm7T16YakL1RZSzp4l4p+C3FHDIMmRVM+ckK3FAlDa+6zEabpJHe
rxoD8azTTVhYTgHI802r8iphEB5WNA3shXiT2OKlGHDIAKpQ7llYiqtVo+Mcvf4le3k7f0Cnqb4N
OyHQrk6JVY6xy3qkWndkntDsK2gF33M9nw2UUtWRAQbvHetmb0W8+kLV86+XB0DMXyH0EYsoaxa1
KTMqXRZ2WSxJySzSFz/f2m1OB2XnRI3He3whjWlOEBC4Ozo+u8tx8ipbm43k50pyp1L17NLfTZ5K
nQuOiQxbmIsDV8dXDWS5OQfGKuy+RYx+FHlrNaNWu1smFS0sQB7olWp15sD4ZdUpboTD5oeZtJMp
IBd/qTDq/ym/CVlK8L9lbvfJ88W2hjKaGyDR7+e4edro7T5jYtGtU4osctJxRieDL//f1eBnBI1I
OM7YaHOxbNmqJAPJasbiYmdLNrmvs5Uho5EH2QL1pqsdCgYcZXbgzm8FoOy0s23dx1j7kMjIxwnj
L/8yKJjsmsY8zNuZ49PM2TaiCEH3yXYAYvHjbylOKSu+fUjF8xjE1aZA5Iun1q7XqwLXGny80sAy
ShK1ojr89Rq6xJPZq73C3g8A5AKd6kikc14qcOnKaB3KI3CSkrmS6u9mzpBOJoTWesVfF/G/Zw3n
KP/9SCLfTUsgU+Oj5frIjP6N2SkilAJ7EHxqJFKDiGshWWqWpFKKITX9mKO1ODLrOQbdNGu8WH6i
meAf8js7MMDN0ZeWULFg61wPK9JgzrbudafTrmZnzwQOSKzMw4b3ryoPptJTn54OB3WkPXypMfCs
RMrd9YJZTt4+6J5slC3UefRbe9SM8CKiqmx0wH5/mmk9uR/eCdqi+zoQL5H6ENhlOQk3ajRIvbcN
dAFlWOgmRvxmLvTrPtYu+xSnDy6t0wjlI8rfCKBANWGlNGDoUZoJO99OmzkPOa3FqrbbQFZwECMr
ebnZdb/FQpenlvBy5lPkEymb5p1dbiGaTG0IZUK+CeDGX/r53njaSrVHGO3tmEGq0CokZyyWxrCE
6mwKkGRYjbl6mEe5Cp+9mPgpqO3cQqq1HsH33moZU5TCN5BVppezHeB5Z2M1PAfinYoA7y4dWuMw
88d0FjO4CYSo7qdWKHrxWbizw1RAjb3S6Q+TWzlpG5qnY6ihdXAvjNq4xCm0Jagz9O1WRC1zavYW
ezMyXRXSrtowrGHgcU+ogVD+Q70phKHDohJHlBpD9WLD3zV/VspwW64DkaM5lJWCUaeAgAb25eIN
PHVczo4TIomcrR+Ul5ChWFjz9wN9uENsZIqX2lAIdBl3mS8Q20VJmCPe9SNC/tWKnFK4bunqjHvf
YomjqZ4oQ4m3iYO4X+NngryUs7844s/p2XwjrJgxFZL1rJGbVDRQxqjn1TJx6elOv3LBVR4BysuM
feQhWtlYrGxueoqpQPde+XsShRGs+KosuShug8IZtnf6vvshhEjxp3Py5W/W5c6qnNpluie4Iatp
AijY2IICPEm+6zTX2vEELWLj8FP+N3zdKV2utAGKrvoL606eWvfhJvK5XQftZYxMlNqpPJmRUlho
ipZVRSfZqw3YVShVf1/6xGHujESdDXRYqbgJL7Ntx6WiBgfxuTKQ5Jb7cKInSj8jWWz2PJ7s7dbu
tKgrIOfEmsbqFdl6Vu8rqu/qseeHvtfN0svGBCdjquOVq2jvVPGOifRQ6qvcVx2oEZv67PKf3EF6
L/uCnYLT+VWykh5W7T2vOgwx9aaqf7r51LIkeRi+ACVVdfnw4vktywSIJmVeKl9teDEVMhP1bPdO
q5L6TK2g2/Fim02CD/UgHOYOv+PKqfoTy6eKc69Mp0TWFaZLYcNRi+nkTbeWlO+5wUOQkwX7HfKF
2h27upt5rMH2qTWbRT8895CZKACVf0wsJdEmEelCynbRuOGAe1gvR2Fwx3FSA+wM99ogytCJRmK+
bJRx9WDb9zh5KOfknJo2Ysos/UmXRvJ62ybBRwbVzkZVh9JgUNBpbGhwgJJoqte21q7yhDd/zveq
e5CT8wxQzhYvYAiyJS1LJQXPAEul3u25kQAGveCJn59HRUMTN0jwza4SMYrx4zMjW+AD3SWxOqcw
ru2LryLkH1F04X8Ub+ImaIug4a3Oqjp0fiiK3XjXQyxE/CKqrMDtUrYHqT95CuT/HA2Eq7d2C2qy
0tymHpZvzz4vUaBsBPHLNDzUaueIVkn9II8k5piHnFqgindNC4AfqunLJDzt68NWiNu+s3NkPJI9
ihp/w54n5M/y2hAfACJHxJZwAEql61yUtOVjut0RGaJkptlrFVqAljYIqs8cK2+k8mzF4Ep1SYpa
Y/Ytdpaoehzndh30NouptnLiojh2el7xPNKtx7S9tWcFSoRP2hSkF242xmgtdU8z+FS3pbJ5EI1b
zTHxNXcJlXC9todvjOa/a0OQpFA535KQDrBalHQ6y0aOCrCquzb76ZkmqeK9QkAuP2gTEDw8beqN
Jxt3S6FJca0rUmzLoi/1SDGkockG6nWUSycFhXCMOP+nIBXBIChuUYVAm8LJ30MqDC0mwxNbytmn
u9wGkJSr0VR5qwBAmInlpljLmLStN+TlTeoKWaF2dRHrQQjBCumxdQwWyjlYhzaavq6KKwwQ3c5O
NkZuWUhjhbwRYdZPg2PwirslANgS+01QgHlzgtYNNkGxZ2JbHgtTMHiV2EqGac3Nti8iWpTvUZzi
oYxaPNAWy/v9AjM6EyVd4b0sllh4sVv/Q2WhzxOqXatJCANRXvRqXK7RaDdg1MeFKDF5Uo3euLIc
vfuitldF9vX5rY0aVm2zzs688G974TP6O87fNtLBZqpkJ823VwPkZ6Y6iKLFh7GHxpAxpvoZSXII
CKRmNe2m44FTsBNvlebDUkutyUBorvi4zsb1/4g0DZEe2Enmnzu0lOi30uGPBw3ylzFQQ9rNl5Xu
KzfO2au6emU3ngQnYUhL5+IMe5VkupOQxdBMuxGgTR0swdqup8K/02psoBXtrNGdGypxT0KP6/xR
w+DMw7S71GskXZiDmGVObEZPmV4MSx1+TzH9I6wUjUc/V6Q2BjtL/ZxcJgl4UqrPC+XfYj7vpIyv
ePcpXcYiSdvDWJsAMSU1Kp9g3KuGyhN5bcud9JMuo+4IB83rGFnNQrVqSwHsL7dF7TlGv19SxuWj
5o2K0HoaiGznkrWH5CtwYOewD2BBIddggF0pANQAhJBk5qn0BSJb9z5IaOrQx2hnB1X17+5ojaOd
bRSpjQR0vS/OMqLDxEGEZ0FwtmVPd/v6gVsUaiD07Jftd5HoT63lfplCJcxnakP9jy3R+MNZ6aVW
m1GkGdhrKbY25XU7oZu99Uq8aX8KMAFBOyXdqeP+WJVX0+isPB1yE8FFM4/HlUSxesULwDanVyZB
FPxYl3Z1ItNP70FFEh4NBbP+VOXMQWY8/UwzTGw9Gjhfqe+2J0AOJ+shi/+e4i4h7Uo/lfgV3tw6
tkDLVrsGNt3JVazxEZyHNCmDP3aJsKU29BydG1RMrnPh6kc2ttAJgNnaRAh4+rHodtVVoO3TJRxg
OFM8XgxmQY8CPCWGpWuIeANlIFLx/okv54m3noGWHoHIT/I0f/5BtrJI2YFqOCbFlMnKqsfFVLya
nIm4Ln6oYCVRotDte86+Ukq6YrPIyxlW1SJ3crt259M7AteDy8u2jNy9aMxpkSTNEo95PVuxU0A8
o8yT5TrWgj0sDXOG6AQ3eEA6dV+GVjVlNfnf432C3JvEJbqlPCeD7VxdTnvzsYhdZflfyM7g6Q5k
iCx/WNdEcuD/2Imh1azX9LvSxRQyh6F+kum5ofKzOSt460RlVmFkxkLz58YODNUUZoz8dwXGK9w4
eSA0klLKSa14JZOGYw3XTu/e5eAHH7zDJUDHB0saFFtdHbKQb48Cna7lS1cHvA4UWk4OBENDww0U
2hllRTnyiyM4zA2b2q03g8wOr0ddR0bilx3LVpKhO8TpZIWhWEuCY2AM8gf1HNOj8a7kuxE+/vCy
dt7rTUoURkmM2gycwb1XH1RtzUsB9mqzRNO9Tkz69CAfScu1iprdQPOJ3X1OrwMT3bb93IcmYMXg
Isv5BkX8AMs9TOh6zzMmnbIgTPAATTk13wWjR6fWvbks3QTLczC/Ccqq+0ZPe/C9Ty/6klKTEXD6
h4N1h2CVv2b5PJuUZWpvIQXLJx4TzVrKBK6VciIl9809AEm14MLIv713NMN1JGNas8FEmSBhyIL/
BrdRBdU/Vjk1NqYbUcqGJoi+D0iB/lEmue0d6zBO41U6X1W73JWGweh5/hBXXVVuukNIsyWwJ7KX
ZPk72T3+rQWj3lOo+HEd7l5VQAIwcSXvXSJHdO75zbxSPiY1nhfMp1nvDHtOVb5vNfZjtdgSgOiH
jnD3XapyHlQp99+e6O5w0qLe6REdmFaAynIBPVybX8dFcC0Nrf8LDWan9Za6nvzR7pXzCzKC26hn
zXhlibb4VMtjFmQCBykph9xBQNdLS8HhS5c3EUEj7129l92lXrzj09F7xd5u0VXBKNfFH4Tryjeo
gOX2iOOz/6WYmmNxNDhv8qtNZXAyXHFrB/ZFCfqoCCosPkEQbYj2TkN7WXvwP4D+ya0hoX4TRTBC
5QeBLSWXAD4uXZ+7cES9Kk57s5FoSbPgJ/T++5D/4hs0Nog/6FtUHbkrYo17jfEMD3DGNB/FhabV
4JXwVcOkCZVTQPOCibrHmjwh/wP9P1SKXaepVDAhkjBNjblfhhHxy0i+plbN29hUNzXjbKhCPJBQ
+8D2ceFBTL9b6TJEg8gleNr8ld6EJj2muBL+oqHUHsHMZdkMs8NqiQVYkM3k3gP+7WFeARlMEwD8
pcXy9hmc+EtUbUdmzQUVI9QNtK9if39q6CT3eEIgWw6xeUF8AjoKI5lN9SoVmwVZ/Ouy0lXAq/PS
TrLsb2/NKSxvpqLu307vi+nTuaEHEXxsEizpz+MzaisGwM8+FckPOgxybeuGz3SYnytgXnZYqwF+
l1rxOF5FLoc/qPqcx7dDFFANwucT0x6w+ah5mTqtqVrp+u6vntkie30+sVZqQaR7+JLvRa42U9mi
ImF4TgLbf237oMBYkBGKEstc4CKf6TKw5xkfoUDd+aoT6k5fDuxK+9HEKGagO6StmkI2Zbh4tFq/
k/8z/007ZNf1wJ/Use9UNRyurFP1XuMzf8rJKR/A+JPXFVmY6rzvj58uuCM8ykCoO33A9i5/rxCl
p4k/at4x/2Jkf1y+SCZppElboPxGFS6CceEbv3p1gC1ahgc9WM5+QYbBMlLyaGQRzbOrWeFAVB3e
7iLFq+sH+RHvjExxmcI6SuqRuF4xigSqQQlXE9vCiXP7N4qtiAc80gT/7shDOKGU1rgkttsRSybl
ww27MJcoTis5vc0RJVd2TZ3LTe7iEzGq2AFGwO6okmnrRHWHr/prw/qKPnfxFJ0Vs9Alnb0FPDRH
4CxgQKHvYpFAev3OKGRhVBTEMDHUAnmJlP9QuLLM4sn+fW3TvTP1NSWl3MGo6ZrWC9d1Wwho6qd9
4BN6YbFDOrS4AbH/Tv3FQbtFa+R6Y0tiIVUTqjAb1dwkeOrx/o4dmyfxnXnFjjWeubsy30IHilU+
B7+gTKcncn8CxKmHjU+ezioCgHXDbpEzEVtyqVvL1GarZOmqjfK33Cr+lOq6pFYuaF2wKxHF0ALL
WEfRlRAsFqyLP2aIm4n3FiGmyrMuHXQrfWNkVJHvmYQlPjk4r7AtMRlH6M1BJeJnwDsQGyZviXyD
x9d6nwVPXYoS49tlhmSgx7mfMt8PsOjXzzS+N03/y4FRk9ZQ9iqaYy2JhChqn1/VJKhQKNDhdhnK
1ytMwGAunfCZIixnLfO54b0zLvajHHPyMXvtE81ePii8cmiAUW/w6tZIVEkeeSK2AqMvcp0WMIlF
P0+Ka9IJblKigw/iJxZXrE8dmu1gocAGTTAQD3vhef5glmAjhiCZ+4syt/634tQBqlIsTdsmKaC4
n607cAHxXG40jh0XCZTP8P3v8answFJIeVXCPFcQAp+uZ/Cyrcs0vpR/er7UqSgXoMqw1Uwb35F/
hbmoMp3/U9eQ1xX3+6aFGjMTS3D5wnhGl1dkuMZpoNS2C8AZf+yGr7/eYS3rGN6IP5u8REwfJn66
pEx5pnK839O7AC9lyqd5/c+pfMiQgXfUiMZlh6KlNGsJmkBkAJLS59rLdIryNm32NX/3z8Cz5iz+
103h9Ds0pvhvom/qNxdxLK6Ia8vQhOpjVLDqgENr7lqbEvT6fMR6xO8Zv4PLYGFIIgpdCMoqCL+f
+m/v2lS8YNoWuLHgFVgeWmqKytMtMy+ukl9zU5j0qe2TEbDHeYhY/19A+V6IfEixt+QrUmESyKaM
2sfclc7bUW04PtPacbdvRlwhY6KKVJlzkcFdIuHS6uLYJWolEPsQHUNr7CaEnA8jUYNz8/+4N3at
YHYrQn08WwBWlwo+35JmGK/bs4CIQ/iIMpWxGAnad2MH9baUizR0dx5gl1EJaLxQA4xJOT77ZiGZ
PvWFaaSAueTSoO0nxVjlYLxe39AqcmtqWVhygKQr5fYRqD/aweSQoxLrVkfa+lCYleFh4DIUuJWF
t4IG3tcmDWdEXmEMXjHTZgToONZA15LxJ3frkvfhDsyb0aib2Oq/WfVCBQy41IB5JftMgdkaSmlL
nDzRIEkH40g3TqTEq2Ps3J7H+u79IPTZybCVhc8Cdm5rvHxnvuo8FQ9BqFdUgMuEAfuYTrUmzkNR
QPR2YBRHXo6Cknvr+E3ol/stjseRfLa4ACEG6QXjq8v2M3X9Os/51TmDuEw0sKbPbkgYwj1HIIsH
7nmR+QNxdHHj8KraYlGW0Ltg/LoYG1jhetU5pT4n/P9FSEj8o0bvdfDw1zXTIH+Z57tPWZc0mfPh
CdPeVwnC6gakut2iKBm+Q6saGYORb2qI3Cff2KmKHJBrC0SOAA2GlXF+aMandwpUfu/g0KJSn0P6
EHhKppvyLwiIZWhWgEJalntlDSQEoaqucIB7rn4gDYBzxlD8w3RuU09r6a3ojtyQ/kuWw3deBOFk
GntnnH0kODO4anAzPeu4cyDgW67h7gg++SKMW0t/LUEj01a9tMK52nZTBZw5VOWe/1VybrIszHvv
j81kX1CliLvNde6vA0BAaZZnvpYt8mrWiLwB2coVcdDSzduT4YBk3pm31TpifqYPK2xVaFnVkJUn
p11cynll6zqvtJSNLzItBwbYhPWirigLQktrX5E8hq7UtSan38eF8swjkjUuLpxpLqcG4zP3r4iT
g0KyuZWkjt18saO++RcLEknzgne7O9N93aPYv2h8bu5m15YH/6I/A2XiLwgVdMhRwrnz5BUNnIT1
Ro05XcD1eQVek2YUx7xYBwWdDhdff1X1KVaiOLf0qqmykM5vujeN3QXyK/s1QINhxeQ003qkm3dS
PS+1DoXDCswaQIOpq9HmeWyL7x6bfWT5BVmh9N1Sx2DThC0snyP64m/jHejDeSVXyh+gyzRN7NdQ
zpa/ZPQo4bUiHsvP60CfO5+QUTHjvrwZbFMcxEN1ixVaT0ytor723605X18qLb8QCS+pqR3WJBmF
5VcDElNDQA0IGwqDQ2i7cUrGmG6W2ZAxUwgspD8B2DlcX0YvDs1rYEU8Id5Lkp/BYrml6tnjm3ut
7Kx7w6t0oky7K4RCcB0adFzEOUyIvqGf3hBb+lhMrFEk1CpApotau89hBJT54djHHAhVJlVGAG2B
5hQ/W7Qsg89DWTErQWVBRTNqI2XG/4nilf4jx0Urlxc5sD4xRfums3ZrXOJrZqIFyvr2bDF5z/kD
uJoG1Nf7mLXolbmGWEMS6K6Tp9ZAEh7QW6y0ODux9yXuSpYhTzZ5+pEOUqh0kzPJDsAIgGucI6cN
MSaUWS4hQheuy+oyTgL8/z7GII55TmO92ReiuUtE6Tv4RSj79XxCqw8vYuuey6WPKmGjWrm+Ir2i
mPvU734vQR4OtMTHT62Q76Iy07MQXkqaDQzAKVok11mqpvAB9grID25k/bg4QHq4aVWLnNZ7x7so
vpglUCHKLjiheUsefYwbBh4FZOYWelboSaKPwgHkV23VsIlJiWKVCQjcSCmZXpIYyxxm8Yz9FXW3
a3FHaQZ5eqsByTzC11XKbpIT1Xgj4YvO0yjhc8SXYQ3SI6AjloxVBXB4IlnHizQvV0KvrnQBqrJU
dorc4Sbur5D3a50We5Owk3K2YPfMar/9yvnY2WhM9tjwWfLPYSEjg8VfLDXbeR+g8rxUS7rDtI9o
G8EIXfaAKh8UPWPWzkUWWtI4fQc+HJfcn9aYRJqQnKagdIRnE2nCIP+H0Mn3zBtf9l2x4zfB1mq2
8+3vNvWAw3ru7zrw8n8dqAoGpxEU4VJGzWsm7j8LXXvhr2dlm+CJuINtMV6yJ2qTaxYlxokiLPxZ
VPvwo58UqU+ZQH7QUVBgpbpmhaD/pbFXBRG8juLoat0jA3+Aun7bg5hxVuXAp1VmUkmjAAqGcaUd
o31Vtoofh3UQAnAys529beHv/rTOY4+6IwW0oIT12D2Xt8LFGDJxDxqKtELKuUyggjiWhhR1miku
Q2BC4eDLhzhlqtAjGE6jG8vMQPF1k4K6twqnuZagpruYe5sMlODquTUPxHA2pdJtTAE9InLJ8r3r
wRRv/SoW+9VAGl3fAVZj1kdHPlXsUPsHklXpzs0qPhcGDI5H3OhlCiTW4rBSGWqSOjaMDDwsAzGQ
66tj/jL6pvRR7mEfXNtXYHumLNip+fvD2BSlHfBTG0r4q53LXrYCc+yz24RbB6K42PQRXJnvD9Uo
phwgABJAodkxGRa2vPNsnQJtAR26HTN1W2CL2t2f8UxohIXwRRoLsf9EcNKhp3DoJAlqbh0aJ9Jk
Zp5m19YldrdH4KCqN8Ub8GuGyTSVUfJLX4vA+TVLpSdmqJYZztkGmBwXl3D0ifzJrgmhh/OE8vnh
V4xaX8fy+bZ8rhBqiQAP0YNtxDUuPrrw1Lp9ESSD/WYUKvFdqQenY9w7lHU2hs1eiJQ8MJly77QS
E3y7z8XL4ikcNm2dn8kMXuhrrF3bWpr2XaJ+0Md5EShXH05c3DoP60mWtMVMcKzvZiIEcXZjr8gq
9SXk9J1HeUk0v7QUWGnzJxSotfOfds2tl/x0GOVcfPD7Z4qpivO2Zyp6TVD/OV6soNBrEf/lom1F
u5anBb0YLSsFU6NSFzIDkfv9BKcHkAn145/1kRUahLC1Y7UMajEyEkbZDfoktsbPOoyTNvTQfNq5
SsULLarvCU+IpFaNaZLLsHl5ehctbUtbVkkiNW/2HnxFWX5evKKQp73awxZjnAdcoHY4n2hi9HsV
YT+F5MG0nyrobjHPlLev6Y26gQJHPExdRb6vAoyrWEPjkE+ZnLAw90AyaCw86B3SmyqNUtLh7mve
qhCzYaHHHTRPAm7khOdrM5FTA110U1VEDiBaEMKDlzqJIkkEqDk+NCSJC6esYSMmfPg2HhpZzjSz
uQc3V/Uxnsjf3w1n0ihpVP5Fa7R52F8whHHWYCmRr7cfFJLuWf5ar54mF0C1kyk/n4w2YL1QQzh/
ipTHqsHMWzQn/M/cN973cIx1G6hiNUs+a2yT5FAu5ITbxeRkOSsazoBIosN+SmhTjOfgmmjpswYu
3Fv/hwRnWvCOZ5z9nlvyp/O9gxuQlpK7dEZ+5UZuTvV8Kcwu5CTi42umWDxFO1fgJa98R1uIExs4
hjsvYQaZ5m4WGDPMZxlz0H9vNZm+ww/u5KUJaxxfY8pXNOxae4XWv82dwPVTlut0c4KuYiXD7GTA
5b/PXuTNvfQ9pPjc66bgbhgYWA2SvS0TWbWiHhVUV3KD1E417Iczt3L8/7hoVH7l5lrGPMlMopZR
Nu1+Psj6EZ1W9ZQ3Xx/46RMz8GEDVZV+slX982AaKvaIhMuPNl5HH4pTR82rc7dVNkImtA0FU2lF
/pKGnhzU0ROvjYEMb8rdrNNMI9woAoUgB2MGqEd6HPJZY5EJgyH+rWd7a/tryxUAT0hindRXj/hZ
BGa7L6QeCD5pQXmpAjSoaJQt3sFIsWFSL91BYl3j6b/Z0lylcEECSnM5LQEmLWjrFoDQqCn9NBbZ
OdUAIa7nI5ijynxVsLosIP4qv1SRbod8vjz6PxY3Zbn9ZzdtYqOY8iaUvtKfx0wQRNMkZJhoOa6x
gxv/xrD5Uyt0Qdm69LhUbSBBMoGu9Y94TCfXPQ/kRJtAI+zQlDjcUHWMyauUaCxlFiTbDK/4VMbI
AW+AUjSSRNAkaiCjzVBweg5VL3CEYuFLoUqXv+Gjof+8lYCJWTkoppIkhuXnFqu+GCN84MvbCzbe
i43RzBH2XqRNIKffKsYKghukKlOwldnN9UUqL8vhB2QDVsSvGEfpJb4fzgy4gI/3SHukdTFjLQHC
aybShxZc1XZikt/v9gq8mwxRLoPcIvh67RBIKhiAF8plP3Ob5oQrSidH5aduKr4mMkdFnpm8za0V
sY7mNbh+L2vVJx7BmljFqdsPSqFiWWJj1a4M8fJsDV6eROl9E/a06G2mcJ983GIHEw4q6X11OLeB
jwZgt1ODaKmHE2bfRdMOOw7Cdqq8PTl+s4y+gETihUTI+IX/DhuRzkCev84d027qj1S2Pn5HPNQI
r/BF2nMjTf8FU8GXcm6kP3ajoVPn3FkJ5WIaXV66yTw8Lgm7e2L6bHj5v3/gKPktAOVDMp/aMQDn
HR6x5BKtI2MbvK4DEILttT0f+33zMHhqb1Gk+9200zfweTn48bmB9xHec5GyQsLTMQ2v47KYB127
uVQnJQHx4xHgtIgt0UVyYKRVjn9bXzWRQ9YzjelBOtkV3OVVL6Dem0lZNBksYJqNgzeAoCy+S0/5
CLyxKFqljPimAE1OW4MIFO3UCuAv+moQn/WCsx6xUSWzVjpL0ups+UvYnhpTSEX+NbAxA4g1250G
NRYzeFy0GaY5ZxGXbnCqhgbBJbJBL/PNNUiBtEEPS/GXxmtfMUVMXVM6n80wEVYuPcBU8G+y4gYR
/Qpg7QA/YD90mIWgojBSDLb/sverRhzMUGlmR/XRf/jsLvg2/+4MM2P3arHGyjDpc9zE9YW5c5yQ
8HqPwDd2VRE7Tn9380LInGooW7ktwIEhmWYUYmZM8vPSjQJ14/I7SpT3JmE2qtxyeYgyztiGcIMk
3inDxJlVzBujI4AvroqPk90GBXjl3UMtZ4N4/d4eIPjqG0LvRqsbGSHwPJHmIyvp1bcD3K9rezz2
OUQvG954yEQHpGh/Pp2C5SCcW+dZLvhmgNyV7Itj7KUPd0uXX8hg3YRppNkBGyjGzqCJY7M5a1BR
0hSFoRJpsm+EaQ/o4Ma4BM03RBvPTqZDSrh2/zMG0K8sO8olmmzax5phjkx9FyaA51dVG2Lym15u
ODCmN3zKzxOgoA4LA5M7YYQTZ9+LbcySKBqg26ZFDCgpXghDZXJVmmmbPU1DjYXSP+pQJhC2YvQf
uuue2LGieC/RENGIXP/nKDMRJLcC31PIiU/XiXMctkaFI162v53D5ksWRcnykCKpYPsVt+NPNdfX
z0QQEN03Bbs0wYfvq5hbxEEEE6XrTLfhSSs8iw+CGfr5gOURBIaDdIOrOxCfwshUKTrhhVYnt3iR
7zGrIg4KJ2S9XrtAZFljPd9jRwJTjJk9dYJYr4LUyy4+wSkgYTxwHFaYlOn3CDdB/ydwdgTodhZs
vj1ATSCSXr/sv+1ULsGTRgX2+qnWoQ2OZAi/fx+9p84hPo6Tn6Y5PA9sgXdEM8fwjSy2s1+ZTLM0
5v0lYOeCqCjSuCwfhhmyACzGyLudy42PXU4xJGT0IaNk+i9FTroh56gOGN4Nd3Dmznn4mUV5Irl2
ajjHY4Zql4UIfx4bPV4bBmqNh4xMzRU6DAXXjdC4bTjsyDzvR9sYza/D7s7am5J2xUdxK7bZHlGC
ZjH292mCaHo+cB5bXMfOSyF0VOFDxN6pr40kWFfUuJ47zZndSvskL+hWwnwbnMzYmWvG4rE7/+yZ
QhG3mm6flc7okp1Zx+H2ebX22mpVghb34+MDcTSsnxiSMglOJqZW8JdTjBi+DkYLfhE/qY84kQGH
G37u5Ua3rWlDf3X9ZvLiCguYxe/qUxq8WuzyzGVugYICXc4Tx5aabct+LFEt+L90lJRLiigYhLbR
gVo5+qs8YtrdJe0T9wr3cox93aavTksISzQHa3f/G9unXbmYn0KRVTMT8bJCiY0dvavPzV8RvK5J
fSsIoy9LwuiAUo7U4hSieh4IbbCWM9ByyqXS3tpSCx4Mu1qUpKlnACUvTj2K5JDWH0Hdh9eBrJbG
l7yuMWE71N3+E0DQH4ueqtKkUy8kkw2xrjp8r0HnAk3g+Je96194PfU3OHYNSId21gfyx+qh4hAH
yt1INEA/R15SLWSnYqDQ6UmIgXUtcOwY8wj3ZEzANesGmVclcURQj+5lAzL2me0o7hrDCBO5jlIO
/VV1+Wka5bQTuGdYpN80EHw9Rzl1CVOBdQBh0YRInVMOUYYLvXfrfHPc4KvosEPFbaXfB8eyTrsZ
DnuOlda9ujb6X9sbCZM+tQm8UHtNgGQgenH1w40heKvp9E/U49Kv2bEaqoJwHwxIOwd53gfcQ1QI
Gm3UG/2xQVJA80SneJ/rnZcPed3cdZSkb9QTpAuLRwuZPGHaLDiZ4ETklLmBL6KhjeawHYc47gXu
PsAEMuaq4dga40Rryli2U19lrBcKucHyLYYIuliRb6pcdFKQw9B95RXCKkApMS/ZwIvUI/XZmaKU
18RLbbs3rCrUPi+FpIoLs6VbK8gtr9ziQyTikeTGGIiaFS13FKkTdnkR6WW1O8MIkEg8oMIT+UeY
RKlhmk2oLD54UqH+qUkxCdUIS78xZjDGDVq3/kO/KaZ9Ey6b7oq6KRtSP4w0yac+RtYzMFFyC0ws
LRE3+ItuTAiso5LIqDq/10beom0+kGTMm7rBrCOjN4qoPW2NgFtsuLTe7xBjlCZSH9N7o0fXTH7h
MThnTID/JBqMfZ8qYzCBn/l1D9LcqtPTOiiJouH1nFVZDJ728KqYak905XIjzcKJeAZQwEhEoc2G
lCswqIeHSVmEsy85Wx22gQAq1LL9SRERzdSpQqy3X2ItXtuCrjP9K15UoOfjdKyvdGytvRRtAQrT
IC6mGnhkaLf/67z7q3QMh7e/nrtFlk4QTyO60fgdm8EREK4Iv5Urw5QCRtrRF042l29jYGW5MA7s
MqM+iliVHz7zVn6DWlSsPT3Yr4oPI5hyACNMJdd/TwRUoqJBn7Co5w78aP3ZRl5aTZ9so6paTBql
62aATYLbCNpLjONF7fQM5Ippjnxo5y9002vNI9X4kCVwB13zwj6JI7leAgZiyuCjbz/cB8wRC7L/
/Y4xLlppLBLUyN1TWo2TN4z6AtwO4cTiLaRmQXdxJylLeg5cy1X2hOtHpt+pNAqyiKXOVANHzAXt
3g0eO9l+vOSzHTX4r/+DUwz/Mcemx2dKT5/WDrRMhnJXQTs+rjNYFdRthd/zjgFLMlbMB3A0sCYd
W/e4+aqONBPw5+vtglGu2JUv4wsj1bi8pV7jv8yjLDzAy7i5hyERbo0SHNrt2InnNWIIQ+aeGDbN
QxOHOdLOtsjiuK1/CxnN46kRU5heHKyt/JZ0PpCy5J+Av+go3gxDpru9GvxOHdgXmkugjRDlfFPu
d0YpQe1gjbWtTXhDuFliibTUqVDblx0LEhG7QsSEsxY3DbSpfqgf6cF11TBLz6dhnVKTSMmTSrWk
5Gr00p0wjlMEgSX4CdDNlXyzjZreKnOYNpDTdqr5mc23JvS+w42KEcom8qawPaaATPbatvpZ6JYJ
OMFKc1PII0Hl8EBE0DmyUSEBhdffPo2NtS/e8RJsM2tjeo8MWATjA/aBVG49es80g51yDkt68fCm
HdWDil3il8KJHtshmrRgAZpnL4YGpKrfXEUnq+ynO6lvTs0ti549/Z1xcOdFWHELH1uLmEv87tc8
I1TNohJHGB9rdee8LHvo1N4rG3cn4OQYFrxLosrSttx/fWcX70t4KL9FdIZLcRhi+8r1fubcjeCx
2HioI2w3EIRdFwLNW/D2+nCGAwu+8h64+mBAa7bZ/tUAEt2Ko/+Xup2YLRD5zDr6bru86dywxJqq
cHFZj5Z5DZtoZsf81RKVWNrdm3z1Uc72m+/2O4d7eJa2sVzzrTE6j5f8MaG4dRtNJBrQlcqVis+8
6vL/sN9X5nz3SAR3Hlh7lPgsS7fxbTcTqSch7JLeOMds7UYT3ZtACe6copn7J2KUIg1dMvYa4lvs
LD9FvFuZhfALBprxpEM5iyZUeLvOMPz3lPVXtCNDy7NmhRDvcArfPzAXMupHv37WFZC/Tvo1XZBL
iXDJcooowEp4hzgE+okRLP9+YMKgLMU5VlbdLAQl44KL7sSxwJi23yLjXGJYW3mEhT6il77A9D4m
a55kz7dJ05lg75OjT7C8afuTXXGuf5T3RCm/E6CvUmnKPJEdVuioVKeqZtY/J80MA+R9Cr9+ab3U
+j9elH59Y/MkLHBJG0yNWXYQazNNNzx12WytJqHOafAOqTYcWbjgRGaAe+8c5lAL1V3rdQheylAo
P9GG8vqQEPAHI5j8V2Hh5XnfwlN95q90tn1N4sYPuZymJfHNZIPTu3XtiDf5yZqHoRl5R3q8UJY5
og6CW+NEDtLPzMiHpGMN7p74LkHlLAmbAp2M+Ig32ERk/aZ450TrDmis1kOJLzoAZjALKAqAnSnn
kbK135oKb1tUqomeFgtu3rhKvQuufvGjEBiOXd1BLDxOo8zv7GnuxHZwpoda3uOIuaLpD7MJdRHF
cnBS3FXarsGrKEBfrDgWCBMjK8+drAhMt+O0Wm7BoBV6kZC92a+KG2qN+PpekO/hzLyO/OaXwK05
DIguyEuUPkfCLxhlNvVZYMxh+BhFXpzMcwYeVGUP5GmXX4jUurxBE6FtF7Tnngp1OtDPDIXsgis0
UokF5NVsxrm/N9ABsES/axXlWB/1XqTOYXtAAFnwClBoHwBUfIv2vXosue1rSUMqk6/3UbOO5ci2
HW/M7+pqo8C0/fPYOD+qM45708lHOl694oTUSph/O+RStmhUKTUSc6xgE5Mh+8FuUXDc1BMEH6d0
XQ/EaI3Pmio1l0okjUW2wzEU4bt9Kuvj+2DNavBIRxUK4memkiQsukLPzfmrgYrXeyxHul7fqUq5
RCmiuHDNFj07Pcmm0QXMVjYAxBfMdrylrrV1zVOZzgVA0gNBA5Hg8QWRbhNLHg7pehH5nViq2uuR
8qn42vWiMy++NJyor7gIZTnn0HyWxBH3PaUgbq5Pa40RY+PKUNvlUXbdEMXwBA3zzSAo+UWneKUO
IVhqRQQsYXgFEf5rLba6uvXdRJeLZwLMpnUzU3/+z2hJaaaCJ2Ozb5WA2rW0Ju2H7wtf5iP3mtP/
fqdwHwfwi/N/LYUT26SyXVP1C0uLIYupYSKebqcwON5lpWzw6WqyfPDTemi3641sFZbCsvSLSRh6
KealoXvM7Rnr6rM5QDz4JzK23veEqBG0JozkdTblmXE2Ucz0cy9+XVhGoGGUaHkf5FzNHKtYXP1s
6ppDC6XjxnVxzGuX4ssoIWyHgeN9ENs1to2xIIjRr5ugGrPt0YL7jFBSaGzVQttQqOsqNRc4OuTZ
troKaLNOlw0gEQcH6GvsCW/1mc2WH3vF5RrYAmovxWvrBNdFUsIk69uwuV+So3JnvHGVVNH9MrmE
e8AstzY2yoW8nvqmlefSHQpFDm0WNCSbR9FkSB3YYKs4zjrN8A5YkopQ+Ram6EDbwkufLmIpAhBf
kgByDF1YBA4c63A0oGSiJG0Z4nEVGUDVMB7npyMyfpwKCX3ZuS67+LUYnzP4jBXxwzJchhqVSI5S
xpzRXVyALxdEQ4C56RLu0RInS1PgVLWhVImUtYO9f6L2FBM1IWy+QzBNAT84pWDSoH62ymi8L6HS
rb0InvZ8YtpaeHK8eaBzDBm3FrzQ2xjLlwutTJRwTzclimLfywJfc+Ge+jZc9gtOOv0B5R5cHzO+
mierrWVo50YGw+LgCLw421tFD/YhflL3+6Eqr0xgm5bUw6JwzPdA/lVDmv/omLLvBAazmCGaMKYU
oQMq/mIPr+vx7rmT2FateeCM0ljpC+iZVYMh2rNxm0dmeyDwwIl2mO5rBUFif7aT6p596kb/ipnW
Xkmc/xCXML/Lh4VCWKqB0kncZ1etsiaXKwsetyOi1qHAU3oJWA1W8q5q7PGZ78rFBFQoJ3+DEQzN
9aS29AtkfgTNEaGWUWRSdpJFsih+cW2vu56aKR7VxtoaejIH/YqrRs0ovTSrIiOVv4IDdYKPHlYT
0xHhAVNySQo4dHJVZqfZGHCNKewLm8E1cs5oCCpLGQcbhkgwuaw/et251k6Ls8p/ndis4UtM4+sY
IXApfyezsaM23fSfszi4sPtTt4mlfWk2L9pgnOeXJyN/sXCqQ8DKa05mIJmRFUAj5Hb+o9MEkUAj
KeHuttYoqoyK0Hf0WCVqiKgVCpQAffHtNMTIrtQ9kYWSt7LlP7E8CC0X5+ElWEnlaJ+9WI3kI3L6
rB5P4KoMpxTeWURvPkS9AsqqUAUMY6B6YO7pOaeTCZyRh3wEu/hNSAuycDL8C/HMmVcycIt72vmq
tFf+HYD0VE01lWoZcuRcH+pS/1zz/D4QU37CCzGVLfaejvRmIch5Hg1oRr6X2F1Pj6wU67uFRwfS
D1YJtCobuO9BEjQ1qANWXklrlfD17CCQBDejMh/vtvNNXQBUndRbsjGX6vuJb3l4j2AdMJyDH0Tq
Vw8fa/LDPKIhblvOqeOgj8J5+PDZKJwm4RxgLUigB1vCk0lzymvoRbKFgo4N5UUnywYi4XgxcSbz
RwIAaco1+zEK33GJvVmSkZsEaXNP43x/k4FIirgZM8w844KFNJhbbzcYz9jctBGNB+lNLkuxXCx5
zelEvFDSHn8tCNlv1fqM8Rb/LVEJ2KyjUMosWzKVZk7HriIfQwPE3l45+aJuwApYDdbZFsaIqNsM
PTKLdISH7MnFWDzm8Zdc3nHtFVIV9I6RTcsRRdS9xmyWtTfd9exYzFlV7qCdW8WOz/+TcxyAjsR8
QudUYpkYpJWYFPFGVZgodEIpyRSTs77GOpyMOa9r+M3MAUd6qdoFoXHvQ/PC8g5rSfvRXJlzxOCE
XFrqb0KlePram8TlU7Jqlhv0nHDxlJSgkw2iFz/zbQdNID3UNQEnA15V2fMVZwebFf4K4bqqnboW
mADsu8Ks3vAxkjVjYBCHUDonjF1eUP9pMab40kL/UBsGrphGEZavBYrDEXLUslsA20Jf6/L3C85I
8vVEsUaPhAUte0VJz2eEKRCwIGoR8TTfWAocq+4qBg5Zi1T7dwiUpCs/qZM47ewG00Rn1KHhD0k0
Ot6fCBOX+9NWLghVGpHotZj9Jv74Vna+38rF9aaDN7sb17ekQllwRKlU6yOi7GzaVlE6PFs0VDH6
7k1Dgu/yY4K8oGWfpAldZp9uGEVV/AmcWzQnW0m30p4oJ3GkQoBrXI2bllMbBpKLOTTRt4oJZccT
28Gr90zdkPF3T3d3W3uiVyZ7AOUKyahUInIgYm3xfGIDh+Gg94sDEZLvWphuyvRGZIXrGh3UckKz
XF5m0FlHg8tSLAu7uW3QOjXVtX/9stLV1KW3va6zONmyoYmBl6x7PSxHGgWay5PFnK0SfLiZ1/lP
I0XEnMfupIVVE0/2iefEnaP9tIpzv3lhocMGSag/47040Rogh8peh/VfLFlobSuUCzFHmo35wGME
N7oeYvUlds6jXMRI0zn/b35QrFrU/fw91EEppsodtN2z9T5a9yxZPJFyj/LrSAcaU/hfHlGK6ODd
KHXr5XQuacH5JbKpIAJuzoQY8xCfDQTqzXMqOMkaYbEKdIZtcvba+brN7CYhxstF8+2rFE+cNPpy
BaFNdeIltwfSuCo2gEtIl8pwjbD4gKkFufg2Q95wgIqeoIIqlT7L2O3OT4f2W8s20oto1QTtQ1PI
YUPHtOFOuL22HpedjZpvWjwEuu7+HI1iaLNK4rSDdSiAPomS1Jgu4XoQKk7g8IMByemCi/4EwFoT
P5CeKJxndrXpfYww2ZCtvXvH09DPC1/AssXd4ne77HZ6g4FrbD2OqmUZ+6FsOEN9TGSjw93PW/AP
1Ke9c/pBwCm26TErzaDJnJ7ut/qPPJ+eYA+A5jlL7YaBYTZAF0GGTzho3VKAZGlUtJB9WjTQGXYr
96kNw1iwMain7sdEec1coFgMZ7RdhIIvwAtrJz9QrAjJZCcTdSb6/eqcrPbzEGeni7lc708wsQVB
X+jIfCXi7bfTwcig3BZZrt1AO2SDyllMoxm5rZvFcH4GE9VuIUpBc7r8h2ssTFDiEgLtSN1ACq8z
ks4SjL/DZmFkX2NiK7UikiTyg8EemHWxsKjqpPog+lYMpMTFRiso6BDugd3ms4Vd73BxDIR65RvC
l0vozXr1XZAis9DIiLCoFnwnKX2FhnVuK29AD+AFfy3DbizZ7VBdQYFI/I5uocKRlYT9RIz4AXeF
k9RQ8nq4HJVt5RmXe8ntijmd5FUs+y82jDFaNtDjWumIb6RBV0kYPuldvv0wgbyq1fW+XcIcHgPJ
rclM97LicoHVQWLfcGzzzXdFdDxXklDVydeKU6SD9NV0Jn3a4hz0FZXaUvkssI9ZEb1ADj6nO0Sz
6gg0yDllWD9bQMYgPI4Ib9biBz+t5nM2Y04+x+YXCH2iCrrvyVZ3r/vJuIXYRJfY7HpQ+QGkY0XV
Bn7RcMbtx7H31nCpdrDEEyvq4dQzwzjD+3AVSAZEIgHoI7jyfhvBw+hhGBKmGe6oihBYU8zfmb2j
akXa7tnLkHjP+Z3yERqeNQU+p4IJPwLl1YaMy78zoeoIW3TR0lLdZFXmZrFGvsWWwqerTq5hkzCh
gldE2a9YrKLDc2umeFhSrYEvbGm6kGCtoP4pxIuqDw9Dfw0ssoUW2vgXKYc1C5nmAU5DgMewnKQl
PhZU0EgAPgl0IRx+AD9Hpu2k7I6jE4MLBcFDWvgsbnS1T2mf4/mkGt6wUyPUiMvFRqh9vrkLmQU8
gcvdd5AH6A4Q15bPRfxLKeW7+G+AaUWlGl8OVwXGLRApSY3OzJySTF5yoeamSwl0GRJ4RmKnN4mk
DOcPFfssSO71o1FHN5tHamrhnZloXbOJRAA6tO4MH6nJG6zp0eGJPB0IGTpsbKxKGGYv5l2/1iXr
PNOjo5nYzAf2jCGhdsXUkn8jRtCLqDRHrkuT19arTclI6L76I/TDy8ji5hMXsYN9jgDFucABErZA
cJ1N2IC6S1Q3jrsacp1mnMQwtbpTjpD4QsP2eosSvsBAS+k62XqkbbzgvDlXhth47H6rNPU2ifLh
wCBsgRReQxk098oAS4vrtZDZUYDYenqLrfqajVYjvB+qGG+iq64z2KvbFPoq+fLlLbDPF+GijP4a
rew56oUvajpgUPdss3SDcrVWL842ajmJauWMhMVGeZ97VPAjWLNyIE3XyT/94PjN9QUQBnr2lJwT
sKexuCukZDuSqKw6j1mnkDxQqU4QDsPByv1t1tNOEgoQHHxWx4e7x62bVYGQ9j8t9FlEr4RqRIcK
zDDJOS2PYkSbMveOhsWJs6JrHKcyBgPvcoDGt5pVKF0zqI4dPBlAJJBvHxE07/it/hEsHPnoxLQ8
AACwLgWIyORkLhtpc6izw0ZRzzTzdsS6llgdrcjLN/oWrViSBPhE/FS/CIxvP20kjXDlCo4couV1
UfusHWOPOcey8WvINpvj2hKRU2p1CXcCkJYA2f/Qf2wFCOn3SUavADYeknbvthyvz+wwXVITGz5c
9Wy/4O8OzDBV6JqJad9kvXs8lV9EwHXSHngKHAmrEpREFGJfyu1EopRXc/DORUckeg2Xi4RzaaTM
1KEtUIXJyz+skj7BK7RapBZM3xWAi0NTk7YK8SRNKzJ041u7KI7fzHB9ZGLQpCcw4H+3YwTX+Z1r
G+Mlfr+8GDhsq8oAB+ax6lO4LjqzbJiRDyuk4vWp0+RyAllkA5dBvzTnh6z4AQqMe8DaaiEjpDct
gwWEx7wWDubY+LUaDCHYVxmUYYK135gcygIV+kPa7i7MOChb+8gYEmNJkB7b68GXYdTzr7+PsS9E
PvTBzdan3ycMp8/ftLBi4uBXuJ9Gmun41c8S64zXuoIz1KnkieDhAN8OeLws2wsfXx7gR8sKhkN4
kPS0L7wtQyZ53wKSjQo+EBYPSsRSNwXBTIn/Q3KpwhWWR62m4neQX3pl8f2lceLQda+96IbrE9wr
NlnQYBegplnylCufpz/01UBEzfG3clpnbdu1DkijASYYSZMHlmhKNzzr0wVe2HpbYYkP/1iP1NfG
goPagIr6paSkGqi6QxCYPQ01ynTf2/rcMZjinGAAhGOsqt9VaHGg2KJNPpmhlhsJdmNH+nTDIvAV
7tCKFlTv6EQHG+MXtFjE3UFaAog1mGIax8jvsc+1PFc+pJZKkkJ/BHtelmkdSxlLZtvv8LGbBXX4
SXUj9LJf4tJDFd2B8+oD+lkm4IuvSLBp/J5qV66Hhx/7wP7ib8FTYvGlbp+TsN+KH8AuodWEUYIx
cQDZImrpBdNpKpewKHVkpuwXLAbB5ndi2iKRZU3eq4gvr2Gl2IMxW0mx0OX+hbRvjaEI2PdWVk1p
Ss5Eg+ohLG2dbuvFQypnjavX+uWvszO+uQH4u4ifTaQ/0GCzPs5ps34mpeSl1naZ7ApdsVFu5W95
LLtKTqC9pUlaQgLzw3r5a6SGmp8IKnR3deP7y9yq5yC8PwscYHeiNpgcIqgmsXeziXe9qacTXRQB
VPTZN6jyGMSBdVgC02vG5wCxlneSqx0qDPvkBFeCLuNs2QP5OUM+zeBqNz8anMofpnaISUSvkazx
/xwUtaiMsl4XQom8ogr5DI4bqz89U78vRUDq4VnVsKxycNVNDaPer5hPOzw81jyAh8Pcsi7Aig6Z
zzvhX4nwn6vRW3VIduv4xkUUik3dyyGMGAnGRHGdTB/m/WS7UPVcxzGHwZIrP/vWRKarQg2mn2pk
qaREgHqbuF5FYeJ7tsBK6af3Nt2vhtJ8Gzz3/WzTE7JmoUm2rd3MqlVmioNROS0e02VX4aULBndd
xM6HUJkeWPeYuA5xq7tNZVakJlNO26LpUpVB4JE5ZhKNg7nTL+6RBep1fNFbI31iKm4T7H4oDwXc
LIjZn0q7Wgfd7JkI1nXk145fqlBbqSjrg0ySdmSCOkKNHcaJlt1NPob80Iu2mQRX8A4jiv8/dTTz
3ef6drGn1Fx9oJSZvorraEcQwz2OtYIeqelyCnUCww+Fdj2zwnSsO7nqBnYqzdXvTIQf7ozPhgG8
LTOFlPpxaDlH6V16O+MiQgNhpMlrtZgEQGEsCEzoJfbS6rZ1JezG5obPiWXhqckYt9JXcJSiqOYM
36l6kXH2t2uPTnLlJzryPFveXSvcmNrQzA6tlNcxDi3IA0hD7VZan1K4dz0NPt+1PNRYhAhMfV6Y
LWu/XuYnij3OMM5msBwVrpMVziKozV1T55D2mUh9BJDg3IldnNj8Oco5SdEbtndtsKuYKEZ6FQMp
6VvKIgIO+fd9JKdeFGEHt+fGftive53Vm+tRD1WM7rjVTwwJDQPMAdUMI7NVmHyGhbM969EsInnH
djWywAwAt/z4lF/y1vMEoweb0W5mSd/6Ci9yBzmtgMCWN/10iMgYKD82mTqVzjTH2w3GrPAKVOht
V+omQsxuMWj4DtcpDBAvrEi1CaEt591sXuD4htq33Ty0vvbqt2AYcuw8Eg5CLYfEYORb9h1jA0xV
HljZ10p+dWF+v/FXd42hRgbVtgm1+7yvDYVbZyo4xqAgIwgnOmtwaYX8VvInJIpJPaxqAqgXXQoj
TWuHmsqJjpplCJQ6FS7dGS0zOHI60lxklH9FFofFT6s/ouwQIFMnJScO0f6etaoF3h9tMHfCsbjp
lCrmYk8jUVDG22dBw7FKe5N3StIcIFyNj5zAyZuI0Z1byivbgUHKsBWn+2d7pwXrI5lKwqgt/raD
uypXCzzOVufKfxboh628LWu0Z+6UKsBtdhRPcVNv0TJ1v3ZSN7oT4NdeZr0ObZMrvoiMaiF9yve5
HbL5B/XryAkizS64NiqiqHbeU/Wmpg/aOBE2n5fZpaod0XeJmG9AZK9ZEkPgE/zOvRxfOZIASZKv
msdKIwZL29ssmZopucRk6azpPnHy3lsA5Tlh6z34WR7Q8lgBsXsHvwiGHBU8nOtfbAl/WM6iLXOH
oWa2z30Kf83IyFuXdk7aQImrgXm+yaNUj2MPb9/l33wPxWgUe7cTtbfVUUFkHZc3rxS5xyTk9i0I
JuSk2TjIgGKsFxIxpSRYbKaI4PVJeCJzwoWblLe/kUAqWpzhnxl4lWrQrvU2G+QbCY4bnRXQ4drO
pZAGXXofYtzMNFMAe9ogtrYzHajajcG58tp5gii2ZTicHUAHDFLnIax62PYOs9l15mdkWVROFeK9
7wITtvRaM2TG3edOVhL1bHazhEJWvc+RZt35MH93dLdXFdL2YQLH1KUVdJZe/gr5mqSDQXsKMKfe
3HbuRmlClm9BDfGW2GJ8+fwJz7iSNfI+F/JyVFazB10u36whWZy3IFR3Y8haoY9YWjp3Gooiys93
m9KW67yAO84kYRCMfs7/k48S2I9C98tXhRA0F3LhVjKE3t40utZYcqkmyacWKjFfjfmGFumS2ibF
WkILvlaiEJ9xmGzq20MU2LfKKj2+bhAF83WvbznwD30t9OPr5N8iS8k1YZP3kf7txFer7z22csWu
lZfYRV+9YqCetEIfdtyK24kMQAPcEv+zurDHOvSvmdwfQDG27Ta/vLZWxzSP6YNzy24Btf1d+XYr
qvMDFdJVlhWAc+46fflJMK/XEyxAr3zU8qLi1Bf3nGdBvvCWJkDFjjgUVY7rn1kihcbmsdQzz8FT
FlxI4C5TWaJ4YVv8b7SgUcs5IV8gDGny5SSoVfCXuRUvDxVU/A8M+9h+QT8yOFShgksdyBaepPSA
BO+DHSYR2jQ72AInnlgkBFtvFmSrV3HXWw+C/2G4spXgU0SV6uQnEB91XdL+8Rn5UQrpDZh+K14o
FXYFgFMfRCWU38L4L0TZG8gyjjBmIH0jNDacvPbXcY+Dh+FU3/LrIv6jfAsiFSgNN4UOjE0IQHSJ
sNMICPgeW4ze7seN34C1sUPB+WjHpLu2EpavqkThz4av9hjxMyAAXauZmCE2Ci8CYvQgOok9XNTr
chmAlgoaXuKV1weBDNaoA6G49eN/NTETVQQlyX2xxZdqfbvspcJSUH3vQwphy3Nsc7s6NWSUR3MU
3bVyfCXPDuuiAfpyc5X4fqlhn/if8AHMr3zATwaayRkVUTOBX7L0RHoQwBYS1bg7Fe5nRWAr1fYU
zcj+E/+LiEA4fBSgqxDqV84gmWYubV4fAK5B2OvJVknS5ZZ6d0Mnqmjia5OwPAqtSdr0vq2cK6hm
yDo/4MZDA4w5jUlvQ+T4W8mGIA4lw9S4JDrsirHCIqWd2DmuEKFb8T0GQ7thSK93CO1QAD73ZCJj
fMMrNEmglWQelfhfCgnhyUEq2dT0T1k62XUWKMEtiPavbPWTP1DekpPPkDNSSzgXSBp1EwGQv3wG
R6j68j6XH1tmAHFJd7yKn3/4U2UqZowsFTc9basshKydQTllXSo70oTeznAxiIOdyJjgCJNtEj7y
VoCnqGuCbRffLgB/4KFjf/mPNH2xk/DTTuaGrghsogJ0xb4Xl+/pJewRmDT7LNYwqYlRoQafeMVG
TF4jWbPEYfquIgD/eD2YPCsCMnJcKUT0OmJXBlWvajrHTzqDU2xYLzkJl/yx+v2xFwSN4kURCNz0
NojHxSjXITfWD6hBLsS1x6vDH8F/Q/1eM3Kh0hcKyiyo/89hACUCJW3OtMAZZ0HtDF7CQBsVqzOw
fd6XrWE6eklVEJ2Gbfx4CFr9goJ9GetqTFRtVXww5wDIL4JqWMdU9THKMJmgVIILc+4icZ1z9Fqw
opZXBnA+Kp1AYFZn8PKAENduLDFyAIXp4zZ0ianYLpvob/Uc0SO/wz6HDN4WEGKp6PE0vU8e2UR+
vFONMI4AG/yQQWHMd+UYqP4hJ+NfCKNSS+C/iPCq6MyC5g/K2ZL0HBbowAr3fJO5TVRql2n764uv
2fgSHWBt+L8L2pxyq4UHYPZi9Rc0sQZ4BT73rZSMUQhkKJPmVmPyCRrLjXH24k6GfNu/rld07ivp
jiIOnb0tHJVqir7VHkhi17X2fXFk87damqj9OJXP1ZRs72tAgqRgTrZBmEVFuHiZ5RN/C/q9pcmp
XOjULJHY2qpI+qHDVk0p7/v0TcGQmP3b4pFc4mWXr+kHV19P7xNngoDSRM2u9mrm39HqtrO9rbfd
pi6iD0XUm3uk5qxEvgous9DAAMarbtUALRcW6ei0Fl+XPZtXbiCblpoMESxLSZpuO9kBCHDZ+GAF
am9XESsyzD+Qxnv2PVQ8FpLNSW6E8gr66pj0D7VAa8gp2MyPwr5dnhtQdcE/BvgTl4XE3IuLKE5o
8fDhuqqnzCHb7I74V5M4LeiscEiACWiH3q5q/EoMyWY073kU4fskUGTiTWQ5+og6UGFrhGrPltC3
hFmlZnpxbTTiZtOKcYCQiEXvcLwCcuAwAzZ3wA6y9KJblB2D0wTWQz7q/0dATPHIwrxe1rtu04LQ
lBWml17c+6uab5MRgHF4Ln7GunrJLC73yFfSmbNrMUVXWwzKXAEfYtSFqDgFYJIIt7uaJkAa5G2W
bw6hYfUwBeB3CT7KNW3VO7QIWAsjRM2DB787hXxyb96UQ5Og1UuB0OPF8L59ET2zb+aV6jRKjvQr
Pi9yvqEKBrI14R5G9dr0SM8bY3MpT1x9wBpGBORTSG9O34DHxQK/Q4TkoNSzHgtt0Ad+BJrfanvm
5SiTntNc2jo8bT6fwCtlf7hHtwvxtiQe/Sw9TOrEV2vwYzLvh4C76cFxKbv6UEU7NE1udXK46+wu
IyFQuFNM9b3tqPCKpzMnAnvMdt+X97VYJJP+w3Lq5DKfDTc/ng3doBPkPA519Hoh1svZrPGntHub
CbM7xcMdptgMZ21DZKtDtISWDhmSm8lGzYIYtyTfUH5fwH6Tkrkj4fjYXWAbrN3NEcraiBu/sJC5
NTBF/gPqvGKoBRYDuu8mQvY60gWj5l82AppTB0svRz7lynjAo4EQTqAQStjrJjLvLVnJfPQ/nrum
cf8fWG4Sq5Ka+WurkfGviP/ZWmy1AOyucMTEiIM18U/0PbQxToMyNKTffIlQw0+inkveOYq3S++s
Ii8OWWGx/olcUVzkQuorYXCxmInxjivy86DJ76qvlxNOdVcr7zxuPCTcOW69IHRNb4iL8mdfuj15
wey1GGA2QMgj6KMXb9+vjgl5RVO8T/PvVs4MaOSvKCtzyn8J4Ph7ZmkwvqsY8MUSlRSSB6Aol8uP
qExX2TVMKPD0Wke6i0hbzGxwn4BFA0SsVyqsAvDYa3G+Qof6AfakHh1nrn/KIVTiDIyz93Pi2izL
ZNoVJ62YKOrwO/FcnjkxNmIUIdlyh63J54KLGShPehOrlCvSvIOESy80k3ktUzc7ld6ow5aC/3Zd
pjX5hWy7xsKd47UhSGqafhAvTj1+BusUfhsm3eP5JLxxD/R68hsPuN283mB5SA1b6CIb2rLXAkFn
xLeLOanyN7Qyta1lh+PxLYi8KJflAdizorb8gEqcvgt4vIwfuf7SsORKNW7CpSkciv45mTVPLmzy
dRE9WN0wZtf9E62ufDzXXYJ5elH14CLb119fzfhRy2Fb5ulqRUH3aJvTMhPBIXh6T6q6tcXCl14F
RoamxIf8sOGQNG8nAOeTx6MqLTLbeCjnDheIn5hymqXEZKgdHUuRhpW0kvAwI+86p8nN/MIdwjGN
5NBA9lek/+LNDX72xsibykTRhnbAK1OY5Obdcd7DfMQxn91H860VMzpa9lxHz1nj+WIRnHGjafyH
1h6KPkilU4aNbY2KC9iKEHFW+WLM+R3RqjOf4m8kCQ3r2D4MRPW+QHYfYA8nsb2b7s1GHihM896t
mUokL7Zp+Xn5Voizn8O/mNe73SGyAe2abhmSF8wMUwXT6Igqp+qwYj7CjyLBmCVgq/F9oVnM14dH
MeMLtV42g1o/Txzc33qKSHT0oH88TrJIZv8BgkiPlURH8WUyk68YslbfFCaGVZVKQC9Tdo+JAdxD
7/1VZopAgDR8I9u00x2ueJKbYrk62bwvY/L23KJVuDAIylnpWq1sc3YEtpy/3uGky6/XQJyRgHBj
VIJsoK8+CcHUrvzrTr/f8GqmvlrhO3aPUtEGG6zm6cFHewqrUWRldgiEo66NBETv26VemfEygYCL
DaoV+kwxuiQBV5jr6IMceUFN6FpJdNxpIi7GVIPRKD8dCn+Fxd1Xc5BBK0Hn7PgGhDgCfMjwD3+y
U2/5WUTtWgPm1XBjgUoXm9MexS2AGDhNhyfCOMBLBMYQewk9FhbtiPdh+PiKxb085kIo8HL39CaS
zL9WCtgrdOGsYEOLA2/4x257+wAyZ55Ak87a9t8dO1qzJ+IOe+h4MSzM8nyr3AkOByfgb5H7U6KB
M6a85v2tUBU5vO8OtA3aRB9vzo1q8kJvweGGDz2IQj/4wggcYxTxfL6W/ELIBq6gUBeVl70unocO
yopb6F4sMBF2DGHKLl9X5Z6HGdgosXSfTKejDlvPCbO/83tptGbyAKqyHTjUfPOong3fG8wUkv4T
X9XgvFGylC1Fwfh2Fz0DgXwRqdWV22hqnKe3NrfreJVd/dHFkNGZlXHPu/6byFa/vHWvxHcTnXsM
lWK91pQEe3/TXcCTCP3okaq8pBuu0JXYYuwBX/qtj4yRVJzioBXEuqIp1MlMExkVu3dTcjvLNJ6A
oWS/d++R81sb9/CmisdWezzK4jClH1+mCjrxVIe++d0p74v8yBUIpWJ/3tr5XM4uTuSFdkvDMG5R
CozULEP2NAqgkD+pd6P5QSLujiEGq6uJys1EUjmPVfnRbKdPv+YEO29d4tGD6jOyfjhwFC2IdeYn
L7CTxp2HkyqX8oQ3COazc95OcvPgOiQNXM2RN5rgMaAVf08QhiRv+Snupy6cDm7hKqSst2vUl1m3
juIv303G+4oYLvjsSHiU4f/dnvP3mPYEkjNkrdl1+zoy+HNJ3lJvWuazPSprV97oMsaB5lNZFONo
6hgSaF+peweJs+kN8adztvG86n+znHSqYxrNUPBt2mrOgR88uILM0pTqzMfgkdUnM2wqmQJmPXLL
PH9Uvk337zGntQ3oJ0iVlQ6gd4E36NYJUgzV6doO9zFKVtjBFDoPP8ogHrFdaBgi0yBxcjsorFZD
S8MZxQPzOIyI7xVtROGNKnd/0nwKJYIpWMDh4Et0O9cgAu0u0DkXCh5uzzdWxDiEDryMBZKRCeOa
5XvPTK1mEhUxylaTxWAlNsrHn5u/MVtoGxlvBvPvdeRjkaC4wN1zX3M5PrUC9HJ0y1hjMSd0zJxm
o7opdCK1Yo5hUWADFooR85Arqxa0HK5bX8yeZHuawKoeeLy+2D67lXOGz+vsLWFtJsDzPXVMXX2I
IbuZSPuKE6PSs+jeA+rAP6KS7jJOd7uGPHaQhodD8Rg+RqjKIxqphv7fC43WyWwRf8LWCb6ekj80
/g83pA/mxa4FRWVDqqOVrSRaNzjLm7vVKbqoeO1I8Pq/slbTNi/Lt3Ymyw7tK70+kgUBftnGj+kk
/sYuC/feSfYWLjxT6snICVKMLPzHkZLdXKxa7GQbSqo9ddTOJum69GbWm4B5z4Nnr2OqLXl7k8v7
a3fvRfBTld2Ufu8SN09meV8p6dkOHG/RfDDMMQBt4d434hLOT/aikOshmlWjvVXlFSctKM3cikOw
PGMZMc34+fw9TGS6SkYYAvCLtcf2G/vcMQkYa0SfdL84I6MDVqt/FdQDE1WdAtD4iquYVDuYLc7+
fKamyM3a6srXxZVaIcA2bOKxOhG4vlfudSpwj9uvZvi4PVazub1HSTdJIlHMZ7fztMkkW/FmpB0R
81Tm2mBn/gTwS5G2Erpkv1FAKj7zCHoQuMrko5ShmbeCzhD7UNM7le62OoOISHGas7lAUEtylbUj
IixB08aqDU0L2Mj6vid0KLHlszSnLFSFoi2c5F7xuJ2dnTRnvfcsEq+ZE7yjO+I538IIdAGMmt7T
6UeMgPndrHSFU4WiQ2RKClFpBFp2jiujA4UyyZVzOydHet11yoXai8Lyn3GFpmh+g6QfkORcoaDs
KWEMFA7uWkVGClNIDhK8rF2BVAPApIf04E2oAEZN99iRzHTn5lBPbH+fXP7uwTvnpDFnH/+Z2/6h
nLu2UtbAGX4TUX/2U2Fmx1ccuNfEe2uCb+j8Ha/jM5grLZqXN4+xeHIV8KXc+okBx05V/3KeFrWI
fN6squyyhBTauQIHcIsA8qhlordueGWgBiPLhJlsxlElGOp9/JUMMhNamvpMGUOoLti29ooF5Hq9
sHFyxCyL8fG5+2IK/mQcbKzVenSJhN9fB31DWq7POi9eKHOPYJzP8mM+0wLiS4X9EugfMMfTCe9L
nLzesiWqIndnfBPl3UKLrZiSPCdfjBewnHY7yz92o3VFanFaG2p6mSchysLQtYQlqlX7v466E07Q
ld2ZFU1HNvjDP+4Yng2e1wSvMlqMbyO/P61mKO+nJmtTXoUMtLEgNiOrEWTq/4oUoZwqMkB84Jy3
UDK47HWYalxCewpDgH7cW1kPyFfv/9u+61iVnMBWddQWVnH90p4T3hOiKxVXp+MW9v0MtWMjNsJd
oUSKUzxFjkpK3pT/UI8JWJobSQkeebzKkDK0HfUp3Zn+qW0kLAyRzkaiMXbVD3sbmt+mdRj8i6U9
fHihp3Jf7Ug+T++MFu3x/dWUqjiXwQLmUDccKD0ESM8BJZBtvWQaj5RrtbkG7M0208jj94s1QG1j
+fQ3pH+6rESwruQoBXonNpRo7XpNCHG0vsFt3saRBq+jVkBUyC6uQMaIibDRHcF4wWo+R8UUUK4M
+AQVqpvmaIfvDkH0QDVSZ3T9LbikacuMLkoR5LV0BkxPLKAxpfCd73xjv228M76q97gnerLT2pTB
V7y56YaarBQzOU1GKmC9yHY0rqpP65g3ZYcyM1Q/rO2diQwprQJWF7VAxrdXL+HWoOb0gZ3p9k/o
zv8spff2ALxc+sicaRmAi7GVKQnsLGUPp1WvwU2i9aPh3Tu5VMoHzdKU8tb1hOsIQs2YkjXeRz6k
2ADuYdI+5/Lk1Q+Ph58eaG8eAvZ8sDVWRC9laL0LYYKmG6uC2KHJp1IU+F+uLn5KIp7VT36BECkI
xo9FBeSnzoB6YMVUiUXmsezkAvX37UpVKJeG2eYGQhuhGypwVeiEpA7ikG2S5NqI0zDEGvI+TW1h
Yup2ySfdNDVAP/YSAFxed6lwIdyRrUUwZ61cvCQ336cDv4sp9oVrGOFUuNFVCW30tLrw//fQUfr3
T9TtB+Pz8gk/2oVzqU6wYVuAiurZEl90ZrFfrUpYjGq6/EFLuR3mTl5N4gL3frLxCROFIUFAV/WU
7lBoxu8Vhryj0eQwQmB4hKeFxpXC0Z/dgYh6jv3yiftGH0MmECTg1qxFNlj6YoWeaZM7msTnYWwB
47lqYJQY4dA+TNCmNjhkaymi9KN2JlJ5BNkZ4HUuetjZEyEbKwUk7y27WuC+PokwU/MNofsWO5WO
bdoUpHHwTCFVQL2VPNQZ62LO/S44kyn7eflqyyakdjPAwIOgI1NZ+zNt9mIo4QDEM9WUUvR97Fla
y5pN+vvfsRDXab4C+3bZjTRduwdRshbxFNUn4UfG0w7D1GPCTWriZFXACSqSXUMsjrFMkm6U3v49
YFsHL52I4HUlrEg0gLQVpzyIWEWyArxPn0hvd9e7IEfxIeOWzgbx5rJ3DtuYwZ0cD6QE9+rORVuG
E7CBbPSshpX6T18Yj9Zm9309OgETGJS74ode4haqrUu9fYN3H+c89FL72DN3UYdOxjynMwGAfYeC
t3l87bv0r7WSXHW052wSNVQvUXoedo+MiDu6V8eusYUACBsvlKwYZqffz0WxCfI476JBYkjuIqf1
vTt5BrV76cEUjlwZxTtPywD4SMVf8KhKVmSLJFyP8i8s6re9mC9plXpulOMY+SCNOBVkhu/fhI3B
t9Cz7aPfYaBAa3e+57ZWeuJMx6r/24/zvT9Ua7itMYJH3h0EFsNKO67rjc15btkgHjC0WZx0P59x
qv73+OCtIdxKwJJHbCxSPtegABNR1b23Io2S2w62D3wITqkSMyxmvwUetYFmQk3RfX6o8AeCvQ6K
fe09msivyeQ7tT4699ANLGH5fpapHA9AxzuKcbja5Qq5pMJm3YGK8OUNInDU4bML9qaCSATqtoWi
8ugsd9LNoELr8MIvEajsh8Xw5o9qsfLIOQlwFSvN2tMcp6ZTr+47LHPDls2v/o67zTVFnDvgN32a
vkqmUuXEUhneFWFLm2Kg4A+2FyFwSZRJa+x4og4Ujcx2w68iA9+v757EuITmIk0Kwr1l517GuHL+
mL9hEQ5vczZKWMuKlIPJV0KlkZueq5Zo0t+uI95c2tS2ZJBPVOuEMRaTmD13VtLRkByuqG9qet1c
1wcj9RQPW4/J2CRj8SbSMoiAvCgMKlsHMp3gViCr3UspKc2bCDFfm4Yt8sXFvJ02M4RAtOurZ1s6
ItihLlfTktw0JQmCD/4ceaI1qzpFeRHsOMnnzrrPTmY6LCKiczP0NWfPECOpqCzA8A3QtASwNS7q
lGLoqRwsggiUH/v6H1HdnpkyneUVJIwg1rmyjr1Rcner41wUMVahWk2u5r3dF3sNRwqACdkJYBxk
bfp54OTSuXaXbENhSKadxigIATkZVcYhBB0qwmnNWGfvMa7k8iapRcU+EQliBcB5L8WqQOakqhQu
nNQtgYdFhP/FD7NODKg9yXaD4203SnruF/q7c+0RN1+9wtqpeWTGNvnKXpTH+bIW4g7/QSnAgkB0
XFqXj8kttTvFbcoHOLABSlzoFE8xyX3sDhj5qX5YSaJH8PKByKmDTcX2byk7LUNpBJn7lSE3KLoi
6N9+Muo8bl13vdAny3Ki72eDpoV8j2ZgfHtJv4eUN8MnnHiFmMEjI3T87TJl1v1DflPZL0spcBW7
BVPqtN3HZJymGgxHwbd0pWcxH/C7wwSXdNwIN9FUEmr+NByx+Hc+PJl2KRimt3JWC4QTW26yoxTe
9feSNS80QuO86GV7E+IFfW1dwGAOoNUCg9o9gDSEx4uVbvMxzrKRP345Q5ZOlE+lUARntKLmMtFW
eJOJILFb8XTujy9CDVlEYTJv18sikWLxnY1br3xuj5hU14yYmvjELGu4KfHSmMtRYH9JPwDelbW+
FB+i583vsegokv0hKf307yB/l77LlBscVXjyVa/PTM9Iudep9lJO1NqlTH8e8yN62iPttUcDzg4/
itxa+dYwEVpQr2fo3p9qVs8Ap7tGHjIU2GFJkOXUd6zl7Q9SP0egdbPfkKc7KOwLE6zJossNHJZh
/FQ6Zk9AgfTHqu+zRGWBx9PcHUYHtlAdX+6L15/IdifnA8wx88Lrj4VVr/jEGRTt8z2U7W+xKSa9
//HVo4n4uNEaO+nci87SwQDmJ33NHfE8W72nws8AhrWGwKW3TWuL6QPZgONnScn50WRx8sqEzDtj
d2u5wau6cCwREOtx+OlG5rU53dtFboOcRHVpEbvslJTe2J1bIrBpmgEJDmQm2FD8SvhuNG5/yCIm
PqFjKQGVtiMPbEFWfsoJ89bHJO+efoTOgYtHuF6ww1gPqMiKC+ay4CW7bG0DmJtW0EUcFZZcIHIv
0m/DRZDmedFz4vFGGEM9sywjxReZoY6e8xGenB3BXToXXhXzcprto6/t5pbMgBLcvKaWCrE3xHcn
BLRV+mni7tkfyb7ff+IrwCLBa+kaqXqPyMZPbPLp0mVOKpaG40ZC+pgXgWwnMX57fTzYGaT+VYRW
AArdFd5fCdUUmS0bJY5B4jyXY5QPMuRwZOJbihrSbWoraaLNvH0a1BVcVj7YePm0ksrbIhiRitTL
1V2JnNMJdLkZECcdDB3tWVzSp+29J6W5jOoCmOI+2JQntlnBO2kHIF1nP1yBwuCG8yp2B6hwb/Om
Ck8nLaVL8AfvFZTse+ibVk2qV94D5vaNy7aPvl4syRM5wqMB0zFJco1JioIetFyzm4EjaDIaubuC
CobSrKsRf+aFBA4ajaEcuccZSXdggkDUV1Rm7BhTw7lMgSMkTynaLVkjWYvtWu1G0l2s1AUVQ+Jn
RLilNJnfOnNyzIhBDFcHywNe3wysuSWnrs9jxckTnVEnjwnUjs9FSzZwqMC7N96VCo/OTCyzF6TF
pnRrw5ofaBjytMCLhZrwEZuD/MEKdvm2wCbj4c65IVeaKHPk/4HQBuBHfVvwN/aSXa6DDVdqP1er
2+/Um2ShtScQgFxLUC2zwY+8FTNo05s0PqU95+njSFpObxwUnTOkPjJa5MdFR6kkzzIZoBLJ5sJd
ex63pqgjed9P26393dNE0+ApYOvOZuTqahyKRRdGF+edmGbtI61b4fdp8YDtcS0IsNt3Xe++eq7I
lhrtDh5Joh54f6S79Y4lj5q+YLqXNCouPwKazqj3MRq05e+VPXnZrKJkpYqj/znUSQQ/xQ/VPcGA
3aSuQJxw17/HC4bzrZ1Xu8OODyJW99MheguDdgqPdij9PTH7gtdDb12Qfmi+LscLXvO5hvWDernn
55NDWPBj2Vog0ecn5i2s6f3TCAj1Xs25Gyo8qwXZGmQlG7vqz/LheMUpStVB+2PDfpluOgtzN7KL
QZPWtYBjcMAsnRtYi+RMX2qFjtvF372c2wJPeYXW1OVDndOq/edTx8oqgmMvbKgrF/RmhE0VYS0B
jS0/jejPgZ6aTcvFHaANTAmBB41NLanU6SjbuF7g3VDJ3bXg9+C4+z6gcqRPiqkaMIshHSa/mdrY
Mlv7wqSqxQ4MoJU40M+1CMwSzlDTRKfpRDhiI+7I+inaWKeiiLZSCgBWpriRnirw/JXBzDAzTx/R
JgzbebgM5hwHoL3qMVUFKS8BDON6t7GLSGhFneEbQl07yObO2qCf6XR5xTHlu46Gblaj0Z0uMN8h
Warcmy2QZQlexXMv/ob2JFaVjYRaXExiDzRol4EebisEbMbZO/euidMQLDZoJjYeaOaSguXfo93c
esjt+v3ntHaIwmxzV3cbwTw1cS1sd19hLxnq4q9KzZAl5Uw3cVezb1KzyhNMBzVRa5qrqvXH+zZL
RZx664no5EyFfZzfoMKZAvgr+asZgb15dgTfl/ziKySdI5k8bSpyf+Wzt1IQfwQSqS/I9ihsrRrN
Ykc3X3O6W/HAEhtBFsBw6Li3bjQvBMiRzrGCj4DCxh1hkdB1+A13L42HDj1jsm1WAYCqDyTutVcm
YM+9zL8+tPeH5LagKuqj6B2rEoLPSJu3CUfFGv4F1mdod0eP7KfgXUQjNyimMMeXvZIRuxHjfhK9
cD9ERcNg+z3k4eaa5o61dpvs5v2mJ+RItlZf9gwK+mhDrOzgUt9ZHxIe9qiQuYsTEaHJhOMNGiPc
KPlIWMjcoIQXRbAKadMDOESoV7xdpU6nFZeqBj7fbnvf2SZ0dWgYsP5/o+0rEejzCyfCOdt7XkwU
yE6NdH3HPGnrKin6DAT82kg7Yg4vt8cipfCs/SGEh1xHuPGcC62FoN1sKAgtaWO9vugz/cOpz1qB
/XUtV43/tLLpunAcL6m8ECDmpo9VrgTigosP6PE1vU3hD3631pe0gRqtP5atARCbxP6nGCVrVoIU
JAtfl3E5ARCcarGi78xYhz3HCDE/SpC4ITAo7O/85wO3Nokg8NRdO6+fogrjSxs4ciCi+5TofA/T
woND4R6cGakfhdA6Bmhmxu/hBslVPqkFkI5+wxROAD9loydsXwq5Eh/Iqnho3eXNvXbgOXW8H2MB
1KrH9jHZJ1hfjGCOSVSi4awkvCSjQXrslXSRT28Abu1hEwjW+UKYq2FSLCuICqHxemabZscXemW8
n7XiFgJrUng9n+C09KjR2otQXUyNyooPGKirtDhAPgJHa9nOJx/wRwJDHIOpEi//V8RzOTWqDr0K
w88QmZUAbq4Wbj1GfyxDXMJhgWu1q0AddVUn8Dc2YxwYwVp81EfZ5hhqdxCHD9OyV64Ik85ZjrYe
VVoPkqBHc6cizeDjxZA2pR9tAdkR2pDm/+cHzGwBypuS1kDS+b+9FI5Yzfloh+zEnKkSLnZy8ybh
E4Bw++aDLyE0rOoHcWDMyWm3EwJIj72kp5QWhNVzhPBJj1c3Q19rxMf4w45YEBVKPxVhLpGIbUrB
0NasFIsx8rRm69uo7lsOZkVTlsaf4v65M/pnlGUdKgCSI557C2PhYTuJFhM8kcPjNwRW2HyuRFwR
p9x7muTIXjIXAcr7D9EvltlrJUvjDRdbvGZGYXLpIfcS3a6AfSxgAnwxfw+mveRjj4w1RSWASXPV
dNuD3aLBZjfX8QLlXc8lEXIOLBCq1Ik/EjNuTZRUBmhwBYmZoXqsd669TtIsTN7QbnoLFyAV3nI6
FVVKzj3dAXkkkDo8Nwgxx9YU2MFQ57/Kj8PhmmAHNaZR8s9EPo71bxtsr9lSAuK2Nim6UaLoJlCA
kOrzX0OxeIGKqTJ7cp5n60XPBIooqXti/T6BIrFEelPZKV4NSE3UzK2c0DnEH9ClVPicnx3ybXij
G9OrUXg0HFoAJda5O3ex/xyN2+MCqghDR2o1PUrqQTnDDgKoMroZxHerGWbmmY50Se3g5BWObG5v
gvO9eTx822xNjQIoPB/UK4s96ezg9u3rA+0eC8AFzPbm0XqJ1mNEZ0QyO0S5PYD7CWOgqwW6gdJm
fpTxWIwr0E/4sjf42BMn3xEd4lwxD8EBNRL5nfpJ3Z/V1ABsLIhoXsKp3X8vHC1D2NXudyduLHab
UjCOFNd24/8AH96NS5uTcBoYWatuexXINYlph3qw7U2GGuZtZErBuASScMr3Q/SxheSjBAjDqsHI
6H51EleqqlefzTG5eCaXr+/ozC1WyZbN5z9R2hmA6so/aMJ6CgESyF+vijWqkgUv5r2ItJBIGg8B
mWfda1gkq2LwVflv7rtXbj8CAC36f7Jck2+ep8QLMj+IP3T2KgRrA5QyJJIZpNXaaZ1w1ipmjvn/
BRRHpEG53EVuXqyRVpkLxrUWTMLmOsDMlz96JEC1B4ZKdfCNqQXPyj9S6t4iwTAcCRf3w6jYBYhv
lKtk7FT+EdROd7/qVrtMDxi48Cx5v8nbZKKT4v9EIeeIkJ5ZreYKs4tnrEzPic10//Fc8urVmgwk
+KFqgLDlMaqm19hxGI1YKipLzgMnUgAS/ehRyrpoCsv+KwGblSffLjENiPy9GvQnBGyVJHrYL3ju
Bn+7wtpd56JEXbjhbdvmcqrJDzZcRw5/1i0KJFgt12dEVI7E6bchS+gKIyjUFp1shw4BcK00D2tA
858D7SnSto05GBEuoPwLRgTG3nc3/1PUG5TKf8rts5P6mw6HMRHhXiq5y2XQZaCxdCt7aABkHi2h
pLt5gTsisEEsCEefXvkAXwL1GYM/UF8pu+sMqBuws1+AOUT6r8qar3rtAoBzoag3LW2VXacseQib
jY6q9SamJEGuIvB2cVQmk4egIJ7k6XV5Qb9Dkd8FUH06IEjjWe0VVOYg7DnAaPV5U/7LXNe5qtBE
zEPK5hvu3k6aqCsbwa7cwMK09rvL/yoG73NQmXL34MBi+5eF48hoJGLH2dPVrz6kMO53DQpdmeYe
VLaq48nK9e1xr2u6nho8FeWVUzUuk99tZo47KE7KIP91o+Ehx8RqW5BCLiUTin3EPogG9y4r/JVD
mjQyUdinZswJIXELQyJhAgX/iQOfQsivVavu4A+URnVAOCD++YnG0hvdxAoZujEnAB7x8wT2z+5H
Ura/1g+0WPrHB2QJREYiNgZ4pwSkYyhsNGnW8ZYk7cwaMJ6qaQq2+T6Nd+MRoe6piIGEE/LOJa5Y
UpQtzOBL4u8439Bo3d0TA7Ci79jsSfp4aSetpDSOOi2duuzf2wkfFk5XqOQm34FOxz5roZ8g90Ja
Nq7dfqSUEMBB+jSv0FDuJLJout8L5EJwQ2YlSrhB7+cQOS4d6TOJObM4I8tE9e4D9m3yo1v80t6b
+LIZjAu7uHvq3OS5QGSjFqAO/NMFAghP98cxjo132pIMmhu4V/NaJ2RFNOeB5xKbaIsSLeuDJlHT
J5f1AEScFY1HRNq2nz+EF/vr6SzgnrRVHYBufiz6gr5xid4YTH8VRZ5KfMmkZeqWu8SU+kvosFW3
5sT5Lx4d9W6q+ZD65I6HV4yYDcVinkzflw8SfzCv/PW9ntPiH+14R/n0k5aZTsKP/UQHrYT+q8Ip
ZRcX/+Rc9kXjQH3CLtTw6dqNL7SaHYGnYWOVoSlf/kp6K4ggqXiwukHUPJVEQitp9g9u30yH4vPs
nMdbZ0IYUeIGlcf6o34FfkCtTK0MjBr8AmbnVehu9e/cySBo0AObn4aLYd3a3lzaGYK1007k1q8V
LdNfQNFmDYpditNk9u0cVSQTQs+WFR7jjsVAiuwqxPRjY7mw0pYQOArXBaeJmgruPkByuiWkhlpF
bgvO/P3wz2NlT+wJ/E5iTdx6lkEZSlx/eKG5kFCs9zEIwur3nid0euMGQEL0rd9t9tdZcqzdmblW
mPyUJdc0+O/16AJqHAFlcxbWpzxYv0+8BY9W9ymp3z7MVS9b+bip2UpWjFpU6w2ELN/IbwR3rTkM
UFD5hbU/xAkhGl6P6bP8AA+GTBoTSTpKh9JSQ+bzWs182xH8PwymFycknO5Pts8irIqyrjM6+l93
9tY2qKsY1SctxlgAXmX5bFNJ9Q5KxJK+UDhg5kxXxgGQRZGDRO0mAmfd8eM5fnSbG1/YuUc1K0zO
bvqK6sLIXpxpJHd5XA3QW2S9W1VoKgmjeyzGDTtQ4AheP+eTtV9/8LsriZXAn8Ot49lZsXcZ43QS
lbfxULFd3L/PuCc8FAKrLDoU1wrxvkslouaArClZsHBw1d6LsTg5bakQ3GEQRd503rTBiugnKqlT
mFkrlYDYwW7xISJ/ojKzDabuSn+6Ll7BJezPRaxJ2j7Cxo8GWMXuaE5QeQas/pLz4+EidVGAoysT
cBu05FVfEu56YyRNJwLCFf7iyKkojmK/6IRcxc7r32+shE1ZMll8K1MmJhII2iktZcuULXmGby+s
M2UOzbkGHe4BckmqZHoGstllBzA71kllnGlWdaX3VskzK6XVAx+hVr4BvMjkuV25AnhVuF76T9Y2
GTM/TXDIov4DbS8raLaiHeGtqczX0+9JQFJU7ri+T8a8aNHLDrd708N0KtjLLLleD2lLG0uthz/W
l45CzRzoU1RF1sHDghisfZb7anq0tDzt2pNPJlz0TT1Vw8kfHvdYKG7l2xJA8JWOERbIaen+jPuv
Fu3TqJMlm7aG8SPixdtjcfEnkZbY5OgwKk6xZ5xIgfIOS2IOYPK5LcvuTf9B/tY/q1srBnHFPkuV
xWUAM91aYnuulHl2ZWMJHpS0Jb/91SSGOzzJNkQRuM7hw93F5ql0DhADdwJys1exlb8OAB4GeUBJ
+91uqNyOqO6tcXFWWUGzgBjnyeBC6Yh/xBHXTXy1eiy8znw7zuqMNLLQ3FpYkjZS+7uX4sD6took
MU7mnEuGa+2A+rRyHMiPVKlpvf/x/kE13YxMSpDDtXX2evLhKJrsu57NOuigqLxkBb76xkonxnxw
umZPBF0mo/rYUIDhz9ClDSPWCex0kjTRPWhBdVPpot6Dz6ijlWugqgp6tvWcDSZHrZ1EdG2TzpFi
QviMX4qm6wMf/0JpzOReBSy/lv3vGTsPPBnX01IC9fW9bEhDTuUmZbuPA6oCxtjs84q02NzNsLmV
4Kam1CPlvy4KQMPQ1gKTFT3ZmPzhRLFgBlrSh9wznevfzVCE799u1dY558KCJPVnfcyjgiJew20R
0OJu4dbmjUUui31U2uHV6a1jXQ+a+QX4KlX2XF1actCtfPwiJscS4zaIuzbukSftmk/v/f0cEh1Q
A0LPagp8IFKMFgSIMRtUvTAi2gsEDdn5doB5GGngeCA5dd79okSpllh9ZlUlo41LAb+CUjiwSeUT
EmH9vRy4WX6BPPGBjo1OI3a4vYh0Lv8+Amimomz/lJibMkAkD0bEOwYTVzplkGaUBRNXSD6Nj4CB
nZvE3VjNAwUyCZ3lDUNiCQhU5kcX8qdnoa3tuTjvo4nEt/JFI+uvqaxXKqrWY1Pdv1W0oQPDUd+H
3iW4k+fT66Z9SQ9NdLhCtUvQpWID3qzGS2AgutgLBqlxYuMRA9WNtbklPTmOTr/GiSu8QNQRd7h9
WfXy93baDXeauouhsKWF+4UW/0HWoIFj8I5vZGhetKPEFreljgKq9c3AWunXzVtgVMgfHfu9qNFF
7Oy8NocnBFeE8BhJiXoQzRFM0y9dPVhiZaB23KFX+RE+j/31AdtNKQ5WkznNFqUvz3WrtPAkFcNw
FD4C5ng/+tcKch9XVdLwkWYz0pLrF2n8aAChBzyrU3v6fDIB4Mwm92C3V7CY59Z6FzLYTdkLj9Bj
qLql8ayW+Gkkw/8VvIqZPixyeYWQ8u7IUjFzl5E65h04aCw4RKG0iMLL4Tv07LpI6iyImN2bPsju
fRVMcDbTwtVNxEKN/NaCdfJg+ou3Rj2Fh/8s3vSjhGqp/9TO8f4NSUuEbmyFBvGfI8slontkLaI1
Wmm0zKVudpNz0xfov829cpPRL+oJ8u1AfgWFb30haubi2qjhipuajcwBruxpAym2BV4IsW0yWovu
VNCWgSthQNP7+C0EriqhNzwf2nEaFVpopAPMhM78y1Xd+6TiQGxKvkDBErpxdnwty9yjBKbu4WvG
3raQHNFdrR+myBxXocPUuiNgNzF68mX7fXix83aYxCZ9RD7CAeRrThWb171h3+RulD0XDllDoIUr
ofwrGE/6Faz9lBdxwkV5GNSUCXEkG8ForKbqjTcZCfIcqhRUeje9rA4jsWR0CV1O9hXvWbVIWnUq
+71L6n+9ul4X7gKzR62ubPmNSKyzmntC3YPU3eJVUuIUz5I20Fvo/OwHk0onZRdu8uk9TRb+zcid
ra0z3r1BLBeICbVB5YvOKILcHVou99rt98yaSz8i3rf9jTDOUmdVH5bitgdzUoKg/WpZ+pdmX1xU
s3wJpYZSC25v+mao5v3rROc1iPM7VVJKAVsoVXaLWzzoPd4BavRS30si1m5Ki1k2FZmNCyar+nyh
9ZIUgOz5PGRw7+cwyapupOXRFNU11q2hTQrgKndCqCHXDv53MEtv6p9Y8OlSLrVsZU+Zy3Rz+FaM
gYtVUiezZ1VjwpbcejEEuTD/nq/esGYTYR11bGOerA8g97CkpFw2sSADryhWSzX36eSmxfvKPvu4
slOMiuXNz5CCoaEubqsh6Qm3rdwqhPeOiw7g16sVsu20H+qzFhkwS6UK9+WMt5aN3HnjYQPB0d7P
yZdXEsmAeqzo7OIHTlEVAm/yfOSOVgnQLHzVFNqFFyzdxkI4eP7IldN7uXvcyocDj+HRBvJkGpL1
NWn7E15tTFc+NJJbSCIZvW45KkxEWPsw7H8vHFqllRU5pAh4UP9KJ02Z+Oijgo+4HmW3t73OPjup
mgW02axGn4kkM4TO1j8GYrl2rZk7fuPbUsVNIKogD2sFUHCzHMfCl+16Tyl7QE/d5lFrK/cXCiV5
B9e3XrwgBK4N6jSb1hWSOfB0hqEbkQkPFejdBohp18pOW0Bt1eNKlYqc/iCpQGb6STibYkwHneYk
W+AR92G307i4BYp8s7MdULqZ6Fg+2qyncGQYF5ArLg1SMs+b5jkKZ1EGvlw8HqTzEZq6qbEEy1Tr
3/bcyaHSnHeaOW13EJ40P9mQY8PxTVERo/2k9dC85BBlxV6prpnnoKRiy5kQFEaANAyLyKCV5HI1
emnwkJhGxN6ic4WVeBF4nV25rO0WNFxaxnyF8I5XWkA5K1DaSduyn1EPMa+2aWgLfDRUQvaBTTHb
t9FcQhvMoSgyS1+wn/yPQOzazl0ZE1+wiMbfV/yjaFCeTIaG7NGcChoVQrBgdjnMW8ETTPW4qwAH
A7Bfr19+YDOjGo+rKEfm5ebG5QeB08x0LcHjioL0F6zkjd2ihrgXnrdJt7fRDPuNVtiu6W1M1iZY
IcaicTtgFRY6+KW8IPP2H+A+Gj/HuIeGLDI57/e28hyUHKIRV4Yr3PfSEk44LGUMlF9dJWnbDJo8
9zKWcJi7t55GdusO3tZKzTmoitY/n4ixo0PerJO22NtXSNm1x/mAFfpqYgw8J9ff0/w99gwKRFbR
xvR32dzfKkbveAmDChqZkC7ORWCb3JrE5PZdKSMYtHVmZVbiRysCtrHpUPKcuQJ+jVlmKL0GqO6Y
u4/UcsxqvxhDqX0kDGrQLKC2K/FtECWZWwqM5qPe8tJLYq7EimkncfTpgqDzb9rUPiG+o1cG7C57
oOdHK7BymU/l8g0T0/nTsmQLoAIq+wI0pIGMiXTpE5UrTKbZF7QB7JeU1GXHIk62SFjwKXTBiBnL
rhYCufafNa0owyLtLJ6oibJNUkXF++ex408DZJ6XW9Os7V0O/aahjUMxDJJbVuNsjxNlvaCxgvBC
M5izoA/ktqjCwkOIS+YX+8oT9goY1mEKO4sURAt7g64wntRMMGqr1CES9CIiIVIhhlv42zF2hfxX
OV60MzsJ1jCGdSXtJf9AGqn/WLYKWh8CCcxibGZ1/6hVUK0FqZ+AEn3I9iamOqOtAAkdGS77RPwZ
wK+RX2dy2rcEv7i4FaaMipigyagc0clLsh94IstwEjnVexdF4HrEGNSDF1mmQELLY8np94WMtb+S
m2XQ53kPa3YS9LO1YEJJygPMUCpvwBn/eogLP4E2DY2wQeAlHJa9yygGKK8y36ta/Dh+Hv4WIjeZ
qL86P6xQ95hdl+MnnA6wcyyuUmvux9Th4DVPHfE2hFPLXI5Bxt+jBQlkK9yFJKQeVHkqb7gw0LCz
AC6+5JTz9QfwzOWqbbqiS+/1aj6Xyov+lgDAX3E+i6i0NyRB96YlhTR4Mh6iNljEy7K32Y3Tffwk
mDaZ8pt6L63O5X881fswPljKbOLSwXIHj91kmBYkyYLeP8EMaH+urs/B+Fq323/I+U5yWJIBXbby
DonjRLjR0pOjNEmO7iuvWMkRC7jnh1RzjXsx25Nz7Akf4ygCFnNeAxaLfj5DRuFIIIvXDS69gtBq
JsaxUBN7MO4tfYnETc1envarznELkz40Py87t82g2dt6SLzAz8kpxwNzfbRR7vyqiLbRW6lVoqWs
WnqDTpmEr4yolvu6fkTlHn3IpKnSSzI1gwTqrFymKNPwFzTh52Mx9hAJ7kdpZ3A4lSuU6WnAbZxV
uvK8DaXONx6ol/nAp9e+zMO1CxSp23IMNnNEsXYH9bN03r0vsZg3ZJeX+AT9KRtlotQSyLDFBg5w
IJLR9/i0rqt6En00p1uxkTu7v34bVZ5STlmeYM2zmVK8FeFLvGyR9CRK58zDrhMFr3xZnq6kjRRP
OXEM10z06ReoHjz9pbVWNstInhCq6uTMFpGZ+xORGHuGoktbssexVWDeZgKuICla0j9cZ2hlVR+6
6iokjspjr+KKt7SlciY5MsyHIzDD4qY8h8eKUBplnCIRV61kt8I0iJe23ea3WeKyX3ZYJTe64Z+4
EYzVMm53mlLjRpFjS5MOsN3CTLWe9S/J/Y0cp6fvuqxc9ZVSsLVr9qjRWnl4qgZUUNb3GeVxzS1L
XecNXjKGhzN6gL5eQcJBTPnwPVnj/++9zzxNdd4kt141Q3K6GZSWTHZnlK9qI9X8jaZVjHR5V7T9
nWKYn8vB1iMOwPex5Za07iSmI5j+ieqcowsSRWpNedrVvKG5jtR8fm+r0Iq3Ep0qOQBY2PbEZPj1
Hv3w2c2E8sIYatRAqF6oaDaLOPfvuZsGpa3E9CQaB14q554szpRLGQ2Mud6Cc3Xw3FXqWFls2C8l
jDpCZo/W4GGR/M49Gc7+4ZeBmzN2HjK9h37EMtzFVkdEjfKvVYFi18fs/983/z74AMZc0+8C6wxf
xTrg+4Rmuj+4iW5vrVXCtSnjKZHr4ClZPA5jfK9HYbPoF4yv+PqINX4PTzbKze9S8O3YZvf9N3GG
jogoi/MfrCxOU2STCqQuGpp0Z5qPe65T+Jr3HstUn5cQNiIaZgaXJ57f9UbOGe1SMJym7TfzTMO+
pz3bb3WENJu13S7NHR+srNlI4m/812YXCaoZzFjex8diQIR1k+yFRDvnHwHUCkYFZsxDvNHYuqp1
kYkbXDG6RDh5SkTCpxm7B/rKI+RYA/lVefw9eBGr1ZaKZIj2ygObdoB8fhtAM8kn6PXyvgH+5998
dlwJ2JaI5SjWPZgamQ6/JJa7ulIwomsfAGb8hlYVrzIzD+kfwh844A9Oxxsz2oA1s8YABSEfmb51
0dP4suAdTQ5wdn3pPzDh/0CbADmCoHAdXR4q3qNvzk3URf98fcgO/PEPwVp5wRHE3s2yYrqY0nr1
5Z32zfhsGbXAfLdQkHlWnvJi7Yo45bVlpvN+ZZSlHQvq2w9dDTovAm7mDm5M+zptJ7D+JHCJYD/u
0ueZ7rzLYjujNokhU0YkCXAdNceBHjzCh8LFs1ijkxVGmX0SB3dSDElc4Pqf9KCMJgzs6CpSuNMP
+KZwC9wnMXUMO1ZioIl41UZu4N493JXFZJK9RInUgunzCxL7yKvPfk8+VXvC7wt0Xdm/322UrHcP
HmrID4CNBrFSqJ5XOgD4kkFQB8j2fLEvQF0q1ZdTAGJlct0oFgMvXZdjKhU6l8s8K96+uOnB/yul
jg/5AnF3IAvW9rWBl6WhG73gmiYxUqGIEqNRL///C5ftrMiYfEKJI2VMDc36gMQkBJqkWnb3o2iw
gQiPByuYfOv+XjK7wce0DW9IhMTUE4AJaAo4NslJlRj9Rf1atqVwzgRyk8LQTHLHKUOgI8UmgzXd
W/Z+io2YxTDqmy+3tOk7+NlBz9eCvTfoHjuXmWWmXa6eJCYucIBpAiEmiHmT4wfCk6sDhg/g7JqU
HKRHGRSYVqx93cFEp2REK6lwEbatPo/tN52KEao5W3R4mw6tTp3IHcnHsZa8yolOpGwf9HZHQ41+
jdpHlXiMEFjgMWgKCagXUUEfoofebdBMytK6qfGngoN2A3pMCQzuAvtk4JfvdVbjZ4VsiZMddMd6
PWwL5zARYnWPJ5wzfKgADO//igqJUJfTbK1j/jNEAOZZRgTrz+7EsnT0eb/bmJAcDUL9+N/8Qpg6
JX+aTJMqsK+u6+7rgvIesXm+e/d+pmRjrM6Bi38/8V6wMobSnkdOeIj//LDCMUuws5jxgVxRCH9E
NPZgZvAu67pfBVIw2WeU0J/k+2hKU/kTUnDql4BepeL7Zwjb57WzbftD3GYRcQpSza9PTvYefcrr
ZFii0/jwSkOyT3YrOiaSLasau0VcGh1Z8FQz6BH5q09P/0zRN7W3LVifoX/GqEcDaj1vKnlPA2xt
clU3fD9Ps6mgqGpAQ+uLuPWH/rXr53K9rdVZkvH0Lgh8MIuYPimp9EXOMSNq/E5uTTYXMYvBkaOU
aAy19ckumfpvPWO46UZ6qlh4vOvJdGYkbm/atTSfMpZeDfQTG5fYB2FBA9Gh7AQk1SP2t8m552xS
kfixPf6bMB9wWoOlPBjtwmiaSCM1pjkxtyBtVp26/yScFhR6SRRiOa+t0aCa7d/JEKtO9T14hXKA
fP0Hew0iShAmDQW1sRXfmlDuNEBU/2tORGgPHVxwp8JPzXsmvGSjoxveyKbQtIsC2W2qTfnIMp/a
0S6VOxeIzOVd8Jg/s50QvSOb7HIlEfbRfk2s1AO0D0Hgwg5QdiVEn5giyukjeTCAeFAistePA0yK
LLFPec+Iwe0mkMFHvIDzOSjztt0F+AZ/HIJsPFuh9UFpJOxQscIzUEUaD2ayFtrGd3pqXyMJi96e
2wXRjl3HvrjuFNtbegWPVPEaCZtP1usxqBhlX8y0mxlH0JEHcLkWFVxU0vOMMjbZPstuI9je+UP/
kHtYGfPzD+KVKo0T+f+CmqsiPWz4Wra3j3DD2vXIai370pxfas6JdCbFZKI7R+2oxkGVn2ry1bNy
3uBGGjfCdPVKJ82HlfYBQw0QNme8gVCYhuaUjDeG96yqVLGu3tKYnkZML5fObXZIC7b2gu8B7b1Q
/XQREFuWz1YEW4l+JIibqubAe710KIRTw/ockxKJkGMj6JjOg/uUByKSXDkkpiZUMWTsba/r+PEs
ZeEI1rOq8AGsL/Lg9w1dsz0bcyIKlDJH2pC78EQPjTNPNlMutJwULglE2Z9caXTYeFDGRKPCvFPU
kXkEY1HMew3FECZxV84VqmmP0ReqytZZ3HGg0iieP4vOGq1U1Cq4QLbFqaYIFxtOpkjWno+ZKT/W
AkmthTrtYkr9CT4JP/WvKHSObizlM6sjsaBs4m3LfcA07vnaejzvkSVXxcEY7ymE4Q+TwcqfsA5U
AhodGHEiGS/11hNFU436blfqQtVuxVKuEoprNTyXduEBXnp1rH/JzuKY8BNxkJI9aUBnJ2w6Wer0
JWKjomKT63QKlRJXXGSmCPoJ8NuPD1M7RQC+pSfSp5C9ZehTFmOwOIXZM84qxNb2lwRmE6ZEjgIu
8nmPeVBSjd28gubyj1JC4sSAJ7FmSn5X390vvYZdJKRJ0XvhFXDI9HBouVgf+V7haiXbVRX0BmmM
PeDpuXjrBtAynEExn5x/XZ36REo6v4S+7NgpBtqvbBYWQgGH5rz42zfar6+HJhRrxS+Yb0cieDVs
zxcMOtqhYDKEb9quSssz1LvzrmHbQugMQgZtK8v+4CzsEbvpvLM7JCBC07bZ+wPgtIjH9r2ja160
q/l+blWMlmCUKwNfS1pVYQNiMuEU75djXYK3pvNW+/rQZ9VRnEDvzdyqQTY/B9Pug/lRr/YM+ZmF
uw6lBXGceq7mjRsep49OU6VFwT+V/FbsYyOEIpOOMziBfEy2F4Nv4ysPgGkbtrxsUymAb7rLbq18
kgwiWqR7NSbkn6hEu52m6kdnQ6lblia6MuQbOtFnzSshAmcYLyW0cb5YKC7L8UJ6aSLP4nuOnzW0
aso30Q62ERaA+OY6KNcGT3xz/VTHIiiKecJKXi6HM/g7rJKrQTvmve9UuHp9Iq1sgoMMYrU5pz/Q
MNLHZBJ4QjHFypbQkB/O2Mgth4lDP6n5K8Yrs1uck1q+6fRjQ/VFNQ90Ph2T4TjeBZytutU4NbLX
kqgkLq4Z4gCskghjEvGVh3I4jxUwOhz6vTGG7bm3lMtU+OFlNkFQi6DWh84OlZ+HLvSBpYoQUfTV
BVBoZVzrxokCtfr3AgHrmnwQmGttjxXnNcbtNmJ+X/PcuKCEyydZg+cPBTtvHr930EEQVzjQkUhh
VTF4J1E7kRD4Tw0K8tOodF+cJWdWTlQ+NiUOeLj/A80KB9nSJnX2STvpDnj4NDVliVRjqwsPmWbv
AIgK/LnPn0V4UlRvNvTLnwLxWjKtJuqRRpD6KcupFyyHuaIAy5Yxcc4ALhyowyZ2zHFRmuvqy5PV
Faap80ts+YdZlWT0NQGsoP4eCUgmmMUGu9jLPJfbhGJr47NkEqGjC19LLTq6AEsKg2ypWbB65O6p
75cvh2k4nL9RAmcR4m4mOf4F0+eyIeK64FwBih2xQJkQJKjX9IvF9jhyZuSZ6FjwgrRVAiB9PMbf
4RZn4/OQnyO0UMUfWvQcQlnKRzwH9TDW0VX+Pm6DN1kICzbWslz7eY0CEfI2H1+1A7SUOic9fMR0
JxfKqI8RzDvzAdL5QFDcxRwPDfWXFyGJroGRrXzH0LRa60lF3Lj+N92U4wG0YEiFG6GNez7paXZv
5x9pqM1vcd1C/Et0JJ41yM0R4MBIs8l33UcpXR3VjSSM6eXslxjoFgS7od0s27vvYPV7c/+kqHHi
tEiIyDJNA5HdEXcQampVXMpQ/EUVWIEIl/BUV0Ki1y1TVKxT+ejzWhVzCmsyTBlzXCGw+uYtUF9M
2bMU6Sw9BWcqgo5ljQgLBjqm5w6Lwr7ZuWjfk5VU+rKBbI4wMYWnrYdLlqVy2qHNZ3Hq7CvCmjR2
WEZYnL/3iJgwKZcu6j7kWHu7Kwpetyl/Hh6SErjF9DitJqCYXt8rxmoYzURyTC1nQxLP410hul5M
yOk30C2FykxqvZYudN/rPWKnC6YkQEXlr0YnEBzA++BevGBRD+bA4XfFHqpKbymiW9cOAB+eCbMH
awKzTjM/+NpqgFItN3kJz7u6zeUv3wrRu4q6h4o/uJ6xC1qJN0sS3SXLn2nrrutlKPHEvxdsJCFU
i/PE7qBkyWJFEn0g6a9LcPC5PY2hOe/ZqkdUpyUiaRjBQvN04tIK0Hfqn+xtdfnA9o3W1FSwEdO2
8DbOLzjOiE7dz6nLnhsljCLmuDIVq9lHoc7aH0YA3jWWAyrr/5uQAfVNRLQJo7qamlOTKCr2vpI3
UrJQSaJstwdlkFJr33WV8GYCHIoGKUbbhAcXnnJjVrgMBQDiAxxQRvvSzKv0S2IzNKugZtkyffyj
c5aON2faOBmFfZCzRv0js1DEIvToY44NkDKXv1I1Mv09GRsk0ObBKjOSmfUAfVNxaregb9U+/gke
DjYLzYqlCDzuxj9paqvObnFjQCKcPWgxoOCz47srM86C4t+zE2WGgudKAmgNKKz5OtehulS723/3
c/bCwo1aQFy9WXtoptKOXO7NEB1kyJoeuPPoVw9EkNYMRSR+iMvas3cvWiHMQ7CIFMiEoc4D/w3J
eXoxdwSoABL1TU967CPwpWIjFVSWraMjh+QcbVfbeyNpRN8qouHpXX8k1rIGEEZSR/PpoyrLxLgJ
ncChHdvqn0hw2zlFel0Rw93q5coA1rDRA0nrGKba0ONeFS2RKOIwJ6ZXGQqzGiqXmTZzsSior8X9
x/8Wz1gGWpGYc8dTXRsUPqaRw37xlG+HqFdlWcIyY5CJTUWZ3wWd1lk02QtpJc6UFSwGVZOXrCjK
XBZGIf7FQ0Vpar/hEcvtx74zyLnw7nFFu5xDMgtBDg7mu8F0Lo2gMpXM5K/exehHfLStwoeWWLW0
5wSXRR01kj/dsuaCxpgEECioLlVi5qZ2V1okU1m8MhTsT7skAk3O48CG3QxOimx21Y5n3eapiuk4
LFxz0dJ3Aq8qLIAMXtDwNALtM3PZNGDgkw/GpL/+YB1pOZTdaXDUG9MGeTGpxhYcdcUzw6V2yPJw
g98q5Fz/O/rtA19zYhQAlpLNrCiStlRtBIjq4k49xPZe6oCMQ1e0fFOHIKErNl0SkBZ4tItOUfxS
3RAdL0d4QGj3VTaQym52sEFxtE2oxrVCMDmlMyryKglRcS7Nq46o7QqLkeMLJOwp6O55zm2dFRLB
pibBSKANZee/cVcs8arCYQyEVIp0eThcJwUiqrTcZdkuBcwARUaGNwZPey5nC1z28ZCCNHPZTyCE
eCS5Zvzjp5hWKwgzk7hNl3TtRgKPmoVY6UW4EOZTT8bfoX79Fxyl1FD2CYg2iT0Ly+YPnx947QLE
9EKesiPbEuTNVGOrz5kODxJhSbTxYNJylzZ0N0wkmQSthu9MfYimnuTMuybXUPSdvf9iV3oULWAf
5d7F4VZALJCs5iy6liyI2fDqGqrzrKGCuaGAbeGDObCrg/gvAbNswCQOgPv5ZclqXUnsY8b9s9R5
hT4D6ZMpzKqspUuCgGqp81qFTygfrvdjE6ZyMmy6exzJiITHAD+T+2vPEIItUIODxoIgJxbxd31X
7QZPA8XbS2TSCDzibG8dAhHs0qChhg4GnSQVn+ISqLlyUSUs7eBEXaqdct6sWmMJrx1fvRlnzR2b
okFtef1ZayjF882kKSV4h9CnSyM4OScDm3FuAQtMm2P9bQzSG3GmOIFjIPpvr6UrNRHPpE9rqb8K
zC6e4WI86W4H/Go8fvfYHtICK9sA5XvlFIAPfdGGsqUfMvmq2dC0Q4kNig1GldLS8yUGXxvNXvWp
UMe1Xghm97Qn1QDb4CeHT9WEPTlbczf02tN7aurh3FT1J7+7/RaEdHQ8rxiRDW/zmXXm9urdaoHX
hHtqiYE2xpL0blt16DCevcfTeWBqZjZvY6RsYCQtTJVk2URHGOjolYpCzoVyf6Z51QAJHCUIHPoc
bZdOJLP26gkBW8pz8kYF2QK3ntbb3YxSCxiBHS/qZ2TO+sEAVYIt1tKBgssijiei+nRhN4bZcxVp
6VfmhEpJOnHpQiqni5J1V1shybh4Mn+xQehgpO/MseMXwFYNqedZtvYp6ZA8Cd1iK/Tm8k5s3D6S
nMGxN5Hld7Ii2lRzmiNNlO6lr7Dcc1TUarhYG+WGOhBHAnb/gRrzdv6GuhxwNuzXHqJTj34wv7h3
WOoq207KgGYcMCn+L73AZAIQc1SnhG2bmu5LZSdwo0QZeqFMlGTYgA8mTfWdQq1SlX9O/nGgLVbH
Yqzy0l6yrnCk4rslQG/EkXg3TlbWG+wsCn1Wqy8B90ZvskFEXwVTcf/Qy6HhaNFg6XrnVnwiNJtI
/pdE/MgZBehsi4+SwtJ19GdL+vY/XjrZ+wwcTehkjHBG7aViO4v+bh8MmQBFzG0kwX6iL9R4FP2q
PIvEf7Mr49EfitvV15fLufgVns30G+C+ZPoSAhtAxxiQHn1tOI3SVtdkvylKFMpM8OnSff/I8J/7
2Oq1Wm7RQBtQT5Vdn46xm1ip2FAN4Gnj52V+VY20GvAbzG1xXOQ6UxyrZCYDhV421li3rbwLYtpW
Pb4PuGtnBFfgT2H0Ak1pMTJzaGrd2m/XAlwh+uwgVyiY2bmikgGEG3u6q6ASgiYMGXdGLmGikacJ
kz+42jctc1s7XKjD6PywNxRs04CdNdTL+WeJLggE+RwpMwgqnJt/dih99yggPpGZdvLTFT1TvvLD
N/iJReRWAzK6TcowbkIHMV95bJ7rE5Gt4ecaw4tDd4k/hEqDr34keat/AL6FY4MkHcsfKIMVNkWg
OgdBZfYYQW6t+4boTRp7SVnA6XxBeBM0bmcN3e4hsAZf5xzwjH+FxZhcNJxSYz6q3wZE+ddN3h8d
ge30HFpU7fsMMngCTLBmNunEEcJykSp0hfpp15P4pu7+xygwgAqHSpIW++hJMdaXhJigjXTqr8fC
doMrycMVLeTVEGOKe+wu9hj3rWs404SWW7tfkghQQstmRwhOuDoDauczb24Lgn1/AoThqYkI3m3W
6ee+ZL3QpYPnM7z9zzuEOcNdNtx5w9jEAbXknQZpQcZWSglySgdXiZPE3tOJMHwwc19scP/JEz5u
artIBZI9g2k3CWdeN77chvG7YYNZQxy+TWpBSSwiVJUZDalI3wDUjKgwGKehCI1uU3MdFZGK1ubc
HwOgLyXftEaFOphFHUANblxJ+OJR+Bce5f6muwCaVhsSuDOlLAS+gWHg5+/lmU5Q4qQql32pgL3X
/976fq7YRJgC7GY0Xwzj2buJsP7DyWqxgjn6Jk22CQPDOjqKl9v0N/OFp5pzFEqqmZib+GpI2q7q
XoBWGQtZwYdG7Z2XPwAnY35xLR0JBQ7vCJfNkjg6oNldESPDcJL0n6TE03qpwOdihw2ABQ/G6Jh3
bz9anVg3LSevqNLGYhx4wwWUrDJ87d3/XzvpPLuFg8bO/kBNZ38rjp/Uisyu0PtMNxrCmM3tCxWZ
Hnd7YS0B8II9Xpl3ZoAvu15/msVZBz8qkVGXzQaj5075W20VABrvo0YRIfpWmeaoo57YIXUPXtBW
291JEYbHCLqRNKHt266y5KMHKjpiRl6k5ofqapBsztMcW+hukB9QenNq9Uz2cp38k+8zgWVdmFgt
46+Pe2IutfOKDsyJV4HKGmB9VoweWeYE/7mCusXQbq6a/Kse9Nc6cys+LrBLNxV5GqoR+UOA0BAL
ma0u9YrctnP3Uu48lbWNG2xLImEIosJI+1z+0uNcrrYIp0P7IYTa9+P7zFjxJs7CZrHYVJI5xmdq
OGnwLluleZGSg8LlG9MEjjga86I5L3kfx3Fi2uKm6Aq4Km6OH5giKzXGpUdxNwum8A+Rbsy/Ivev
7o4pbdXdIzQ345s3Lk2HBcTPCjh+xah0h6GgJGVqsGM/wWY6wX+yVFh/8rdFTKogRTzdE9OAMYSg
1zZPSIIfUlUfGFwpjOwh5Dpbzss7OeVJ39Rmqd/V9mggOvtf1U3qDJUAsO+vZcaKekck6t0UNHeV
zC7Yc8pv1X706RCyUAdE0HLfsaElcxso/zy2cv5EptaAN3x6PRnqk31V7bCVg01DYRsm7L+xERsb
UcrUamI8KZsh5rNSC4ewXGZX/48JXid06AttY3L0hKNktzyYPBXx8uLekfgWnnkQguX6rAwMqHbB
BJhU7eK6JLchSxXa6RiHBEyMzwvT24xfgwPf3sF6vUl+tULhFrI+RHZmz7sjpdZYxkNApFUk4rhk
vqLUXd0jJouhp6ULKSTRSejEUZ8WsyGAKlm8Q6u8i2m1Z5qLGlXlWTl0OHHBXOM2GgZjbFG8AXXt
vSoe+PMPfncvn1HSxGcelSrvj5XYFmxuFUPCUzHmWyE9ITC5HwmKOFwTEAOc/HXLLAkhO04xerug
+4O+JViDNxmg24PJlHGbeU4TBQ2WYvOrlOsLQq8g0G0wakZj9gedzzV94+zWKDUa31k7QXUTFN/g
XM/M6/CuI3b5qHdOhPETRXO9m4W3Yl0axSohg9YgRhXcegNp9CjQgBUE2ZyAKW4ZTVtDT6SJMFvB
2Yac71zw2eA473OnndnPQGL7JPeuS44NxYdZTx/+VkxA15sHByxnpzDidY5w4NMFRfXfl+gU4DTT
vqXYw77AzM/i6QrfJnKtPKOJPymmnJJn/1ibqF+MRsPuMLxcB9KMN7KDWkMN3I5clhEpEeM4Vw8M
LPyNKgafojZx+eOCVbCgtnmKYgHPjmxO9IwkOBaSGlVOJWYL3N5ucQPUtY+5QBEIfIciBnYH2rQx
q2POb2YK/IeRk3LzrVtr9lXcfwaZTBL1TWXPVYlSSOONcIRTo4nmgjNTq4kfajO1QufUeYy5EQLN
T4zaZCNXnPDl1nZK+w1Pwvh5L1Z9W202kHC+1WNyPl8OC9db5F+J/KN85/yFmLXpVA3j985KlDXV
rvVEwFsC8NaaJxr8XeiyXDOnm5Q2/RooDgUiJUKmjq5+ZZXcSldg12Egu2qgWOipIkBMqUu7otwN
sh2HhfKFbeF2pIvOjfBS1UtVuVu6/QFG/zkWjRK9s1yJn1CyVHQu0DTfTjlwMVSSQme5Z7ejCVUC
9yga/4Walo/6OpnWXCRlA4op1RTEK7xgG/WxZJYJY59PL5V/X+jhs4Yhr5MPG/X6MejhtT5QEnLr
LfrCtmheBr7eeTuYFI8vnbE0yxbOLpNORo2NkO0RRVrYKEUx8cAN4jiz58m1IzSy1JrBuIqWoguH
UVggDWAqT1iq8TadTe3x5hrqlK5ysaU2vfbAipb/70G71myt4uIM9jXeiEv0nQwWn0eyo4LKNhx5
OtzyJdyAvY/QK+gL0sUr14/ha9IdI1fj/XGYKiJA8gk56HH1SoSqde539IIXpARcL9sjfcGBOz0P
nCoLDauBXf1BQtqou+abjzIg5Rnqm6eBC+sxzq+kvCMCdxaAuYaHaFxwREejYxUxLb4mcdEnvAQa
lUtmDyqqNGobptebZ4U9lt5uveQ++JKvRal/X56+NX3FgmhTDN2sHKZo+PK8S1whF59zap0GT6JS
NV7guXC+wCiNmKQsw1Y7ZjjL2znDY0a9ItC9gqRGsOMke1vM94fo+FbAuhvHqOaiZpkbXalabBBj
u18BMCEDg6igbZ4rFY3l0NOVtzpARnX2Nob7ewdTS4rSYKXEpBIuQVVfSxI4VF7G6xsAZeo8nPfL
GmI+mHYLzI6LSLznFIiEva0/sbs/s6qHQEIsAQ9J/3HJsHOJvuE/v0+BPYfcnUUpzHE8MS/gMu2G
TR5yI+BAROWavpGO9QuUDUk3wuiWBE7Pz4COxhZT/BCJgU2+Hh5jrjELalEELo0FlKgqr/xak7A/
fAHTN/tItW3zNk4lzSkVh4PwvErtVypE3ei3DvSXUTzLTOPYiQ1TJSFi7CCCF7vJAR2hK1hKec4B
t26jyuKJ+o0wbEwueiypX92XWIFRm9aFUuGL3Q1CO87fl8eTvtRAxkC7CbpNp2fh3iloMX/v0h2Q
yNknlzE5e+2GE3p499R23QV40D2T7xwrioGBXiS7kLivkzJglJ024/OlxTftZnblCdTNdtcilryO
lJ8Z7s5av2Br8sOu/231aEnWmCFNe3OsGpE23luYxSlLbwMWaWcPJJG/KwY4bwtiDudHPoLnYvgP
+1uKUSDNipdG2ocr6Ip5SPWQQaLAPvnC/oleNmUONkMNZhATiRIpNYaaxB0pBSma74eVx+FFf/wn
PKIjPVk68lAOFXMePxoeoWj197vmIUQXC94f599KQ48TlNxfR8e+ckwdY0vRDseBfOcXsKOTBuAN
5VD8xmVzQNbwg+pjRF0Ss9vh+qYFg4MVjcMrQit8AE1XgHUhRpDODzP7GWbZaHNbb5XkMmgpZmOP
3eRPWCyy3aGsXkTpm7XEsx/UiReVNfxkQQlL/tnCWqzzPCt54ak+wfdgEJoe8tBSMeUtER0O2yff
6/LVkSN3kMafulsIIdCrL4S069Daq675lR6lTyp7BvAlhT50O1//UR0dOC0rZJkPkrQCjcMDuISf
OxoUkb7nv3Hl+KsAKnEQvQIxjYzioTZEASIEs1hUX2hmfLQQJEDGWH/85pYh32rMdH5hP1Zh8H05
nAIR5yocqyVvz9vpEcV6FsH9YVElbEg3ikEVQrhO14vG76hZlgKSB4vRu7nSMmsJ6LgWNk0A4T0U
u+pzBW1nTGgQivLKZUMGC1d+h/3t3cRjT+xDgtyPilNYtARSaLOXExJGWv1w2LcNWNiiKpVKyblt
P67Vog+JxjRlMcYiQ95qYGujHz6WQWxMjmVUEx7BOZ1f7gRTUG20HvH8IJ/v0+Qw0cmrtXO4F/AG
FaIFWN3g4TzjZ9VCIeUj0UH4KkbtKg/hIQoX++UXxGjAN40gUi6xvFDNpS9/PeF6suI7qxp2Xgtc
471qu9z+qUf5U2YFuOiSMwaCLMy7lNCA5exUbIjCPyvOyhJVBzfqcdOvpnDcXc5PhmSgU94j0jjl
Su4mMSciVVXfM6YOXs6WvKcWXav8ZZRY1Er94kpwWJeGhGf7+2e+PA95NrTu3AWM+U4VAKiVOvPO
GVbvu4oFb+wgi0FwDMVB5Jk06Cg89sA6/l4lRGPWNoXSkiyQEzpPk/TLWVwz3k8EjidA9s/B7FUl
UEiIoPbmsBQCgdDBtRSVHO1oq6g/GDDY/MSGmvrmuZ7Qkt4YAKyQxD9Noo6UzfgLycwB82TWGQ3/
N/nvdoH21mgVPDtGdPaMyO+pX9QVhJRplXy2+wbmB1FwS+CmAngNZ08HfLoKDIxhvQ0qnJM1wnNm
8CL1oFRp6yG7xj/1EYqlnLbDlX4LJDyaFXhytNOu1bTF39omGC3Ew5aH8U/9O8Jq/lt+Wlq8TMT9
JQ1gGq072H6enui6zCgGTDkMitIZTZxR2voBdA293GdRtk4Y3hYKJivWuAJTC1r6rDEXd2Kv9rcE
gmggHb2XGFxJjyh4KOBwu4vLFXJX6hHjM9ury7Tsidr3OEt+sZi7/MEgWx5A+JCnPwD+AaRwqVht
cWkSb02iozf7WiXUbSgmy5fwyoNZZX8fKU197JDNUwjGnTOhQUFU8Jf1VGlei3R0EhtGplqNEWxz
KLBdvHQ5Cn8J7RTSLuH0ruJMzS8fr/sRiYL9NjC7kwCv9px8Co/wiDEYgymLHrUCICP1SaBS2Kjz
9qXpLFHO6PHDiomsdxEH4/JnJLIuhPl/f6O+V9YVx+BziyU+G4OX1QBdJMFwk8793DQZZYcujqsa
3IDS0s+h1jZ6B6gDCG3dOzWnPtdpFdAZUpOkRIyJJsL62GbLMKIcDyYvhZXk26BhFDNfwN8GbpvW
VFTNzyantQEhFBJ1cyyWxIB6MFfUZM/zI9W6CioHmkKa9i81mXnJJbyKXFisyGvY7HLwXflOqjBR
v4oqo3vc9ermdzqRimQ/SZj0beCW43SIh5Kwn36SQgcoT3XNJKvXRPn4mjUGcf/yoEZzL/1Tcl/y
wsPY5u9a8B9xGUNK4riHkUEckewXi1rP7aeQPeRtltZ6ZRnwqkbbUqUnwWCXSKe1cvz1HKr0FsZS
7o7JW2j8oSM8YzegAmS2pJxgkrFV7T12imiebR2gGFTvhgXNcLjQknBM5yiuig9ovfkGJqtC5BPD
2/m/5/Pc4pT4HcJSK4k/Hlr67FFNb16B/YB5eMtwWcgy+NyPXjNvVqPjoADoHgbtJB2+rhyaTmmh
vp0aUNztFv5ff8PyoKD/YJ+gLi9y68xxki34Ej9DzX3s5uF6B8fOAaOIAkKbGp3nJ5xIwZLavhdM
MgDiBCj+0cewBKMDPV1ZbaUk4rExhuFtIqdbynuoLC70MFjQ3Bm+3FmDQUs9c9iryU6oDQMePDjR
WXMdYojYB0DP1PZFmAQOlFyufS5Tj6U6oWztLoJIBwaT6lgy4gyq7goerU7/i5LCGhrge4lwgYIl
7oJVMG8drSk3s8xziZnCuywpDeaDwLsq7RPCDb8bJTu2POxlsEiUJp+vRzVpL4GgP+s9zYv0uyiz
ars6dW2JByJIkjs2o3mf8COlKLHw7S92c5LT/i4JvkY8WhwIPbko+0GvJeFwxMug/OXqp/myvVVq
TFAYcnuyvb/FfBlrbSlnCm7tiU9ZGpa4evpI7z43/+UJtHrIQOwrl22T1G2mqY3+q3T/7CkMnOnO
OTOEuEuf1cM9I/0pMZMqfu5bNMIIUy2RreNfCsy3N7bTy7azZLWoRBxtKihSF4P0l0kn8WPWXqkO
bmoQX5gHz75f0w4bDcAkc9AuSG9aODdiHyMuO0DjiRDP7LiugFA+KjIcBGaxZ681Hi8KnANTpxI6
0UZ0TVxAAilAYaY6QliO8nx4n1iqv5F6B57z2RggWu3sSL98rYLc2a9tvDl2JNwy4GHux74P+qk/
VOA65G41j/oe/mnt4tsKgy3xY51rogojxcxRDhiClm4kUmKfytw0Fei37S9pGaIcIYW9Vzd9YrXd
HXNhGL1UXX9qhUYzyFmzWVF1EPgxOQlIpbqS2dbHwEHifQdVFZEv8sbSa8RXwGF6p9BIA7HH3bdv
RK3F25lb3NhNeTNF5YU1/Hmg2U8M6fEsaCAATQkxKqxsyhioGQKzdLUu5EEFzK05kOLYJkeMVEzG
P11MsdNyXq2r5iWhOEt6GH6pHA/2pyb1FWLrVkdR9yI/hBpJVitaqP/xHfIWOenIJQeITKYCYatO
gxoL147bt4W0AtYroJRnS3PQcEgAxXLq3X+FKDYmUhiW1HvxdHb66gsnF7el/xctFS6wLAJArknc
0A42PiIxW7DKsfnDs2jWyjcBeO6mPMHndrwKGfmVKcM+BZXizjldR2uan2QXfIOVNXBYYeq39q4J
cLOx7x7dpcPlSPCJq2Jo+ST63hPaTizVX5dCP90/LyPY/LcZWcsFEp9s4ZDYZhigK4OkkXsnlQYe
+o7s++jA27yKb7ibGqp+Rny3EKjTNLzBxPVczc3V5yOQ95rLtVDuRvxMS5yJa5mTbSOvvHOP/k4E
MADRbsTgPZxU1DPDpCcPUqr6bAOY3o32lH408/t8wnYvrzVsolcmauhZ7wkqGhPUkeOl40pmfaFL
yQxL60lEDHLrt23P+1cRadHKzi5fQWgAadvyLpx9JUL4YqjMlRAwxLG99CUoqEmLA3YfW7Os2TTn
8YvCWtbzHH4rnNbG6iQRL+c6E9CANPZHSJ4V00GAVEqcRB8RDhz3Cw2c+Gf2HjLsXULC7Ltfsi9E
2xeHk0nIATZGKpwirxwUyF0EkWozyutjmUQW1xdr4Nw4FR8DHa1x3Y0NHrCDHWCGbd4ZJKgMroKP
badqN2xBqMp+Bz2N5g6eOtBiHI1yyj2dzaKxsttZfcybQLT65HDLaiEVSGh5be3pyut452Q78Tt/
Pf6FwG7xY6hSCMrDWOBeopQTQSEjZ59PemeTGQS4bHnkWs+cDvbxINoo2Kjn0wWWIF8PHaTEIZrk
tDRVXtRX36YxWnJpLSBFzEnLYUNMjU12b+1L+C0ESDdEc4aN4xqOzb5tvwj5V7kh65P85Fqi4e3b
CiSgJcGTd12sl6+Z/SbNGrul9nhwCjBlvfAtjrkzsJ442mNWzdt5I93aIjwKZGF33gBiYphDr6uB
8lWbjVtwkK9wF/mD7pjwygSmZ4I3BOZlU4TBrrORCT/p8al80Vkaweh7bLJHAPlb1wLqL/HsTxh9
/GDqKyiSricCzLusMRx8Lv54fwaHRY55+0zlR0TXm/Y3nu5n64VJsgtJLB/lQGrXtf6X6doLi3sv
FTNmL9qjRHRUokVfuqNyyq0/rGYiq0DDl7uJr26WGQMMQ2vsgRJ3ygWaFB1l70hNgDv28hDFxPF3
eMG61ooiNzJtD0FtieeubXzZF9fE/0ckHfvvdt7t/iMo2juuShPqLEVE/UNun3EehAaXi12RkIqn
sYSYUgmjn7D4u0MQOQ00XTopQvzJVb7PgvnpSULR0X5/tDZ+FrhCMBSwWIurlu1cLdtQ+mcgAdWQ
qz8RaIAKJ32xiumyHW7nFAFSNpQsjOOFtAKkjPzAMtrySv2EtQxOHSyTC43BUAsjTFlr9d7MAY8p
/rgaQ2ffwkz3a9GJ+K8mKjX2Zb72DJHoLDcCZdBFamkY+iyC7L0IpXx0xk96f288g4qynpNug2Ie
wKDTy0lYQlSaceDXdKzQSJijNRuhWDJ4UhY3ryyjfl9aDnzl7orH+uFX+MF66NK41IaBIFir+Qso
rOMqutL7JuzrBV8MnfTwsb5HyN300XzYzXDwqFZDAtuEXDfqWI5PiYDOdiBa7fLJ/2NUIs57cOSC
iNrDF+BHmrlCZHLE/XwaKPkh8AABFfaI8n2lsoS9+uhWReAyvD2ilnHkOu4JSC6Z7mwt/VnkQziz
bITOXSXf3Al7QtaxfoK9zsSxNryPMx5e7SfVFhICvy7VzE8aofoBjw0l5ACxq5yx6nuOTZsUwJTj
xG5R9efQAWb2zJopboAJnmix5cxtylNuLkyCZ3PXAHslDdqotOXWnk7QfuhCfCC/f3L93/ItPSh9
BR6FETYN+M7G+yITBnJJUIOpf+o7hT5k9E4UGV45F2yAPF27sfy1wTpMZhtq5KLYptZjMNegbGsx
d/+kOtYBEbdK2niTYXVaCmIddMmWJ0IIMLlZa/OzP6ArwxhQ8JOzHON4rbMCKEhE1arhm4q1l1bb
T6jYM0dBeQaDQLrkfgU+Ffe2QIA0n2cEp2m+I/7puCI670XZZjNjU09KGLf5IFlFcwn/jtdfKj+A
YJum+uupgFwB2rmg2GF+7paIKEIgvv7R9OdaECTrO/gcDm+sXTgCgekPZQbUW5wF4xSwVQKh2G15
R1MivxCin7Jenv0neOgFdX0RVuFj9fbtTsu/OJu+rZfjo5dbHpJ3wBIuq0d8Shd2BZ/DTYYRVAe1
uJA7x/BXat1v8YgZQD7iWCyaHWfNNWw4+zMPraA0AZskV7I4yEPQeuAgq7nCZgYltTkTNI9kOVKk
j4weXR/hEF8YVnR97caZHEdikKf8Ml3efQ28I1sA3m8XF028WSOqw/7YtllVFSh/hci69V2Sry+s
EaPjXKgl/LaiWdE6hi9hdLB9eO0DO09FaPlfMjOWqWP6eCC0GEE5I0+S5tXO9wSJeM7GH7uVH2MQ
lmTiJnHywmuiIrIuXow7KOfsvo1E5jjmTJ9O9w5QqS/TsoY8RSR5AIhW5Lx22T5S0nN/JE7Z50m+
R0V2LSMBoXnRv284XlbKWFuxL4FK4WbTfR7oiRA7QBkzcVWh2tulmSQarSjL1mGWvHu8D2ANSdJ/
LI+QROBhomPBTeWXY+6Slzl07h/mQRvUI3e/oGiIdo0oBGlwLL+YTCmAZrTGYaLwn67qBWdq4l2x
D5DYEWWtaRCZW0JeXUE15xaGYPT+7OIqv7YWF3Oa5quimK5vgmx5sEOHPPuYcM7ajb7/N4NxbuKo
Q0JyohU7RUJsl7cCws4ybzMkhxlinkKX3Xq6RVXbLg4/OFu7kSIVECjU2fHsuU5rEw1eXW5hRCzM
ps3O50qCeiVUEQnPfGoP+qq4Y70MWfdi/EWeNG5pxsFp4nLSizGGJybXqmDVxbuT/CTfF2AtEVs0
po5MobKIyg6uR2NRBjAV0Jb28+jNKJ39/yhxxJ9ADnZYria8dteUfqSeit7z0QKl6KMg4FWE72mJ
furl0OLq5jUJlt2Etz32Padq70Sddw1lLWUZieGtQnxVfuBVtW6tcCOPsjpr52V2xAGPmsHgR9WR
N57EolpU88wpjp+we0Wk2fzCheL0cxF5lKio2g8o1yvkV/dWqt0+YQB7/O+DHuSTsNfOLfD+w1TR
p2209NDO/mg3CDlr7iu3g7OQUzFhxjRRcNjBOTQ3P8bu9qVmht1kqL8vKKZiz96tjNI/xdRduQO5
/bIve735z2FP1Waa0N1k1REwDR2zgcA189mduk2EgHV0BFz+7L/T/golJMcbnZ+toONSVtG+dsC2
zEcfjc4uRBUdxQe3Ch72UhAfTLYRHhdkE610XIpr03/HKp2Gn/gs6HKDU3tnfDV5kSYyRLAbClKP
OZrM9GSX0RGGoRO1enrtoQVLDoYYYJ6OD3xZgqzVP6A+v/P9BCAJC1wp7VLcxXb3cfYTtVV4FNgF
jUnjdGspUnjXm7kxqGwFkcaPXS8AGZT5F4Hyavli9ACtFklKCR9OjkWcZ+bkfypzNDtSC6pIno8d
n3bfIVGz1nTF8Icf9610HfTqAsRC2/ZNdm+8mqPuou/Cx9y+oSmgcbekaSQoRr12Lv7Yazu2CXgS
zaScy50uY5afLlF+7mPnsRmsGE+/JtzSctYoerCt6+TfaifLJdYKZFj/5XCF1fJ+c568Qs72zjUD
Z76W2c9JHwy7VJjIUsS9ABeGZNdeWIzrK/Bw95M8lx71pnUxlv1SBl5AAtsyPY5bbyVFeYWJnOU4
gTakBzjxi0BdIAa01Yz58S3xgkE+iquB69cNFf0c7ru6lnzlXKvF7QpkGWD8ZGON9BTc52sgGRfc
TdyKGxbBcJPUoYY7+YzW3AH8RTvEvNeLc7ZA70qzGjJLeP+0cSQ4ORmw6SP8RTjyXxFTkw0h3sn3
LqxivmpTfYYkekKcgAk6q9VIOl4lCTxyk/hmZf5s1AxHNE+Cov0uvw9/TThXyBk+MIouIMbx90r7
wpahgE+GJSkBRq7Pj9+mM/Q2MUOaC/k3mran79tkqZrzehXiQpuPVgiYQ2UA4FPjmvI94nkirjea
DPdxFjAaAV+SKKfXGYv+my/e2z6jXEYkxRcWpaKlTtpkWaPLhTbulJbihwBID+J8yJp+ru6/o0eH
bjS8r30VF+pTZPml4hyrujrRkOiRG6z3ZsgoYbDawHVa+EYnj4XmXrMOfui2jo+QozFqW++p1Zjn
rvzvAuii43JeI3ZW8o9k7iyftfprZC9+QAMZ2tMhGYyrdDO1YNoXNoBDxcxFrKU6W7tn7M0AonH+
YURAqvY8VQebbh6/fUEkhbimM1YvIldkQppPRTQHTRdkW7b8OVr8lHg7EEYPKcz6rCTdOJzIndtO
FGGrEhT+ND+WiCIMK2wGGEIm8ev0npR4WqrAimV1d0qv6NhsXDy9IfTISuXs6X1RBrPu6eq/fs2g
gByfxRo5M4p+YI8IsPgXipKEC1wly+Vb02vikSoiQwuO1lRJAr2R0Ny6rn2V2f6rBCUkWZxA9m2v
9DM2xVzOEgrThCG0He7HPj7GzkWGgPn5n8VfoFI3NvxKhzspqh23kprrK86Ca6J66rApg2Ri6+XK
NnzuZ2GkDYGbgavrQ1hYs3ZwXiuym7P3qIf2S60B70oF/p6alWrWZJNJxgTMMxiagNqtIZ0jijHr
wR1ldbn6f/R7Iq490Uitk98Ar95wMLe3U4yfGTZmejpgVLjgtMQkmQnbQVhTNtcP+jQ1YAN5+KxW
V0QHG0QrGFPhaGh3MvYB0oyg4wuZJw1XqL7A9LPklpDd6lFB9UdLyJnkMtNLKBZNFJhZeskDFr0z
Swiusr35Q2HBSsTiTHZa1KSGjP9dB0Sqs7TeG8EMa8egKCoD4jTNlyWfH3qheocEvYg40NmNyowf
CxyUUgQKs+mOJBpQ1k5qwP2nCf4DlBm9+sTF8k6/yddgosS6EkSHLeNt931SuQ3Za9xItNB81XSJ
pVuhf0/SlA34TdG+r97afQpQKpi3iFztJb9ZbaxGgJMP6fxCy10ow+Z69gWQspgv4LCosQcqWCEx
/iEeONf9pYIiDtJwXyaj98JGI5Ff4FsVsGHEeCYrdMob/w3g+OKChLABLRbIwML7zjqbnm5bP9UN
Gh11dt3q+gpSXGlnGDZ8e6XxxxxEvyOTx7eOx7OHUn3kqQOOTOKOtXkAQRc5iFJCoJZcD8Fl0/UC
FIG32YcH5LSM7al8Mg50lEZ5n2CV9eFI3bpJB8Bmjq2kcdrSEnPRr4wtBHjYBTX2zb1bNHpLmULb
kHV1GDs6igfZVs1kqOvuVWR7ZJl8t12/diOIuBANS8v9W3kYB0a5hNibWZhVwtQCeeEQSbktuiqU
poet2XDxmSsOT/W4xtBXdNxnwBaUYEmcQWa4AwcKwAV4tAH9BuCvTTCyseCZIZFlCZ6Pq84HjWSk
rmOlX4eQgEAEvD0Toz1w+xQLbqZABRhdst5x3caLhsMGhPD0x6b6zcrQTNmEsgi+lvrM6s9MnPnm
3bSsSarazI6BzVBxIDoKtOqqoPoU/9rdQ6mN6x40QF6C9lJS6meiEPN1L0T3EvZycirNDVViQP2F
dzyDhCmMcCXZZgIIW+xO7WdOIhrwaZr/9u9xlX5OrAjyW5MSW1MZIIXh5zuvt7kkiU42y8s97PDz
aGvRXHjSs+yra/WeX2iowwba1GQDR1tnefm90Zh5+5ndPIJTUjSCscPBStG0k9CtCQawIDcWK5C+
3QWdaWujbPDetloQH3dbIj+tDFRJqIWU4qNTA4037U+mJlzQ65jQ/j+OSKILHG0sieaJGgCYW+2u
wpt5y7Y0xDFlBwu44o+xIVIQrDGdllM0xb3Gsy9c/9snX5yi/VVjHpocs+MErK1Hpvl2+JYo9gye
XjCXnonI9ZaJeyIOBNIMzZpM/xUefqT2lWHAkSpbkwgriVC9xXx+Bnjao30/K+XmTF1B2ALB8P9M
qwRdhDjfm9QhwI9zOFSXe7yMnkmrmohAyU6imVkh7ANRB4V9zK2zvUqjE2Zzgq1TIo30y8CDw4On
owz+qEtovT95ULb2QfrFEgoIUbTsUziCXeEf+dyLqJ72Onhh2sVBHCw7c0Zr0ypiMf4KwsyuAoFV
B3Xi9YZraYc9heoOMPMfXenkF7ihiQuwzJsr+1gIiEqNzN4u3bGkxBwL3Nto9QA0yxJ9Mq94t+uZ
pJXE2ewuYYxtUbJ8CXHvCyT50ZI4p0JMh1E6xAp8I4mtbcJlZiN8j2nnKp4Y3cy5rUBZR8MtivY9
dtOsf1z6attJK2StJsJ2c783PI8xpIWtK1Lw2zSIG8/Tq5X38/wE4Eec64sEYLhL7IM5N+XEpbyW
y1Gazx0bGQOW6SM8SY2olvTPqHrAUx/nMiKuTVRzT3me9A2L4pWZB3S82Jb0cyctqF0iDwUJJ+rv
OOg42DK2+DZOWj8zjKkT/dDXaOtG2vKBz5hW1RQffkh4AkM5qgdTxPCfU/Bi/mpDKIew9H7LRVwJ
glFc8Sr6xikPvGfJrjWlKO0moX7bmF0dX2C5g905GX42GOnIEL2DErjxlQjwBIRD1+lBHoCM0n/P
Oze2dlIHysK1nHOKbxzRcuCoABa/XI320anBgBzoJq1S5rbv6SjepsBuxJe3ieSCg6Xi1YikHeo8
lFUCBId+tDUyqG/7j823t2pW+Rx0Jh557UjjSaPtq5g6Y68AEm5dY91O+3an7AuUrx2aXH3XVahA
R8htSHgRQPY8SuW0aopFY4xNSVyeROxUAzMMa8Fl/Mz86ZH/0WqKCu/ROZfIqlhU+rrJSWKIJnGY
RYsEdBjVK/0G7q7/vtRCiPVc/E/oZ0v2vqDAuE0ptDFDULA26tbgQY+knD0E1tifN+svRXDrp6d8
F2z0tHBCpDQTd4TS/Fev1/PSB+vvFtm/8olgJ4iWHxWR4jVFCqWk2xEikqRKFq+lOsA0Ez+uKaJk
N0IbTPKb8gZc4YAn9tsKHU3557nTUrkIGBXo8OE90mMb1MgpYEozrK7xr8Fywv7bF6YGxsQmCyDw
zrFL7H0evEpYHFJMckCUapH81s/oieFp9a9mAlK/H0fj27R6KLrgdUN7KaUax9Xs/ns4tFAF4NU6
eQDkIvRezgJmC5TzpG4RiRqblniNI2V9uY4MunOTWN3X43QUHQBKJquZWqJp4QJWMtYA3z2pfjea
Mx54n64fQtkOEq0qulCzdf0EQQXJQi8i5KVCRkLd19EinRUwcmoPB4xT2sq4su024uxfvdAcSuuf
/t2RQ3dPyCflXAjrZ3CTSSIodXwqwFazIFSWKuT9lsUlwkbbrMRMsh5waaIgwKsIwNRAmEGLlKCm
DI+L94WFOJCxRQ+/2xV7E4aJ+13m5lCrukBhesY2nVJTfPKCr8EpSnW59Oa+l38BGICHODuFvPb0
/IKKqH10Qt1YZqwMxAw8cPLQXjl/AxKRRavNkp0sW031eo84VLKhqujzNmo5cYPl8L1GwJPImFpG
vuQe1MZeyEbrxvNFaWe3GVV7yMj/eQ6HEomRpPlBfKAfiTKi8PQ4I1VgkmyJiCK/pblHP+32wMp9
zR4LOjk7yhktwhqK/DH7llpTG6Tc4Zp/6K/yPwKc6oHhSHnnVANxCAWGVKiA7TcycnQpDNY4qBNq
B3sF8xxpYEMZcWzIbYh19JDTS7z1Te+LrymMDbj2y7+mHkTZEwHHMRkr9lUxqZyZaXb9OZyL+0go
D1DErFVs1RLNXO0UiRv+ynMP5b4/Xi/r5NCx8qcaDqPH4xElh1du+gKwvpLrtD4gj6uA8U+BMdNy
XIOswnRqTHlPzd2jhXOMJwGAspZdaTGWK64PsMToFLQ0zgbtcqKv2cBJy8GvSHqBC3nD4KaSTCGS
aSC1fvhA97XGm36iMIRVRLvyJjCWdiOpiYfcDUe49qqtytau02iKSmeEMmjeFar2fbVEuGwWrhw7
PVjk6d/23O194QWuCcrQS6wdpXcd5PhkLgU0JRmRvN+9Kl7fHy7C35n51axEaQOixHywUQy3jIyO
8aoY0mja80uoBcmjIWKmFx3g1Rn0pmEJz+YUOb16TSvV1vWrFE5pk0nM2ZdoaZ5rzUCDYI4mhnhT
da4jumG+79MemoZsbPBiD51nfmSyn8m7kqZ3PDyonwsFdcWhef/4Py+vepOTfFk2t7aUGyf85J3G
nGSm6uqSp4ej/2ExgRELTByuh/Rf64B6T7Q+jkSW7YFZDZF1+jKDK3rtEl/zT/y1FvZy+Yj27KZH
U1WByV7TzrgRRdodmB6GAXIWbLhJlG8UnkrkYwmqY2Uz+l1ZjaV8P7jpnDI8tN0cWhxogunYzvL3
XxG+GZo/rY7YbA61NuA4IaM1Jj6AmfL0stoMf93/Sy+1+avsTi8LTR1zEdK18SrxGmK/p4nVO52M
q/S+qjHIN1gylXQrhX5o0fDDwSlIU7SB+bY+5UDuhDCb/CIEGrG6uwgf1j6V3x3F5Js7BnoGEt+x
Wan902KTBxlMeBBJmc9ikP65DEAQMLnGM9s2u0nC92scEhpY/FKB6zA445yMk0vcnxKw5qFt0KVp
WkFzOPQuGqyGssTu0zwtyRQPpLCoxKw7AbElKsjmB6K+4x6tCWNor2mLM+gQrPW3P+F9b8P+vRwl
Mi8dcFD3OwD2s4ruAymyVC5A2TuhKg/FYxpVhJv6uKN7Oxt/pux21w8g+ppX1ASUF2sd8D4FHUm+
opYVKkHNrvdCjCPE8S3qrFttFOg731g58VkKDT5SuaYPGLa/IuNPh6uU0ud6Fr3RqZ77cPAciUA1
FlHvcx3wEEGsR0i7gu30hMm7Ef7i15Kx3sbJo+H0SkRVrYwVv/TXXE2CfVsCNqEF5r2Vqqzbh2jh
SZM/410Vuj6iotxB7i/hGVW2FmycHfwKzpbjrptmUkQyTHCBTpiI7hD4ZMzlsdlGvmRx+m+qp+j4
Xd9Pd2sR2SdY2gGU7J+XyDYzRz15BdvqHE55f2rDTgA/35k4VjGIOnODpVfY543C5zTA2mSgBvBN
2Y+Mxq756OUnFPPc8fpNMAILYb3ar6ay2L5TjTsKBNpDAtQuO0HwkqWbCvmJkc8c4cJbGKqI6X9o
U5mCfvQn8pSfZi0IK9mEmJ47K36vSv1pJAStwwUgw1B5OkhLpAEQ8qEUwr6a1MUMej+qhIbuAQMn
ia/ytyv1SBtSzA1mqIomLfBh+ejFg7hCn2x7db/8JtQQAX8sKRNNGL+4jM0ERwxJJMYZMmKrHDZm
hR9T700cL7MqS4FqZzvR6ZbDfgqmwvNSpv4umfm/ENQxUDKE6bs75uUXSE+9E/+cLMq0eeF0mxl9
WtD9mmH/cC2rbMvFuYy4wRRPhqNrJ/sNKTd03ytc0PQzDSo7QyhlCZC0K9M6OzPc6NNXybJsrBWO
bBkU+TOB2a9voxL1BHx2p7N2hR9e0EGQiD2hjDmKH0YXSLMfo3DtM0xjcc2C1cYRK2q3ORC+4PjX
TpCnqnp/wXs4+M8e8I6PyU+VFSzNF5xI4ASt5Bz3vQi0cPzRJqWuFT7s1cKDvcAFnh0A1F67wnrv
IBiu6ZT6pkwsorwXEiT5GWGSFFgoAfl5yVYwRvqFEdTMziyJAzjLXHSb7dASz2bgcLLyqs7ONfqB
xvFZd0hwH4NksJctj6dmfCP3k9vkVojVPsOQT0AhS/I4FtcJLCteIdo+NuFMFlsfw+GTj5E+fOLA
er4RiUTBoPk9xSO8zzfP8RpOq9zFOJunuEjRb2KGMau9gDk85jxn0tCVl/F64XC6f+MgjU3sKmFo
pkVIVrhkSKYLEWTjdLqt6wZ+zKi/mVIeP6yy1Ywc711RZBOVljx0FeCNL3L1SCrVmXuuhsZy9vvf
0iSjMR7LTdmID78/XnZFGk1N+qaKTyrgWZ3aK7VlhrXQyGKaXUdq4Ox+POOCt0CNzbnArYqV4lKS
nT/CRi2F++gAyVFBjv+oJXw0QFWuHxkPD3tnuD8r5ncIACS1yRoIAbCuz3L6Q+S1claVrluKGXzK
XftnY/UCWiqaWyzlQvJz4c3W+GpFApNX2J+QwCg4Ef9PeC/z5Ya/LK1SiWqFN289i9SJ4H7dgpaU
dALHXMOxAvzozoaBTvmuL9sINioGZ5+hIE4I2w6+wGG7E2jfTVTqbTbtJk64aozU+3MeL0+gXjad
FGVLCYPNF7nX9bc5Jfq6fPaSPC8kl6E93650WWpfPLV463F85KO/UlK0iJKDl3AtDxgtR2Yy3JqB
qxyU19nXAHP2xrTK+hwuX5zywuwZrObQelIYIuF46sG7PEHx1Cct14MrltyWtwhtrIXS7PQmIOuY
9xg0d2mR5fT8BW0LihUkBp6eY1JVu3OvKsOduCbk+NQvPZdo4Jbp6MIElyPIUvCCelUNBBxDTGbk
SZD/VTeLSKqApcAO1VnFXbxaRE5SHNA7HZOPIOnYYxbdKBnVIOyd4B1ZFTo5oaDbvBNFSv7zZHqV
238bwbnuQlh6ns9V2zUvIndTiqSdyjomYMfFKZ3nbNUbA5sHXhdK4Ucr/kFss+flNBAeNELRdyKg
lvJ0HCksTcXR8VadKUPGcmmd5Ge9V0PegyyrR/vEiW3+5csjl5vW3uZ6oqqtTn/auhTje9QqTZOi
RUjQo4YtllEG+dqzr84+ML+jmZc2PK6tzY6Ta+Uu8HUz1df5pUULOUehVPNZlJdaH1ZqqYaRNLRt
XeY+1ST6FuKqONYGqOU4qJP+P6TCJY70aVRFozRX7WObJplC98qWIMoAe10R2LZ+c3C6ZiAhpcWA
S+l6J+R4nEdk7u65VKfVcbWJpII0RifwPzxxSp3UUw2I/Y6u7xf+78g8IXnwR/UIEXJBN4TtCmrc
beJqxsHjIa0OERfz+HCMXFiV1ivJx9T8dzRxkLwlclapsn89ORq6xhlxCW8r29z/cFji2u0RohDX
iYyOgSZTO+Eun6Ux3LZXiErgQ3w+ijW1B45Vu1Nz1b8uZBQAvGTZEYQmTTZMCvVB0R6tbFNrfxOL
xBf1Se8jAVfQOMn+GS48KC0VSHWMqlgRJWB8GTA0TV6kVHMCWcDDjgh3qxb4LZMmkUs2oKqvkNxd
i12kNqoJFuk+tXHFK5OH6HG+YomQ+QQUZz53Fs6vHAdEb3JAS3IohM/xOfUgO4WDIsf6nAvKGPWo
9sevC8wNWE6HDezKFtjJfIMe3BFO6mxhcwz9+B+vOMQD/K9MJ2/8oNay7nAqDFC2JL1hKFVaMeYx
vel9sSb/S6cZCkW+zRl4k9CNbG9q419lCzU074QKRExt0/VdRulG92SH4T/1Gs9Ob1koEqpRB6Ft
xnNu7J6vqRof7jlrtvIEN53Z66mtTvm0csD0pfiUTQkQ5dPzvi6zq9L3Cf3NzIzU56NWR1SIw853
BLHbJsLIU4zIpcqtTXkawCdxl1Y/iNIFBef4WOQTFjHlboRqU4bde4DXwc9puzI/TilWw5Y0I718
H47aAgn/XgQ7q0OW3Ei5I0lkqS6QLhweevXNgPyaZvtYdEKW1gPiTxdgO7Mgsse1XSzTDtVpIKsx
Hma63QKdWpTr+fS8pmd0KwpcCw22Jg3JHZKfw5eYMziMMO2iYo5gIetYDv/7zlrDysqhIRVM5dbB
IfFL1F27XibCR7a9qD2F1SOD9eHQfIvEdip/Ps6OmrY1OAe1ZJLZz5ROzE4rJCfAotNhbLsM7q15
FjbEyC+VvE4IyZqOJPi7hkU0vQOCaMDVnNEbeSjCFDTUCkx+AUbp1Di0yh7hMdRoUSomYqqgh3YZ
16hHpHmlomiQGtyHe0Lqc7suwkxJqIMSQY72xGRi4TUwUgkykwWdSmms8NECf2QLm+TIlQSSMwKV
ePHFpkVKoaypz/aHv+qahOpXrtxvEU3roYRTaDky7IM/ThqWhqnBjdH4BSCAVO+ElZ4np65EUMbn
XJydMHVsfqOQzMDrL6pT1uGqowjDU1UPto7/jWV5DFuH3j1gHz8FuW5XT23y6O7K8q/gbN7xCMOM
atWFBElcRgyd+Fdt0gLvwgK/RUngWYneRV6Vh4OsrjRfftwGFrmeqhxOv2OjWamzc0aKWmAZ8HOB
d4sh+5wg6DGhy7RTPq4yw1uVEIwkSlKRoFukjDYXgutt2YYTlml4AqEArRQrVLWwusiUCX0lHv9R
GyC2B+O9l8PurW/gsi0gO5CKDZmTh47HLIHi6qD9yE/zN/xjhSS4EUjCmZO7laFYqajdpVitxd1+
1Cne/4kAcrTTK0Wad98cf9i/ynjIVc5NzTYS+MjSXFBTVBdhxaLXH0CI+juxbjwtwmjT5FSrsbc2
ki+8iesmzDXvTRm2Km+PZS8HYBX7ZdZzhm2UTJg3POMsqQhKi9SmLnePRZFnx3znyY10M7e+gKim
WJVmq0+KGua5X1iUjx8EtpC8gyRFzFEfufLQDipcSiSMBndmK6lxbvpRWJxvGzJc2Jqe+MVwvyuz
Kfk50vqNWno8gm85/kyuVy/f1VMl333aQKVlGCJIfL5Cdkr77zDgWVolZNXM+hbdySyqqD1UWGZv
rTJYcQCPaCPl532X0SSOIFIkvb2iSQw9BloVUGPgHAoaL55/QUTHvI23LtOTsxRg9qbD6fk2IiDz
yH/1aYMMAyWybtUJO6lowUz9+7K8DkCCpZPYD+JJTI7LOV4VDkZkoJtp2uy/wmEDkU6HlNFotkJA
ZnNtRA4Zj0RQdNGPB2QB64aPZWyqD84+DJNbLHxaA1/M2lV9YmwgYIclPASIC5uefj+F4mDeI334
rbznRr4L/o4WzTRUZ6PPKmOYTKKyM/DXZLMwmLItuKYOm7ElHRaJtnJOMSWCSpF9rJdNjJIEemlb
H6u3nYfwcumgzPasLGUKfbyi6NWR9vfyDhSzkUlL0Gkw1DVgdbUVWbyEsryM2zaLQKpQi/0gSfbW
U7HJKE/pCIR9/zwQlxZE16iARLsETfhsuvvKkRz0fo0UMX8aakT4pOJob4ZNLJptP9XpwXdcVvjd
lM8M+CSlhUMwWtYFYq9VHJBYeg5YMP/lpjMZ9sgUZZUjTOrLDDmBiVVQU9w9m9fcsKB0ymE2iFvn
vDkl3PzaZprSXgIyfl4f2mmQ5kc6SJZDu32USRpOhOavuegBB7eyMWqCqqVtJa31axaLCniRTpaq
89w65rIvayjr9QMcipNizqEOwDT/4KduwxgwwF6kmzF7Te1cQUvPQ1Kf5G20foP0E8KhX5K8OaU9
a2LaHCTca5xhHXBwS/6okoWYU38vrtJ4UnSfLn3a5tBbFFCMOEIqSobkF5O3xnuMx+S/nIyWaZCZ
V71YMoQhKDzL7spUAG3MZzDAiv7VStFPrlORuCTQrcjQ9UBc44gSGbpA6L9r3AYbZn3EN/MDyj1p
ioSjjckezvuJB31T5QLyqlQDXKSbgM7DcrYzTpViStPCMmCuWl0Tk2iay+k7BKCzTpszJ5sD7c/M
IU4Ccw/7Zbg7cbu4paWcfoamZ1whUQybpnma6fpcIr0Io9gJVYstIRZ4meUdUXReMz5otYCb7oyt
i1fQ+4BtDj5zMIvaEaaJSnBJBVRrKyJtXJ1Id7kr9AT/c3DBh95OQhyXQbr8QDjfO/IPKxwXF6wp
/lBWuaprsumMHS8uxnwsfrQZ5F0O3O8aJ/ARbHn3Ft6eI3n6f0FgMRgbCTMapI6pB/LwylASK2Xb
3+IcCmc1WML9ML0RZGozZClckGiSwwpEJz3CLz1Qfj3VEv/UAr9LLgjl/cBM8Uuela0lxlr0l+hJ
W8n/BiZZhAD8rGU+wWC1gyAE9b4CrMrtRIirCkAlIOHcW8EIpmyQFNrC9tUHPpBihPJ1wAjwNhrm
J8cxDc1pWBxQDZsYqcQgX82dDZGy0j3zKvxNJLieK3x22GCMApdYcmkwCAOQNwR/ORtrBf8zTaET
HrYoNs1by9xqqDnNvp4vd964hIlLfNhk3/0OjkWOp3pad9NBlH68kORqSz4DpaLynnmsElF6TQ76
ZU0YM1eQgGtqWR0+cppcbg0iQGGNMbQHRRmamUe3K8X97vhHAouGSlhK4Q1TRIOaFbmMdm67jBOT
0xqsImybN8oLZT6+ZXimbaUYKlIWLPWGuY+2cukm8zoTka8E/PgDHKB+pBP/FNLtsjbI/cu8jGEA
Q8UO5VL7us23ilhEA6fdSIL+9Z0YPtyPzv0H5U2+0tI3+uMuPlhfe5nWqXnqlVNj5X9bdaIV3hrJ
nBeMaw3s8AtlY44SkHSjrsZbe5YozCm5f84oahlaO7Owjr0d0Ec1D8yLhT7tfBbk6YiTaokNv5ve
gadRTEfPgQoz2k99iNYk30eG30e7f0E9ezYgbe4dFfBJ3LLcxOA2lOdeH+NcXDeywLuJI9U8MqJH
6BYOuJ0d4l1vNLhlUcKTRvMFlyIj3hbxLf2WiwAfkVUbQPERzSk9ncD1EQsHm0P58RCWpPX+9bkE
MibW8HAFNTZsvRVifSOMp2fcTAPgUoETwvFU+FTORdamLscOKDFPiZhxO0RdbO6mlDv9VzYrGxUL
0d7h0/zWTp4Y+iMakoPvN/T1EkQwAzFfd6po+kEvprvnmd4IgdqSCywJIJUamI+UZ9RAikxz5NCa
ktBYWOCKhilaLWuxhJM7xGpElM2aH9mV3jFYK40vt3xl/q1JIu59fxNG1x7nOOhzV4F8wCZ/mYel
VQ2FpKtQfKR9kVaxfWlHClW3GoUKCRavfLLYmTZX7idtcYsUQGnecZ6TTlf/IZoBoys9r/Zsuwk3
gxKtFwzV3XKuE/BqCu/TdzATUhgyTlq3TebOeqteGJca0qIRVxk5M5ZhvYXMuSIvAFAsgKHJGCJC
Wdxt9vWbPTp76yIOZuH6AV5ca6oRA7TW0JxO9GQ9Sya07Cy2YWphiySUIcUUMeIOzYQQfSvNbV9C
7itRxC6vD5BoGxtnRtIl3taq9PrYH38knlU7zgNxhyj6gjDRSwU4B6yAm/DrzrZpiMkic6yGb78w
QadsjUAjtW9Gf0qU17NAJsI3pWGn8wh/e0/dMxmyqSu4Peh2BYAY5oTMyRfXFX2JcaVQw4nuL/63
LBoNNirgJ/yvOXBcKTtCXtJDOZeGshGZO5qmPphG3Tz8OQeGv1ELDPi6KEIfLD/Z7wdpCy/vosEs
UNc/awj7Pwy3eXnsN9n+Iqt0E/FhsceidkA99e7tFgY4WwUXvd3ovdyTk/o8W7OINLqO/8G26a2b
7AUtoSH38GBN95AAnPxzWYAC8K1DtL8VWRxp+ESs9zng4D6uJcMl7PGv3BbcGJmSFsdKwkKgbxsj
hd7QjZq6pD9JTe2urkOEG7/oUI3fCxkyrtGYBil2ggPsJfRq3fpAkLuBbQHIF1IsM5dxhU7rvVO6
5ZSr1GpbOpUpcwpGwCLxLRyFgcZK5siARxMKuPv0eMrtXmoHMtAOZSQSerRmj5Wakbs9evtHCpL3
miMj6u0dI75Kv+1txdniWtmB0V5egkdop4SVok0lZOz/IyDFq3Q6zZNd+45Ls9vmwSlwM/r4avgy
0cbq43wOTyfP1eLy58IowqpkDyNcJUw2gcNRACukr/bfSWefrZFNf4BfSLOBBIY1u1m3OkwGrk/T
VviKYJI5vzuhOTsqbTAnU7KKY2ODcTLyoSRnOOP9hKsXRI6P+vvztMHimpPszPJ7v3z8tN4+sOQt
3Ui1nBqlG+KguIPkD6KelVlmzc2lZO7Zt0FPYTBs1YLiiVyWkEXzY0McjGY6zn7ECXyidgLtcPSJ
OeQNrBuF9g+5QFsLF8OBtfT9UwAR1ryUXnHEDCdDtjdYDg2cN3/YO/op00mYBVTlWfDmgvWcHx3O
BlvuOUP/4GcwqzbqLOJ5SbvG1qxBtWNrJ9wO3VCZWis5MyhodNwLJlXdu5Smyp35trGU36qwar2D
zQMfmqEueexWcWLgMz5sDVn4FewVcowU0hnaQE5gygl37Zmtg+wf1rfeMro4/0TMG2oP5fPzpmtH
jDempLAH5L6FCw2gVR9WrbMlDkEbktHLHX4lSAUQoys6NQij/uE1g579nziaXGfsLkkRbsjITpHd
NgJOKpw44ASh3x4vblnf+J5P+pqu6m4SzGERDpfbjfAeGzfWET99At9qXPxxXxIFKSwsoFCv/28J
MAqJBCTdbZ5yVFPH44JyXtvjA5tpV9QT8iEqb/Nu4yDc6fxKkLIfXyi7fzxyZ/D3ZdGEgBpCJ4mp
kStXXPNr/oKhNR3x//1APULBs2526t8La1V71zmyXMNGpRyoFr6dWTJRl5kEg0W2UfdvfBlj4qXc
Pth39t6eVOmp23fHIK8E9qW6vOkDNyN1EybK0JzKm5IydhUkrmgOnFDOWKmaRQfiDn9iLkOGcDmQ
6JfxpsogmxNw0g0xtmwedWlDi4BI229tC5osRDReKyCRGE4jr6HprPvms+nihFV4vPs+41Dmeb/g
cFGTTNbzt9tGDo2yQSUNkx87UCaMzyFt//HxbiD3XIisdULLcOJbOu2iJRniUG36EG+1Q0uEz4b9
iWDYYb5wOJeFBQPdIKpxTEUYM2Y2x4nF8lpP+E37FPE5Xl7IwP2AkDEYNROzhABEV0sw+Sji9gS3
3a8dPvn/tJVHS15Sb3xTytBkYKqR2CSPRW/jckZ3MbdKSavh7nUBZ8ZwZXjSRYvNEYqgvNdoUWt2
ihXjbaeuSbEzgXR00e80w0Do92ddaNeUU1UdIA4D9Zi+QbKfCNvnUINGx/XugWMiKKVz2Q8SI7+C
PaZPv4BOVzTJYUFpE03TiUkLAoUW8Gvy8sRWzns4vts48tPBffVqpMXyiMfIJxlE49+f8hy6WpmM
Z7sLQf8WDQe3d8B0jnfwYe4gT94Hr5lLmlH2BJjWSre/gULk/a8fpfOYS204PbN9mRbbgUoRnM0g
/Qn+UhPk6j7QJ9qEE+VSYFK8dkxyVVaAxdcfdTqmtioX6qgao5KKHLSGwVHgHF6r++BKbkYnaZaG
ZTQ2iR5m5NrQTh8KJfMZCbtuiNusUlIyQ4c5UxEmiByARKbFnuJfmrunGu8orxrTUZ66Qat35nVo
HQawzi7TW0RkzE3iQfsbxLDDbbCJokYMiBq2YOV/OeT+tvNhdfBeuCFN3jS0lJmrye/lp2D2/JOW
+rOg9whQdlCronkIkW2Ups/gokqY/1WVcINSM1gsvQIKvEUJySzm/rIFQ6RvdVcmm2vpHBB2Cyb0
ApHJuqSFe2XSzmjBA14r19VWSZKnSNjAnm/uQ/cpyQ61UmnCjHue6Hs3AkYMrPCf5ERmXbpnuJ45
0t6skFPnAMxD80+Kfp6PzsHeB18wiP2+Icv8xlOqSg0r/asT3RmH+QMXy8XxC1rFEzDKpRsb6gsn
Os+jnqjKEp0493nXI4q03uRBOlEhTsdpER3AUpCjNKaMcSX0X3ACwydAvQNFhcfl6T4eXNAX3Yv0
aPBfH8TAQggNByiqYfIA7M9xNvXSEXjkdczEZutxufRCzbLIfR2kPwCg1Tezd1SG1rs6ggYYGC9S
KUnjFaUYjdmI+nT9Yf7GPEgT4dF2khGYfCUcUMgq3JA3oiPBfIl8HfZliU9JUXPoB00Uk1LhysxI
r+6bzY28rjXwlz7Kxz3njI88EA0lSo1Fox4ZGG/KVheDrxZV9SxBm2eEHiOWrmuz5LTH5LBnncB3
gsVEL6MWsfM5tnwiBmRifFeHp22OA4ep2PiGDiREdYQlm6n5UCmHFchTGMcC2s9M2NXw5dSnsPx3
7oxja5wUj6QwlsVlQRjIBAA2NYhfgvRX5xB4XXy+qVerMkwg/iS9qNHmoID7//XQFI+d9Vb1xC4c
+hqG2MwG+sDrmxTzu1gjMIUCdAhTWnYww53+sJzoHb96uqdGsP1YuRSyhURedtBU4lexxOScHli4
XaKfuyjI094FGP6sJlcWonkei4vSE7ZdHOvpvnCVj1DSQhxBlVzsUaukYD2dy242Hu3N4JpNCCYm
V119Am6h/0X2DUZ0Y2exgUTeCjR3t0TEsRfYB2qV6Ftqg/h/l4pxMnx/dn6QTh/TiNCSZXme3BlH
/KXaTewYqk3Fdf7BTzPUDCW2w/E7KcN1/tOYbY52PTJU6H+q3ro985Nxin+SsKEmxKRdOnE6QAbL
Mj9bOlcmZ0KWiVGCI/iMxxndpgGcYat7fYVMGtwHetqepARndBmWqQRPN0l8XTTkV5ScRQMlW8c/
6kID4Q5cfcL5+CeUrbrtbWypQrAsPpHJGAJXCwXMhWKSublgHokP9jO7ghXK4P2bLa6YR8JofzzA
za+KSZEcL2NFIpq43fudcGYBhLs5QrkuEOrUpfEQTfQBsAAnVLSWqNdL77Rkm27L4+adsSqOqa5K
IDWcogr6o5JBk8t6ZKP5GWwViWu+QLUeP8xX2e6QIxsp89nx7UdjXSPXs2pkhQnCY49C6j9wN8YU
peFI8SQLYHEgLew8LPosWIRkjQE0zjt085/1WYXoAsIyiSstTQznfSnrsi1aWd71nnStExYEYZEN
NpkM3hcHtFMl4zqYB1NN5MAd0sI9hG9D+yi/BpPAz+XTZpuc8jkxjnUOWG9wDt/G00NzUYYclBsR
pQ5FUuYZxhxHb1Dk8kOiqb35OwQicL5RW69c0Ta6UTLbN27jctfxHPnOuzG9apiA3m0YVmNN/EU9
Jk4YdgXsbc7PpJFoPMw3uFrqdjhc4DyQZHLTsPPQdNrtaRrxTw6pmPiU6IJhLztj1ThnZwyD84RU
hbXQv/Ce1sWBev1ooutCPckeTCdetxyKlruXRHjN5I2cxJKS0I285WNrxYUXljjuCP/T9JfcK8qC
ykXjpDjqsINxnXCHSnBxZV0OLjvsQb4yJecV3ixRNvn+2R27sAcDk3U83hOqeiZQZuUIaUwjQBOQ
z8LOqfsxU93cVT19YK66blI/xyok5NyTfCMUlGOpHWzZEB/X7fLA7t69kjpOO6mknCjyF3i5YHes
jEdmQZQJ6G/RHWbrJ4pBb5sqJoezfUB8YkyNOmNBg4z9lfWZoQhbIRzATv5/teGQMC5kixo4RqPG
Dnbg+lusVui4fsDCVUIbFuhE77c6V3hWYPabyMKjovZm5HbG3EvHyaXD5ZBYeFKRnkCcEb+oH14m
dl2OqYS70UixycUlRsENo13Cybl9xpvjPUGx5PQmM7A5qLdiheLw7evbJl+eDZE/SQFIYqP5NatD
QyGLF0yQhrnpBMfoQ/aXodbpHeCAu3rUM7p4wS8eDsGhN0Nxwz+cr8HKrifc2Bg48WmTHF6+thFV
nAAa0ZzL+hdnjAgO4rfbez9HAIW/seGvYrLbjTQ2bGnIV+iZXHucd9c+GEBrPnYssDAIjlG8c/Yw
dHPnkm2zlOsMCCHUfpHS+JpPf/kX3KiHqm4fid7nvvqoPOajb2Zuw1XKgDIJnyrVyfbvB1b1aqNq
YsQPsacDtCLDmKrMmdtQVjdM0V2mvOpaxNlBthL/WDTjedwCi6kqSN7b9tHmpz9MaDGuComUuXkD
rcZE8zsWQwJCcZhiTEsPoc69YU2N1NnnveIV7FkzBqlXaaGjq59vPojpUp/lPeQ9jQfWZ7NXOclV
1h4I7akXIlG+s2pMRdERJ8ieMrshSoFLbx324YyxA3H/c5yPZ8g7H0a4UPCBzXaLdlxZt91VC3rm
ty9EIO/EnwAk4/G01dFwVKKDZ3K41ifcNbPyYDWL6XKe3hG6fA4tvqZZEW5J7aniFsoVF3owZXlx
cBLdnRehNP7r0r70/s7b4KKRXBbFy9GcqLVF0YBe6ABp5FpskNl5i0REP6ES12kRhuuJ3mwu+40e
Nnt7yzDjhgb86cUU6OafPw5Zi0ki4XiYiD/EbsW4yIwRUoeB8XV3v9GjMhEGcI+BsImTXfYri82M
pwOdRFpCR/4JoH605GNcdUwy2bswbTUSug1rhjReKsxS9Siac3kGw6rpvCSk5buCRQrJKgpGDc39
D1c9EQbOlj7ypj2WPmBhiNh15J9xQygJJPz72JnstsVqbKASQNha23wQErCz1NJYhuxG9MoAz9x0
fu3hHPEnEtbGQab62LGRvG8SNpCpPg8R/B3anlyQnf+VJXOFu00IUxqf+GMUE4zC9gwwTu6ncI0A
LHgyyBLE82FBztuC95u/v4sXWVkkC/coD4VqUF3pT9iHGPeYPTAl0af2E4LkFEqr8ElsvetY7Yn/
8e7L8/FoMsmGq9mJxPwrrhX8uWPy0swicjvWsz1I2EydM9Jm3XERoeL+8XNKO8C5hmXtg8rzawhR
jrIkU3ZaLY97LgBO9GUQ/oTO1MDBTMeqmX0OfoIgJUqeUzdxgfrzL9GHVV3ITdV4kcRmNVwSYCVr
xh1Ei0vNNab81oOspJtzWwoB1SqVj6q/Sjt/etOzqfZedfmM6rmHOYQJpyBah4x07Oteprx79+lz
qcsts8l4UTgggMohxM8gW/pmGZ3zSsBaylBm8a6i9IEwx/Dnr7bQ67NHbdz1RGpw9cdvdKXnqilT
k3+xhST45wvmwY8VqfJZ8smMhISn1mz22I0XyFkCXb/q4Y1j2P7ER0pCQT4rqN4WEtow1w2ovVVY
Sr7FjNQRgkDVg100EXti2yXd2U5dUzaf0oj2ZjmPapOZhd99uoZWPJmK2NWSYbnSS722Kb9eYTxd
P1Ef6GFPT3UjZiN0uo6ZZ2KHUGT+rX75y7VP/PPYiXGdHV+ECvanPrkZo08xthc4e6nEC+HJ5P6U
rk5nByw7Hra71VX3M4NWK4eE7He9ICM+bZ09JYpzTvMeV4x3XW9mqpgTjLTBXFpykMKPpuR9QXj4
XcxfiPP9BpInXm7e86dfmNL8BVmHQBEWKWC/zuCfxM3aZ2rlm8ZOEz9Sd9/5EookhykNcfppSRrW
w/lv0h10k3hwkcri9W2gNgZTyUTY6pb5be8rRjc7mELLnednwjQjOrmQ6yKMJvnpaitIXJiHZH9J
oPpFI7Kr3yVXkgGDgCfDvdykyyaCR/wXA4bSPP/Lz8Y+xfmzjTSEysCVjcPfOaWiDmG6JgZVQN5I
linnPCpCmSAUj+JfI6kyRZzFSz0WCWShPR248OTwwPmG4LbMc+EPo4azqQmZ1/hjEpbPQkv+BWGT
VWvUt2LSG3WS9ztiAh+8aydgy+RZbuc2vUFuihvQk+JCUorOitxNkHkvnHE2VvfMeLlXUwr7Z499
0KoPNNIwWiVUmQgtIk5Za0TIS1jFkhSbi2lhl99949WfAXgZzpgLFeaS7tqHAOa5b+uRG4v8GOaG
SOMN2zOwLwh8CbxcKLwSVI3lNyJVN7oy7hTFxmh9JRGUADenbyPCNi7Q7HH52f79jMY7PIZe27z8
ayKeHfGhxQriUF5bJf2641RxLlIe11CaGBEp3DHo+rNTn4dRLO6E4BnELkJ9P/DAgb8aQ0vfDBUd
zO9V33bRdVDGi54K+mRcHex1tgAS5XoPaYqphzG4blB9XCrf4Zi9zdoSCtc1hqz4MfFlfxvk2yJQ
725DfbsyJPLhYutQdbRuABuoUXAUrQfrn4EGy/NJz0xzTWB+qnEe8Zx7JvKDx1j9dVVLm42kndXJ
/cXr6q91VVp4lRRDUXXpu60bzrR16koWVba+YFYXRjPSalE49CYdc9YiO5zIb3CVbK4+VR1BpjS4
EUivxLt20s7qQfTWzrrOdGpzzfgjgrJabpdk1Yn/xHiMmR0WVTDVNe3XxFNpsV0jMWi4DzTDUcDr
6vwG5IDQIkB3UEjU37kp4jP5J7KqgAI4KGE42WHp84JUOhz6oownkge2t0K5O9e2xPSdxfS8brae
OAQfUbduVCqukD0buv/VMzSTizCLvRqIj9u2773JWm5UXogHkKcHvvLvsV4rB0eXwQyZKZKGcPFB
3E1hcpvVtyYnFqlFIuOssfPnCu8HvFrUmu9N57dnqq6Sxjofwmxi5QYalFqsa4F7I1JL8UP/NUi+
/Tdtti6ADq3BgNI9aRDZGvYmesGTpZCk3u6587P1ruM+vZp/LTBGxmGOtjZBX0PTxjqnaSM9Z32F
v59eQJ/AWx+S9NFaaSWI1E/EOGnhYfpoW6BDlxuoGrIbGSFQrhVfZSzqU8xXr/9F+6qGr8sVWD+S
rmT7xFv00Sr72KMf3DiEwE77aa9DXZ8uS8xf663+k21k4N5hrHxl4l624c/79RhM5eDFAFoB0OJ+
Y7jQQDJFzjrOIRRqi7jV96J/UO2S3gdTzaCy/svdbM2VJUBdcqWzd24c2B8bevYVMYILALYnISxo
LiyIkyzZ2Ym64INE9So9VHKgAckWkNxc/xgH37BzkgQYl2/kMo42XL/i+fvzp/R6yX+FlycaAZau
2EBrtfW0cZJmKFj1uELMJryszquxLFOj2/ITI79ITzg6ETM4/uWiot+7FpBGXj5UDsk+ZrR17IsQ
t29pm05Rwqk73Wbw1a7/kTq5w6cw/q7OD12foy4WvSaKU4MV50D9YGb4b/febewxZ5FTmAGhHPxH
6gtLG0roADaG78zsAFFs4RrwKeSzmFeyAzQrVBVMK2XgELLZWJwEiid3GQ3BwvP9uZuVY2ZGlTDS
LIVKu0L+W/8Hlfh+edKsoeq2hPDG/hhgo244ouADRQcgnBAurRgB1xYVkE/C2UHlh9LDpJz69x2k
KqYF5qioNYMjLRDrozg4W0l5Ea4FVIi17MFeTt5eW1Pkj4DAqc6n0mRq0jisW7tOjhLQa2z9QYq5
EvsDCffi/3ylqRlWKo4lwtyRjI7xA0qJpbZOlyYMyfr1DPNLsaaLXJ9rPg/QDtuoYC78ZLDNrDHi
GBf0zQGhSGidpYiXrftu11ata7atlwJoXPj6UdHyuV1Y+7nmckd+ex6/N3XdZsLBXWb4lp8EDy7z
IYg9reK20gvegs1ZxoPbAJUe64S8Bse4CrlAI5DzQv/RonFAb3r9sD5BvKHNIJxkQNDREtwr0shZ
CjCnyAz8d7rx1B7B4OS3/IQfhoqIWAZaKvp2iDXvASwrm5NUvcRsVlzd9nzVlmV8mQ2VtWVogJml
MitebRHihmdN6gUNcWbjUgDRN4rkqrqoPGBcD7zRqqjYHKlUn5cEijIZDevjEJovYljceY8QSoK/
T6GQ1YYm8/iazIwYhV7N7wjUtkhVnI+trQl1EY+ge4EqRQRXg4OEN9yxJE7foVl8IYekMDw3+sKO
lkUwPRXkszQsQEHhwGAnojpfbqYU1ZyNRYAowf2Kn9/N9wAh0tGzTc9YwA3BqJ3Z52v7okVXcObC
JW2NxfnalT6JXZGaqCupHN+xvGSNTbb0WrViwD6JDtifiv/yRWwtPEJsyADV0Hh0m6XgtREHnDLx
Dl58mFYITSziz/V52HkNcyAb81tqhwGcLYDecOPYR1c8uJ6IiBKxN0hyIFbel1pnyZKE5VbKo+A6
PgMx8R76YOq8SlbwKrVvhjHoOUBhbV5As3xc+REWo0o7BQeDSa9RQjpPi1Ead9vcI2sdK9nmGEmo
O+atdZvR5Ne+ICFYC9yDVjPB6GgUKi9F6tsc1Kpy34yQ4WtPtZwh7dKRtEo+s3+63CBYFZnRB1dQ
F7U53k5mDQINs+5bLFguqxM7/autCRUoKzk43foAy8Gl40vnubFhjTAnE49tZQNhpJk7D21Z3Ybo
bDov3ToVfYK5lNU69TVjAQt5JTkNJqrqXb3Hi52nMqAi/0dE/Sw7tU2FR/n6c2VLkLWpOVJ4C5jB
6Ag1Lk16z1JvFOPgXYjyICDpERuYkrvxptnSk3ypo7wXFDy3WoKDyaa86RFzqBLddJEt+/FsRri0
h8H3T58ft12uuvePOL23zlLOzK3T6lkAPsPlREIJJMgE/YPKb4BoeCvZirDZTtiK6+jvT/TOWNld
C6SaxlOuW0hLyVzmD/06l9RXN2B0GkEVbr14C0UOG/RO0yTUTmKEOIFhgr4ozdp1Tdtq/gDJ6JOv
rxnSqfWeep8YjiNpDxv5986JIJvqrpHNIfLQYHjWmapRTwrW7pBtfq2zUVhSGOjIuj2shwxcj0n7
fUnPoipVHfcAszW32O65V5KA+9YVg0gJdR49FvmqMGKFQkj8jsVJS5wYaiU30csGNn4VRAM2Y9g8
z1IN8/jeks6vnsnoya89GQaqvTsXQ5ZJEvCw6LjxBMSJa1SeViAUUIC6L0eHDOnJ0t0wYRdm4/Yd
fRBQyiHhbf5HwX0HuKUz2GsB3yeXNk/K6QebeqkdiEtZ+nh9gPBWp//XkJXUhvFeumMXQafJEAW/
/h4qqChdMdb16K/9BEB9jMybf0avEckok3PEtl9y/WFOXNcLi7ktsMuc3o4n0MyE3e/4IBm+vkX4
D4BJ1yWTkTQk2J+gobvRs+QNdr1jDxP74ZbB5rbRF0M+r0/gFzPVB+r2h1YzcMCXfPmDKC0Esvnl
26AISuY9Vrtw2R2Ibo+O5M2o6szILGbIiJCMvXbP942xj8wDLdHSIYo4laK+E53d6a3z4hIj7+7E
wPBUXK55/vLfaQ7noSCyr3tzFtvfL8aXGP+otUNQrIz8ie6xOZpVF8ZrCBquF0pbV2KZDHAMARTq
PHSxTg/Ri7dxNc7IEqSdc82qA1kPwNsFrV6LnxWQv1yGcrj1Lh+hE8TzCh16IwTDETFFDhK9OSr6
MrNttfZnIL3/E/ehMLhe4wbIeBtissX33JVo5dPT4kTJYC52xF0R8sEbwssmBp6ILIohJM9xw16D
D4L1coH9YS4/tAVpquVgVGgaB9NRoz3Gqe7MSfmye5MQt+SBPrT8/ymGK2IzuzDjbOB0P6JUotXN
5xCMH/q/pFy9gfeLKjOKLHU0TX7zkf/NHtp0xdqvh7ObnHp9kPLVc5ejwSndtivXv96S4mHbYCe+
rnVN0hHA6/1eQMgE0BTLis1wPRM3pj9L1EKZQ5HGEAz8eq7GGRdNAZIw/96FbRyrTd/rqTcI5o4N
KnhcRWZZfyBzqtpl41M1S2o6ROEgE0FMzSLqzRQtyIzFs1JQMLliBih+hmZJgepA/9C3ce4td2IB
1Dn0DOgwkpPD2mkfnN9r6SSIwdAXCnib04ReC1lobvjHQfXTaLCvNi03M6lXwBvOyePIT0NQT+qP
Vg0BNzz6Jmm/wPB+zZ8o+H9CDx7ma+72hvR5ElpeKcCmnYaDtFiOeeFwq3A6WILYOrlwOWgZVB4h
jAIDAeghy+9y0TeS7FyjQDgrT5kF72hx5AcDl/3pGib6KXVo7n9gSbZ0cjbAnru/9jPjkXpqA+Cl
s2OClbigafKoWoPkFQZMkzZLm08bDa63ukkWLJs2kZu4hZb5dN4iWniOtkTP65srURbgB1Mu8ih4
oVyiR75EsWxHOu0TsOIegtxS2q/TbAvfwtpIo0OB+n1XyNkSgiljgPtJGRhwva21r3QyZnoMTKRN
zFxGhh+fvQhC15Ji06vBoHV4xQ5uoweY3GdFa8rl4jSmZxzqcAiNoDmgfu2owXvpouRjiilW0sHL
e7/ga6VPg1zeenybo/+mYVbQkTDgef9oMM0QjulILxQOpsxzurA4eNIupgfQR0FxRMfeMRL4xnFf
CF9D6Ng2TKpmKEM0kw3kIoBN99Z5u+xkHmOGuGTijVoVeeOV5IjPwDPMSIKjProR/yw89tWd1alo
wAezuSQxNQd3oLUixSNhtJRUrXXHOmewaUsZZl5gJ/9+Z4E+z48uOHBvod4FOXnPuKCZha6lgMkB
1hCuSiDll78xqCWTmvNauVtExe3c5nAv04FeOuT+62TZPu3OY7FpiVccphlMzcAEPSKgtLygsN9W
v+XweLXIyuZQaNRoMFm00Wcbsmi8ITmgCjX/u2I+oaYO7kOGWiPJLBZBBd0ZQBy08hury8N6sFza
E5KKXDR6EKMW9CEsO6/YccRHN7wviitAM+YZKgXGl+IZggAZwaFGPaqQ5dUsJ+idruEhrWuQMBNv
S0SqLWfxewMOrfwyq3z28llmSNeg0RZlxj+HbNU6KUljgL5Wqg0v30wPXWph/qJE9VVjY3iSYxm4
OO4S4aQ+EquaKEHAmb/fgx6Ew2yGr9rqYUBqbZMW9JYi6PM3uCeK7yBvgld79iCKvu9qsDtzg2I2
8mb5abAh/0pmKEim4yTMyxxy1r21QfCfr6MjqBLdrBpJyyY+CJXLZKVSwpx7utV4IQ5V/a6e7/LP
IA664D2KF8tGqbnHSCqBKeMt5IHgGjuxNAMcpct69tPdy9thaV7x1Z0nAPJBimc79JlBdMKkpHJa
7EuL4/tg0dSNryIMSO5v0+rXe5MKZChjsjAXS0tl1G7uJTm16+yuC2bl2Va0q1XKGOnzmrt+jKuO
XLfsntOpS9mWfMAOeXOby5ktai6caN5vYAqWpJSTUgcwA1B9eJPTHUwr4Tn3SpWIjUg7Ik+aDjrj
vMA82kQFbjx/zMwKFASZzzfJ9BSqvdN6ijBQ8kUHthLIHem1JayCmkHF7EgrMn9eJBSjdzGi2EOl
jfVFB8qXEoj54kiib8u9uOKbHDl8ymDgxLmzB9VKfP8RSVDLPV0ar0pueyjd9LOWrgmZd86Cbj30
dreJdNMHPdHBmuKNPgy/Oc2Z5NPn3e5VVGkzHzG/CPsPd5MsTkcCK477WsBPe2XMF0qjFr+/QYY7
J0In3h84oQVfmZFKs0fv1MSxjkg7C9z1dkrE4ssU+V0eurDON9/tndJC90u3SbCH7QI8uvj2JG2q
lgimgBMs8pIX/NTPEyxrCuNUQkDQyC4F9Bx7wI9vKtzTKxzP/AIQ4DhSSXQyCDAfGiWQfBV+LIPA
fv8dlSAkKaO6koZQRICuEkUmqxTeLIJ4LnfnQ4uDb6ZETOrN/AmNneeIMslC14JOK7xpuTPsmOpU
KWGeMUGjRZn/GMCSCQOIb8YCAUtensLRyJkjSx6r3w+pMQd2O30bIF0MVLjueaa+TZjjZezd2WSC
ZOeue0zWBvFST1AOxI+j8zZ6pRFX+VK6H7IxtbixYq7H8DvYl5n4Cqoj/OZbsRLm7MVWBQnwZGES
nl3vyks9wGHavVy082PpQO0kLiMACqmqQCHcvrpA/DRPXBxC+pS2g0b3gdGx23HAzwFXcTw21vS0
g3MwkKThKUqCCpWdxv+0UF4e3BsWvztu3MSRi2SGPnRC4RFleWcLhRL5wK1B5FVUNdsJo4wM79Qe
846yWocqOsCsuyuZttOm4BA0GJGraNkx7pHIp5RVRTrT2PJ52x8BL7Q62uBGOdXygBx9QHfnMoKq
6T+3dCi0XUvLq7MAjtkHwiBKUd5opeeF2TsB7UU6EZ5CPYsz08XQELzJUNqKQX1olKDI3mJ8P6Dr
0wA0XzoGL1uG4/w/S2dlhjYqeg8hhbPPjdTRYhNMwWZK0mxtcEcn/SS1GF9S1vla8C0Ica6m/iiB
/pdid5HQDh0m63ui9zBFQl69kU6eFCfUlicshRutg+iD7hg8/SOVU8LtI7bL+FwWmfWwJlGbPJz8
H7yDl6zb/tEoUgr8qjZa74aW+oA1ycsSYeCYJQUaIjGqiq5qJxTyyoShE89+sbpaWl2sEWD/Tga+
fXy02RNsQjIipuSDMWmhHckbHDfa9+y6NWwRixgXTIGWSHSbvSk8PbBQaa1wDiADyDE3LVIFBEZo
3qWvAleAlduuyNcT0uYmXmELDeNrxfTiNGI0KDfJna8nmHHmEhUnXgk0K/NHnMPPgljToiO+ieZy
DB/X0Pi9tKb8oJXVGD8Ejfpfqj5PYwbtwL16ygL/61NHjHVmQV0QJ78dhwkBkVJYbJLZza9eaJXc
rAo16v822KYMleM6D9IG+xAwoyDRWLOllLgNA5qdhlIncWJHBG+OMiyc+W9Hd/JM/otqWL52VmSb
2YPhjNa5eDpf7o410O7iIFU0XGh6Z8u9iYRR2ZKB2UGoOLwZ23t1qEDtIV7STwZfXoPtWx9flFfA
GonpGXpMtMH4WUW92WeM5nBWCYe2JB2je8RhGmXODIPFut5H6UBiXkkwhDw1mkBfK1oomunRVyPd
iUZ/YhJaJxFcdgjMmavqWw+DKB1XhVqJruQ/gHc5QT4A/vqVbaJQP92JmizQTOK+npoS7yBbgmNL
P1J8eFbsJDsmdZd996Z/I847bvmqQYo2aWkRWbe97U5xLdzLoUhtAj38L8gHssFWde5LfAdD8JiL
DzKgQ1UKleLPA65xGIqeeYpAHPkSuJum5b52TriJdbWzby4wL1UXtTW99VbdmxPtgT5eqCkYOm1F
eoECYn3Lqqd5wW1aXizQd3rqAJJ5btkQ/6MDjipoM6W3aiJXKbRb//xavmBPI89J5El3195be/sx
y4XTn7Ra47tzVK5OG/DF/gVrxlDQZ1QfsBkf7efIYqrj6CzL4xR94B8cIz4g/DHMbkoKr9P3Ha2r
ju6ThH0IWE4ClhazVPptshsEIcVkvkffujvuANVg/uXrzluFpuRYkkHGviNEJxo6EOSt99pP/oWz
CQyNtZw0NRsf4z2ZYFnTSdFDvQHPgzk1mXH/hxKdojJT8ylylrLnUaQPA+GSkEHy4Pg49meD3c/l
6k28Spum8xtWRzN+GPwCCE9hHWNSmWpqa2cKNQG+hD+51PtXaoQnyI7WTf9gsaH6geau6BfsvY3S
x3UhCOBoWMYGb8jr+ULCZPpOVTZ0A3yZzWIHQ52QXE6rnASTApeYPSqIB7O//bSNcAF5AzGgmyu7
qF31mcOlNv0e8qL0+XepwXcfHQPnFI4TuUiEqJ6ijhDKfXNZAZVAmtDO1RUS8towrf8KOti9UuJT
P1q3fVJOX/jjXItrUs3IcYxwq3OXiwPW6oRqqX+rbnpQ8brOv0Z3jNG3xIA+8o86GjVf5oBu6uIz
KEvxxIzMCs4UzwEQ2Yfr8QCmFYnKZqaN51VM9xisEILXR2tkFNaHLR1KKp+JoJzrKhh8vaB2kWIh
0t+lQM7T5VgC5P2/Uydiq8xOEnAXa3xF/r0gF1LA1gfC2sm/SAK5P6KmZsGb+41dHDtEEXjwLdN8
W1yYUiNqiaBP34w7Wp0/X2qRFXNfu3bO476u3rVaO7TQ0ssvmmXeYfDaYQR6gnxRm/MdAzXefkjU
+P9vmw3b9lIJE9g2Goe9+1Y/nsRDlBK+Gwsf/regEjXBBk7KnaE87Rs/CV1+ACrhNCOyZLf1ww/C
3L9UDz9U9l+uXMUbPEkpi1/dQOhnDznA/fVgxnPKs6xC4p5J4ytytrMUSaWOf+aDcBKRWj2YeKyn
wBrJi4DFiPlebeMlW4MGLIIPkfNvzTaLdXsuN6GPuWZ5sPoEODcb1E+w7eAsWtigJzovXPVfQtr7
/ydgoPncoOQFov7TcB2VftyGKuvPXlmELQZtIqsnSTpSB5O0hxdyTEP98PlF4VG3i+bXnCjjDYgW
215xBEJ0CMndnPy+NCuemyKosFozSbdNe3Tr1BIGhZnehoR98ED7uuQeg1CgCs+itqI31OA438+X
M8H6jEbH6LWZS2/FGoezBgGFyqMCUTwGl6ecDAhmce79hwW6rJNTAa8DWsnUxz/cn///5gmNOx7a
ZpZKgzhro1K0amLJIlNUR/IN3RbtH3kpt5PaFBdjYSzAY5jh04zyiLOgiY6qkPk1h4JoynPuJanP
Hscmnb0oofJgPYdLtVzwxhKz25SieFMg5t7RJIMRyS3CNccq8dBIX8v2nRJWoWIvGif+vG2A747s
WgL+SqoID6qc5LUU5rM1LpoD8B/GGofGwf9XYhYDVHG+MRDEhSWP/ok/xLhtoCKN60AXvyDQR3Ro
edm4GRd57T279j1z9mFDcQEZtwyp4FZAEjI7DoogVAm9LI1l/okN+7JXErhMHppT7ccveeBV4x+H
n8XicTcp2B7Ib2cEwld2BdNE9kxQQKd1tu4f9XyV/louSibIZd1t1AE4yr3EHkhV986Kfg2nILif
HHB30TxQ2otHEzSSXq+vWnGxDePHwUit7/uSLRbBiAlVGk8EwgJMASq1zpzSUD+oZCLd589OV0oc
BlGW69JWeIhbG2FkM14b1XOsDgEv2zWd/vhVKCw/xn+eXDwadc0S4/4Ct8dOWzNTUFrRrgnEBvaD
A/FTANfd6WRWLy5GX7G/muyUOdGqx6hv5DcgUfNp1g2+bTTp3uUa8HHR2kyZOEfc2UMR1OHzq8WE
gXGsfkpqyey5+TMTXSk1uVJen3kCARN8vm0XgW6LqG2jvSyPA/bh66HIfJGyX8z8b+MX+fjUGwL8
2SGMdmDQtbUamwYKcxwAPFCCJPtawl2Vw6w0l1PWjzWMb07mH0daK2dh1INwtYoFLvOLN+7jNVZ9
YY9SbwrwSUvvMNpWgBhbZt48qXDf60sXgVAAKooLANcV1E9eKld9Eo6HpdG3P5I35/F9dazRlCrP
F5gdQilaDrkKnYC+fV46vBpks7NEswQNaDIhxsyrGpFdsVkIbVPutkAIU8Urtc3Ai+DOjXc7atsj
KNMArOtghNQALHn1JhyskBDATMVIkQwp2L+LiN/1FvamBDJtYE4i5MOJeI0M/t/Sn1aoBm//SUnw
dmjSnF/p/DpgiXf+2drzcO7LazBQbzgdFi+Dr5A236TX0ixYQQ9fPc6qdprqs3X1cVwRorEL7Hoq
Vp82bZba+yMtXuoEy2c+h9CM5sApe892fVks+k0kF/BGRf7wbGCDXYghWi3mdiz9/ysqrI6s5Xcu
FgzYIYGLFZbVSXLMZKbg6gZj2WH1DWomE34rwe0/rwkey5/Sh9tcwlH7rxm3OZsqVofyV5jKyUx9
1KEQSzV3fglMaU7JyPkc9TSnOid8UrMvhL2ue5VHZhPMoSoGrfX8SGpBE5/zUarpo8LzTaOZbESl
fDlEwFgcqiQe8n8TrvjB+z24KiZYkOzTNYqlc4aUylupXXjtUEEcq3nDfz8vaq/EBrHB80+xOpmx
h1TQa++GZq486nBBsjMKroWYV4j4znxXyBM6qdqavP/iC1v8oW+oznNHOTw3goc//aiMQ76QfBXM
dxhFRK0IyHnmCX1HHRne7fg5Y7do8EqlAfNgTYd20UMEHDoK0n2uylGoZJ9Pj0ibkKJsvvQ76S25
yqXt+B49AbRmZsNRWsR9jhZwgATzh0NTBWEnAl2nCve3uSnDXXwHu+jhpvClU6NevSCRgYNcaQ4l
oq1RFSihnpbAhJb/zr6nE3fbVmq0BrjtNSlTDhWHr5sZ1G9F2IWgZanAsUoDM6im/gVHCQjsevg3
DuCh36OKF6gO9EQCTvSPi4PYLIglGCoWfFPv5htAV/Z+yVMUcfpN85rKE5sbw5bDDIr7QZu7FrYN
7Olv2bFNLzLlwf3GMUQRNEAFIajHWCsG8Py7IVk1o6G7FEUqAICVMJFxTlkTXM8tCT2rdgfauV4d
XyOFIC7Q5ggaCWux518orm8cFemKf3hTRjU9O+ZHBv9TzZDtsclLz7D2I/gLV5+UColiZNb3oFPO
YLN1fHhmNCR7ietwh2jdMa2m6KQt6ZDQdEDHVjb6Yzttf2exgf7+a6pmLWnAJ43HFE4Q6sJqtvXu
FY6aXxIQtqIBro5m0CHlv+uNNa9a9UD1e/qZQGRWggdzTcM1oIpEavZNRVl5J0mPuQYHybF9Zmkc
WYvi5siHiv+NbFl1GKzO/mtX1jUIAPnfLyVWK2XimlefqTZ6KeYDNigAL+6bmVN7DG+shiGWtl//
W8OqoFVXXT5uL1O9HDAvFsr+FDxdfJ7dAJyBGweGJV35Gfj2pZj7+zFB+rYhOSNlhx1im9U630hh
uRAEong5+WVkxwaCGkdK+IO5b44Zwdbdudz9h3BsvE5YV3mexY2RuOmwlVqd8prvGS5HuiuDtL4r
qftLg3vXeC1Y6Sas6ls6bHq9+9hnKjLzAI6AYaU5EaZ5cRzv4370bNgXuyffzYZnY3GYdRdNIdkq
usB6GQVpB8gJBTn6CnhGesBbAQk1dIOiVTVt8jXgVuuFh8C4HPEAcnccWApK35G3Rv4H1w8QSjap
TDOx1oxdIMVqw55/5/e/+Vc6pjX4CilB3MJdKT5JGBMaZdyshahw5sKNRhfGEE/u0M1DJ+R9dP2N
OG6g4AgD9QAZAO1eUOgVngqAcFtkhwBvyOdXtbplD/N+yN1aui7Yo6nSLh3DQrz0FFCaNfD40itk
Xv6b2PpT07pCLc53x/GHDFt2xy+RxzVVroDbz+Gu+qGlyuVFLH4MrJAWEFPpeZ0rvfbz8h0QwzIl
/3eusuGLlJdlSXovUCY+IsIxsXAow4jJu5t7mWoKdRFXP+5IDQJIqENM2BjpZxp123GrlP3gvR1U
x6an5mUhvlRqDykZWrfM77szuwRiAP0CMte2jHHiV4YuHUC4CwbzV8yEuffteWJT2EDWMa1Qs+/d
RiUftMgYsjMuEqGg+2JcoxxYHovRM+gtLkzFGnQVuUdZKhZHeZ9wkvogYqRGE/wKjuyVSFCrFhxh
RfrTpWdkm8O5nBm2jIMqfSQcKIlyH85douLNVkRQc91P7W9DaE2IgoQ4aaneLv9X2IYL1aYOA/cg
Ute9zrpFxzRXCw13LgOR57L75omy0P76H29U9+qwWIZWvT6VLZoryVTMDp4t/AnVHgr/QwGbHVo3
7Zuod2DtAG+UfAlFhxP8plcVyShdYUcB2jfNphe+xorUVy2AadZ+hrjp7UyRyjjVYp3fBgwX5NIt
zDLV1KU2lYHtWXvT2bPFAPH7zVLiYunl2AQqCLC8FveAJK7JAp4sbHgDXxfDE1oht/aD0VshGN7V
bQsuGYxhHW8wONnvjm9SexJsu+A+yk+ajQUxNUrMNwsyqmeFoIOY1Qm3W5ka6k0rEWPKPzzo9l60
UjLXR/V2BG/i9Q51B99YNKH5LM7LSPgKSRCTB+OsayjsM9jDAhVlpzn+zBtSy3/HOZbQkrAmlz7T
eHfxMSWFxwPqkwC90U+qIXBq00oZ1ivCBsw49waS7h3OfOos86FkF2IqWEWIl5WLGfW+utiw10E5
+b2uMl4053NPACvBKOZelVbu9+lmfZTaHEjVRRIBfC7XwN8b5CmR0Sie8WbyMl+c3OA8rqt5mQcB
84fjFtnBuuB/ytUpYGzQu72ir0ZVJLKkkWWXDeLjFTaFyiM7W2PcWpuFxZF1Wz2wimoyq3VslIVP
7zSUBa9IYHkqi2/oawcMLeoqZMcrQWn3Fuoc6MBUGhPgNpppAvuhlOZFRUIbOGGw2uo3WcNWhb+v
syuZNqxb1OsRA05c8Be+jH84oQXWDamA6r3eyn0KjJNbX5vOlhNHnigjU6CvF/Zy8GFCyhv6b5oc
7WByAkdgoLiQaW1NpwH7eMxILd+0clmxAcRbXFeuCCjxAYYUmkky0Pyd9IDeukLVlkf2NeqIQD71
jmnD2p8Nz6B2UdZ+z2DL5LKlZz0ECMmGylQCFDaXWSfSs1n0iyvt5iPTV50gOTBK5qjlplyeZWCF
YjazH1rallgDZVATLCLLHJU+i8PGoyO5Pxt++7TIxX8Kz0S4gAa34dFPeJsREgubg3deFGbAJfMj
ofUC0kne2SgRECf6a8DvDhiEGSpFrEHb+i9xfGR0YKUEkWdzMqEEjXDyLRv55vAu6H+xOYdwrAl+
amNxwgBeFqGQW8rgcoF5h+r9EambmfVL214cz6KmLrpvj08l/hRSuLAskF1TnvDhhbf/QNU2F7NA
jpO8BOKoFEqbdSoEWKq+OvPqqzHGwVWEB6ORBSpFKznKvzbq53/xZd0xvxMF1b2IF3UrFGcMwY5S
87ZeQGJ6Fp93g6GI6TA/MwGfBr6xfm1AIKy44HfI/lWN7cWHv7Hd7xjpI1x0brlxkhTGaOIIMzJ7
jusWx3lazsn4Ta29Be/oiowwjNRa0lBq81qDp3ZUncmUsZXClWSnz1r3AbL8Pqr9pWhBpI4UaPdq
rTDRFF9TCD4D89vGoiVOh7wIV7Y/Ul0nHpaT/XVW35djo9U1IT1sxNrr+mbwugmi4Hf4PsuKAEPM
ACjLFMfEuCBeb9waB8Y8ak4m6rpvie7jvZZTyz57CQ0ci3IacTBd+yFTmNMNWN9+Ci03S+Llz+KD
ird0in+Fjopxdoc8N5tjVnbTeces/WlRQ9qthqaFoot0c4tQAL+k1fi1oW2IBKS9YTByFDYgYh7L
L8FjHmsJk70U6wpxVZSy99IdI1b6B1WR0H0f7i/ngMvPXROMf5RXcbGK7RZ1RVesBL9+i+JYU9RL
a5/QwUAwROoTMPQ27PqEFLcbzM9f1on4PsRu0m5I5YysZgwvqqs06JIBe7EcD8GgRK3Ik+1rXdrX
uJFlGdurCNO/BdUwzI6id83F5Adm9kL10AG3ejAIRWrIYxqROoWntddqwlx+a0mVWK44JH3UXKcy
qUzVvgcaXUZ+CqLyjbc3JcazgLinb2S5XRuN6K1bO2NKjvqE3FSPphY417oq1KkbyMvU7d3cHHKx
OxwGchYTHn+RYU7ohBRWU07csVdJgb8HKk9iWrXzTebD06xgjg7Tf65g7VxAg8ypnlTqwW+7M66y
/XbAgUxOauqDLnL3C4nlRsgg20wkj5bUdgs6zph5J7UuITvys9lfL5IpaGEKcO6384DKX6e0nnL2
dDNyO5i1nsMKDWOlL6FJ5vzZ3mTj6b/IGoSBk11YmqeVwk7xBJO8V/KN+O1ARLOe2koQqLKKt8m5
BQicF/hzXBUp1FgAMT5H6tgEDec8BBhg0oxbn4Jb1YLGtS2NBZs8vobDRFOtinKhjbLjZRZp9yBT
l5OJpDBG4Sp43c7pJwWSK6Nv5blGgcJO1hefNQaiRq6Rc1FEdXQOZmeR2lFW2vNGu6XCtfHrCWWC
gDpWFGGni0IUdvnEbnGjDAx9tozIdVIPl+Xva4+ioC6tiJPpnOovtlrk77lnNdhIJi+nXrcdLNjR
ukFFXr+wZqoRqHhLLpUq9SH02m7kH8Ds3Yzryl/VKofAOb4Bf99zRBaIosNt6QrnqUWDaz+OEmv1
pGauaifkH7v49bl2gJ2NAeqXGG6kBfqStz6OmENmPlmDIRimEN+kFMpKohuskkmlN6l7ccqG5UdS
yEjFtZ6jCEQxAf/jlrKWeSxDUXoCtULmWetPbZUJpkPL9Vzg676z/I8iFjIk7Uxl/096MPBR6LJS
iPuYCvEDR1nHJYfnvbImidnrE4qIGaII8uASM0WetlVEyzPhEupbU7/KN8TeayfmF+eY7ceVnJXq
gixDUZQoAM9rH+T6N5y4pYuvqpCuetZd6gtMzQxlmNLKkZbWFRUBWuqvNqF7Sk9FSVK1HqcNhp7X
zSRMKr5tuQd2W0/jXkfZ3F0fcT/Mlf4UTGtXyFwhSvmvtIi9EB3tpBfldUhqpgm4HgzFCt0x/xJP
3oCBzn2GOX3mwg5Rk3JXmy9KiXLG19kvPVLgvRqfVDVhd6w6BbB9OnerXPhZwALCRbayhC4k5BmP
XjxxnPio2sStPYX07plno+baEUv1qjqWSPjwEswFasL9UzyDNGebcY1Nki3g4jvLsT0eWi75WSdY
1N/77fpm0R6pxfpeFQ312A80MOjjtbsmA15ccASU80oowIx+96Iar+Gigw2B3eCxxA1ymdsnTnZK
Mxe+uDPtG5J7i3fCE5pGvgwcOaMos+a5yi7AOS/69M+FRRYMA2nFAJA2p/FQONsta1xKLRQc/Z8d
zdLavnHVBkojrIo+hSDXK9Dsn9hrcESrM8+/pda0EaV12GMVfbP7YLniLjqbizrGGW2OYKyY78uI
d7LfclHIZZvJMwPA0eIwNZV2EKMECRvSk6UndeXoHn+C7Cgnaf8HITZaoPr9of4c0nh6WX+meiTf
9a0Nyq66NwLlJ/6dHIY7qHW7Y52PbbD3AJ1LfDzhNpctWRFGDa5/67Vx6BhhStj36eqMoy+qQ/ZV
P/eBiGZ2XbZ6+QxGkyvXDQ8n5GDP/dCgYFcQL9WiP4WN8t+a3G2FTxBn4yefrY6EL+X8owpXhBDS
i1dKrW/vCBps0465nFRrBw6f9R26EaW3ORTQkAYV3BWzBqtuoVVrFJOis7l1YrQVjKwz5pxHbOS6
zLA3eBhvxWL/+av6BYLgjM5Hspr+94fTk8tGtfpp2e57Fj3hedKIZNma8EVN++D5A5rJ64b6uyuI
neMIwoOCsxNzwM2QGR5UI/HXpK34lYf2rOenz6wSEy/1mWTCtbXKaMHOFcYWZdc07sNaQB6GAkYs
+qLD2I5arFElhND0KpeBysBE5sQYGTBb4/6YqhZmYtdJlJEC/dcyegViESB4vbJejyo1/V3PLAki
SceErNHgSKr2I4bgb2GgNmXvVoL8oxNee19QZZNi3AiMa/aLhhO8kYiP+L8jIolZLCvhsDB9P182
I4C5LVgOGu5QAu5TbKBNgnoQJ48Ws9MTxnyxW1fHXzDwzg0bdctA8YHTpHe5g0+ZEoh2jY9rYPal
JPLM6pHWKQlPouYwwhSY+oxDQLNkz0sJS6ROPxkyQDPnXafw0VxBSXQRJy02nLKaOpoE/Sgab3+A
YUsF3v6l6FWwHXRd5yfw5CDiBhU1WQbjV+mW8uQTLOfitdgboWB6PNrYWi40CGPTzynjw8k9SIMS
KukCdG4SejFh+p8XH4A6AyYQC0p18YG/5CoshH8KxpFqHHk/Le3oFII8gGcnKlFBJppAD+C+DqE9
pMY4ySnVMwgKXhDRx5gqZrsrc/NkrbW/GfPAh76FTtcA+EWuCNbeWsqFGA4YX4gv88sY1tUDjZ+W
grjV2+jspwOUmYcNRuY8YAJxgNPzjdoVBVqwnEyso/HeZw/Y3pgCInLVzE+kr1TvSEaYROBk7fUy
TXz1k/MtJ26JkqX0iv2IkGxRiHG6NXSBLb9Vzl6Ycn3jA3xiEJmx7si0x7IYCNbIyR5+N6I+WJkq
U1tlFKwc1TSDVyKuUMYzRtggqLKUSrqhoclY/csEQwJ6QsBc23C2kSY4PfHZkbOKs6sozxXuqK/n
rGZDSlW4d8fVENgl+VRA2yA3rb6aZK3qnrWFEt++hPKhhpijIVrwiPIlRJkwgIyO8UR/Nuc7VgKq
S2dc1ESdL3fbcNU2GR2tUSIa4IVkMXvae0a0aFUD9ldaMBxbMqJbZnBs5nN81iGOF3tZ3KM8KzGG
GnnMVH9kDg0dDdWi7Kkp8LzZUavICr/iFXlShv+gNekja46qnKnnOVwuqwwXyIvrDGIOJWu6HuhY
QLSNi7Xg40Z/TQ1B3lmbWfuF7yKSmvDgmqj9KAGiYNj5BtBtDkjVm/LhAK5dflxqT6xGVPrjwTmq
k4wpPOrFBy0NuXRXbfnx9Tz+sh6E4BWT0GwYNfp344eQy+fsdlOaD/jIJqjRSddJ4IOFuMWhdstr
bRgHwWqV09ANn5OEYQSTIj4N/prK5eF+a1HAYkroPMhNIRR2atDQhIMfB0EGVT/yvuErwkF7PW+6
X23RNyDNZm3ArOL+yojoHLgU1DTLjmNtrwXuTzXlRVGi2JvXfEKKE8Bu6aXHuZF7EEbEp3qtlsA/
eRe4ows57qmi9XI+GOSuz+3C2tCF90cNC2uMbzM8C2KGkB6Cz6BamaptuGeIpMwwSN1y7k9lsAzg
3XC7aC7X5uobz9yiYiWRqtE3W/KTbjN87iO4ojcly45+eq4JF1nb5dU527Dn0N8V1bzm9IgknyTJ
CeSHknEm61kt1l1HdC4hFGP1yCTam3hlpmdULgrIJ6226I3MmqBkkVQXRZEQEMvsW1hskMVu5IR2
KtsAmHyFNyUfWUuBl9FA2gMFYRKDU1Y0XtptbxCnpSf6vk9VT2kRQOE1NYcEhJ17eR2Bcd+MaT98
rUiuoRAPvDdZwwViksNtHgwd5cBJPhT8ETGgRR+D7jMX8d7hpEHoJAt8rH5VI//sB2KkD5N9jF9B
zkn8cggMZDphN/omBJYHeeTWKU37gJfzAbrisXj1NOT6wa0O9t9J81mDrOia1Pn1HkdOF7P3ZobK
vHfRi6o5RF83x6fbAZFCeniKkIPbZsp3l3PgpUE4BDIyAUsXiXkIffOFbgfLo47gKcamEL8QBT/q
SLzTaU0Pr/hjFjFza0Xwn4qRFv0WCB97mYrPNPfftla5I/VDAZ3sVUBElAxbjEah3WnVMnIH46lO
SiJqkF9nUVKeIuCiK27LwDN9mSa0oqIu7Tsa3o2uDm/Qlg8sQ+95esATomgk/iXMmoSeCgLOkAiL
cMz+RHIjijjFxPCH5Ymq2qs2iZNMT7Hv18kA+ptfTDjhmjbvfEm1u8kJ4LrC1iopfdctpJbKPNON
+13A0YawUCEdw899//Lt4t2J/nrja0lJvIbpLBbH7xdERFMUoKHiiBukrEd/0p/lqpptae8RVIZv
qwIBLZQm0zFVUDT+gp0/53+weMApwD9HyxKnK+evv6skiIUWquOSsb9s+Bjrjq+UuMmDUUsCdTSR
LqtW8ydnHO582JzeOSNpsFWyr1juP42UpEj5lMBqlwmxhT7NnZyAYbMvKzwqeYyy/HGwsdYj0nSh
90Fcmgl2urVc4C4a5wfHkmqvJAVB4hQCX/KuLf5VNld4jdBTOo4wIFnwMIhxZ5TuOIeC/7zCAY/0
79AQYkpUOmQ3hYY3nWHzY8mi6YANjq6BdYKthEbxQJLJ3Y7XoCUPLqKLLBG28GxluBdXrFVH/M7F
BS+5PIySsibmdGkyuIo6OUwFlCJK2DYxqPgBK4n2c3GU5oLRM2wmoRMsi/PXJg7jO7HdJO/qOZX2
N7hn/e9lfMcJQdLfgBSOVEQJ5ezwSqrPkYBmrHzxU/p8vMWzAlB3Dp67gglDg/A+w4Q7s5b4/8HP
9qow1ZQd5+UmBYslX8oROlgGhrr6Zo/7TJTWRnlbGeACWAa4OgCvMljImL7kiA/fpHZlGzti1grG
xGgP/cHXTQgdrzld/7jFadyWsjp6QoQ2tmQIQEuG69jQDDR1eznBoxUIWNiytgMJt5biVha7fLoH
IjcchKUlQymGu24ZjphL/T4XSmnSEpntirfTcix+ocIkWDopoqMCX8/DznAnjbSshJvPzf0Zq9u7
4faLIHZ84FOJFojGjnWiDXR2lYXN2foV9HQufVcnpa/yYyBmKq1vVUWyur7KbnnDJoBnB+3CDs7Y
ppdwVKTiN6LDc9VgqgV+1U4/mQuAlzaYPShyRuUL3aqYOipbFBpgJSoXX3IXFYXJ/lcgSIOaK8Ie
d/lV4MN+Ce+CR9qxX4KLoZfz9fiTuPRNYNbI0xPD2/yYdAxK3NFt4uppWLqnHAXKaSxhqhV0vSQc
pX5D5jPhvvZl3mk/+FVxbwOG/OqD+EiIrn3qqpFBs6oaKjyL4sqyYg56sISCZ6qEoajg/swqBvUR
jOMeOk+v5x1BPu+MfnxuJIVwIwjJY3b4tc+Vhvh9128vPp9bkgwgrV7iHj0dQqXq9JbF2EP0utp3
8SJI/sa7kyhI1E9aadsbjYct2P3U9/dr6f3h2NtgGOAU4bh2wOPu+Jw3Odsh8fkx28EauLgq42uK
JDJ/BG/LfQcA4HYfhBKHFMflwKQPilK4QIcCIrERv5fTNQWrPdGIiaQouuNZyPNjkG0SCK5vVwG3
ZUylogmOSK9a6e4qCC1vsjB4+TipXZZ5f0D3N5A1vauzGBOpwGUrgDJPHMunVUoozWpweJUJHLVP
icXFsqMDadpZfUOtzx9CWZJPOCs0+X/HplJGhry5e+finfpIzOH1hXNmV1eLX/f3fNE2WBoNErHL
hAlgUrMpJN8UPNx/kbW6u9lVA9Lj0FQs1ntd4prFeTj0V+LVP75s7UNbaYANRJTi+PpkXaPZRaYs
c1BK7+qNCwMnDLYY9qu+WMnKEk2k7rb5CCzX8hEUeonvXPKN2VkcC7LP+udvTm4izoqGb5yP5bm0
1X5VyPOtBpWwFOg0aTSCcG5AXrAmQ21Lro7xg9ULDa8YjeRSh1vu/SwTAUufVwPt7wzm+R5RCBhi
+s/ULHmIOApJW510xi1qTUzsjzwPuPc+A3iWxyqehSIPh82etF71g5rDoCs02MK1PfBFrHbRXOLC
o4APGy29z6HT1DeRPLHng3w6zdBPLPnqRZEeneqLwJ3RSA3sw/3dmH5y8abvJ14+qrmq3cPGGWaD
BDkXDObnpshnp4LScL+UEEilytRv+ybkpxS+MxGjLRiRXJlvXrLdhm/ORrxTKeWWqwmxssgeI7Jn
vZHW9zE06lHXJy5dO8RG5Lme72f2tC20+2S8ihG6SWJMON85kpdRk1UQcFTYvXkdJ5P7hV10hVls
bGvOwZucC9XqYDPl2lbvWMgRx5Q8BCZhAB+QoWDP2GgiNcjQtXM/pyhAyG9VI+b7X+wEGckRDH0O
xUhqVZIKIUPfHVFn2omZX+JwTiL3fVwb4aylAUG7/Xii81DchPOObUYFledFyu20xD2gbhP86sPp
5vJZrIWSg3heJzsIzQsAvdE5O9dWEbfRrGAF8e+aBbjo7/QaaXQUJIpQR5t7EEoSI7Rcw83yW4k4
QdJTzxyGVBCiVOqEUv5gJycZ+P8aNYQ9QqPK6okqxKEKdhSrqdXnRJ8TXTvuDo8yCexTtbm9SPrV
ZhaZQqgE9fSpC1Fse7m9G1+psbSTOo84ce8J8I3AyilaInWLxJMAbvhnG8/TMPOvMjU5fdfrLQ5C
3cgbA90osPjzKiK2YtU4MFaoYlg9Sq+Tryb9OlorPBCCRXx8Flruw0oPDOr6FR6WivfThOfYdya2
f6N9oRADNHhaE+UQTf3OIO249FxuDtF8EJJMgM0yBWt1z3SLWH0tTvrtFnz0rnF+MqvLy65dfoKl
Keiwo3Eh8X9wwzbKTRKQs9Ldhi7sQ4AfLC1LQc7hjRjAjydVGhdYDaDbluc9oECrlR5ERZWvpzEx
7id2Hg+awLR3sgmTB8/9bovrnaJPB8qoKtChe4LSIuJTWkJHJaycGXUKlYJnRT+a1l0TSuuiMz3k
XKLVq3aBR86x2Kh1CahvDjQYjg0Sv7BJ0gUMMK1TMo8WVPYdWuVQgJuDePqJcRXOIZ78vzzCMsMi
4Y/AsQfyxTpIsk4WfGLAvgcae8ssLftkfX9kjE1jwedqR+fhANG6x9ZV/RoMVEzjvOFKRWsHG3ya
MJlyZ/4fIpR+hIY5b3c7heMWlDH0RUIrYXX1uGMq/plJ1ePK/yLNpvoSUDUQW8e2jrMDFyNtoLlJ
JQ3IGLqnyPB6eqmGP0iUzbz0kznTrIaZ/YqNen9g23APKBGDpkxRqZxHoJR+lL5z6xCXIltCTNJN
sU7jeaZ7x8D/sfoJb4ZVm4NNEykolmYMn9KUsAMdwbA1ig3Wg0t/hb/dg91CvOU6M5WPgqiO+zfk
8l4O1k6/mtbZP3Ufkx8GEdO4VCsXlhQw3klSddyQ6m56rzR1xyhiFFvUo62glVu00+8k5C/lE/Xi
PRpQ+C0WsPj+A9yCyko8wbRQ9bQyBklbRvXcEDCd65wQMH73y4x0qoe/qKPotoQvDgdCRkXBOFnZ
k8Rof6/wWJHFO9t3Z/DdyH7LiXiKbzNjQKBaPNskAgsmvR2ASbwrXOb5MsZimxqVg2B7Mx7U+N+Z
XLWgF8aPruL+c1c8S7PFSmqGb1GK8p987O8hJYmACPXBGeZBplUcZ2ZYKhwQcC5j7ahkXTY7+o3B
e2ZuFUNIl/+A9BPUfvsyPIqg+xFuyYRzoWuT1xJOHg1cjs58m15jIfpjZODKZ9Xm82ruYcTH0v86
j3tFixJ6xLXfLUvK83l/72zROpnxzidIWhva4S96dvhif6sveU2y2dOIspAjCIDjN85u/9XF2fg5
g2PPbhZuTXNf17P9VCsyKnI6dsGp/FDXqH7p+UqT6GZuvuAXXPTI7ePtKyR0NmzdnNX1y4BNgu5/
9NYlSrsRgO9K7ug3ytkfqPuhq6wuLih5af6D4tsgLHEgL6ZaXzieDLBNbZIuC73uFeTLX32ttid7
nKK0rQIgKlZn5UVy7LIEZebPZrm8rXtDCdq+DpYSyVjpZe1QOFJ5PuW8ESyMtLP3/YkDQcygdWsh
LeFwtMHljixAyHqL73rF2ofpP9u4YirVGBRumumDAL+TVF3YpIZvJLIg9RptnI6g0YEev6XGonqL
jw+j5kO4NnWbG780A6riQS1Xkqvg+UjMreHZF5kTXKdLZQW5uT/flQVGhas8VEKhQtrNWCOOsNzq
hBivVjIx+p9dCvEG7Zg40LfL3cg1Ag12Iioj+dpsb+6Ki2jo4HFNiO+AoVSjcig/6DHy0RAz5l+z
gHtdB2cAO4f+B0mtKUyECwHITqVsbrJY1Zf8uYk4MyUaUz4hEZeAOJwz6ez7a5dx60W5JNqTPVJT
Y/ir8faKib5vCYysC9DKhHxQpunCj6LPaJQVBLRnQnATBuq2YRMYCXgbbhhE8AhqEIub3gxkTVNF
efzfTsaGslSriDo3GOEPyC2ymEEECFlUR0Fo9l6mEDi8m1BTzz8Ze7kc0anucVTYp+pCSvmbivTX
ts6xW1Wjupb3fWxTIxypg3QLOC+aYuEDwkFgDNnEVY0Yp9rO+Nq2PIgamwKfTn0YpL2+tqqjywDS
iclKPEw6sCUluvNnSHPj+5rhz2kC4ZotsCrdiatUr3iLlLfTujTQxXaWrwV1MiD5QpZFpjF/Zwnd
PHwd24w3Vi48ie7HnnE8z2255PtKAhPYhF0Xw8D7nj9WbkO/tO17maz/ZrsBnj6gnKdQANgm16r0
OTtYoRKdZ6b4o8l1KqrJ+tVnIPndW9KHlsJIlSvdTXH4ol3nCE1q9Ov0sSRxI2OcuZDzgGEV9j+L
KxIlcPmvBmnyNT8Vu6O3Q/qypocVP7CTGeSQEbLSppJU+CfzTsYtov1Dtf7sUDcivjJ5xI8BV2+q
OcraGgffd8sFKJJDMOKOvKZaEO9GLKDoX3VYCc8M18mNzMJkDDsyLrNXiI1ESghkDBBRsdC8rudZ
sRkfMHe03vYycv+GYImwmLJjsAtxGJ6RK9LtMsvK2cVCrIyVLjjmDIr9y4qgnVgmi6zbx19s/fD/
rfdHNHSDex4tnqaZ40NYXCS/3Kb9ta0oa4JaR00ymo64pLX8gs3U9PhTIhkCrsy93qczUaIy5Tjr
/KKzH8MZDYeN2IzXf0gCwsm/cxp40JkaaQHIu/4TnF17mLN75GYkc3cTxwAAoGkFMHg30Cp93+ry
TQPlCwpoeyJO5Zjz90JYILgPIn+hvJCru3tkTwnEw49vZnLMJTzL5ii97bLu7ArENbSBr6FCjNal
eQyTeOJLZRLFGATOMSB97yusFFDP1goCA0eY0FTsA4QGN4YMawl2pmS9blYi7VZaTZJi1Z1TYMNL
zeiGeTK7WzHYLm39RIjnhvzUR7EtRKLWHX6wHN2F9PseZ17ototTkK9vZATiJdqr4I8sDkPqD6n3
rxjVSu2KsAqSnXDo45hKq5dj9PSd1nWvH4UqlrCUO6x+C/DA7NejnQaUNhOSqnqqyPWDLqR4L+QR
wuq4NfA9LTd3rZ3AY+qoUS1UgIVVRnlsT/pUudWrU17jYpbIVMIU0Pw6jFawsyb5lOs7LJSVr/fo
hQ9wWl3saLwzyT/EWceKXFeesITxGy06CMsZYroAa/K6gK9nHdfenxpjQe14T6hoTNbIQ9ylmiA6
4HLM/Au4Vh5tdb6IBVLKfz/Vaz5h4+kLL2MWnYbcBW3T66e2ARVdoYe8rxjw1FF30cvieMHigcB9
v/6ckXtLAxNdmQMzlkLQV7Zxu6qni5CfigEQL5QReszvpmy81CxCdLIH7TbhSOlsWVsoV7jsni2e
ZDnox1bCHCunxzKGjO/hUujIFlH1bhoIpm5jsZVkvk5pkJjqx5XoGi6EemyMNRwiDxBpkQsieOJJ
dbxhPUbUIVCv7UBlPjpZ5Aqzgm7B+4/r0asn48qF7qD5R+CEuwlTA8TKwtFWJ2T0DTsFV5qZbBp3
scfU+0PqN4fSLZHOnpytpxC2yU0XwUQ+MSm/OYast6O2p0vPOINqOvOVBMlBEODSIjZcADvSneXB
4jukdLMRbhP2GgO7lTa2Cbd2JaAn8RaSEQvmceufFW4d1farVU8M4VvB181WQZWjgnP/gyOMF8mz
lXEUtdKBM63WRHtEakiCc2me6E5nmCdoPS/yKGtReuyDvUcCdhnrFqXjz6K2A+DmkWaKw/RNd1XM
oJ5zNOxVyJ/HgzqejC3G79ym9qg4si5J4UruyNne/PPCGNwir5/31iwZTESQOXlbWF26nAVlnG2T
Qh15K+FC+49PXZk6uVMg8R83EjQiWFVc382opw794g0hk2XuJIQBUK7Ev/UP3lUL1BgqQOglEIom
dRw0Dqj4YxDEu/uGFSMaHOfnIXUZc8kJwHXJFKFIA6aUcyNH/dFgRE2dPPlBIOP8ljNiVtS0mLUI
18bbMKI63YRHqKGVnxrNaTblL6MZcc7ox8v0gVtD553h6njpD/VreK1Ee0v37ytp+7oCOSyIV/Kg
BexAOh+7w3pMYCYIg13q2qZlvOhLVR15U0V92Ka9WKoWHPogDWIlIb0CiZ+3Lx2WPrYA3hrKETW8
GpEOlos1k1oJuz9Xs5pSBRu069PHCEW7Isg8vieOvQJH0EmqP1DCwOSjriJYsndmwEmY5kgy+TjS
HTUvVI6wjVuTthTWLfM0SNOXwioCobBLSRMjVMD2Nh1yq0w7DQYkM1QJ6i3aGZQJmOOxoa2XwH+C
/CqMg4AA7R7go4yG7hdf7qoEvkgX4BKPVA2lVv/vabRclIY7Q4Ip4EKveJvGhd1zJeaoGWNMMK9n
ZnTY9L2U9dZZ/heYCx6zTV6GlQmFZgeK4Ub3S4wgNAgJ/+aD0nlpCg5keDt+KWxm7XfSI9iAUMyJ
06SrY2POFD1ekJzYzu0sjzysLPWPMYGAdYGxajxZzz1z1uSP9y8ynmo0m07FFPBqzH5600iFKdq6
PUWTPsACAgKnC5TSTPFtpmUmp9S4/fvdYak+OEppAre4X21SykuxFPnKuKSLZLmxN67bAQvdcsfG
gjmm8Lf1NaEjHIYfgLQBrxPAf2E6FtGJCxZkcU9oap35sAV1keS7BAHKCcrDHAdnR/uCIz+qqW7z
AswNZqU45mlAgC80Om5PtGm+LdN1E/6Nlf7+5aPL5jNWvkXO7rXQLfs+dTHEqpvqQJOpz7dFTiKW
rOaf5S5iyVruu4/aUZaQicc0hHkuX487z+KlyUFcSGDEL4MOWDeSwTLMDdQl85KXjaOnq+bYpzwq
Nb8D+9UCioD811nm1/5yAbFTTn6AIM8iIKy+WH2bDTZ80qoTpcs8vgCteYo3VinyuevGoTSwUZHS
2L55ZTLdmuaidDY0kWXEASAN1pGWrCc2drfIPbaXCtMzPOQdls3uV85PsynamJGWF5XYMM85Gch5
Krt3PyX1/rm3LOpcz7uejwVxsIeacJ3TXg6KsdjrzxY0U5bPkD99bE72bZ4sTLMhtifJzxhBuVfH
GaZkQ8GnyZhMrvVnCTXXU/ZhgynpPOTs+uK2nN+J4D8eq1QIRl3WEUxetdkok5dlhD68slmtLoYi
cU5dt0H3dNd6tTcrKIoN8BrkPZ/tB8xWi1iFxEHLW4vyz69PRH3sVx3yDoNiODjRz6994ZrlpASN
NaMOla+aV46l9bGwyIXSS80h66t7CY6wV6mumkUEtxlPpMmyXSth1NiFxpItoBRfuSp1sPfdpxNG
G3Rv4KgiW+THrbh75D9snAIPbVcKL5vNjEEVSbXlapcOaAYQNBjnoduHOQcQLk0ARLXZKqN6Gbkz
aaTPNMTgvPYIV5zOK9Rj1+BNvO49KXWPufkFEB39VHECqZu9loaM0LxuDN1U6Ekjo2f99Mg0zfhT
aY9KlUHmJG8NsvCEtQN6Dj4qOoIWKlu8u4ZEJsCWYpQpu4zdJHUT6SUaFIfoCLJPIaLFSxTfVAp1
VwLI9T6c3WuNlb7QJABgVQju6hHbGPNCn/7Jevyxu2jB9wZxnN91PCWj4aogGPQQHM8P5CWgh7MX
6Qg+SOx2jGLLIHDIvmJZ4ZMyEOma+T9TqWyWpCOjM9enWay74ZdjWsFsuBUsbHEa2tlgxf265FXg
KTEglIw89ACkyVr8Z61WBX5zY9JW3QOyaUczk5mYgasP2OtbbvcpBPRYWoAtHyhBjBQ3P4415KiF
/Qb5PxN1tGr4HwVlDXQiv/IXIQfPVUiJfSShSJ70dIGkzAxJffQf/fwIf+JY/MYnia+wj7LtweIY
D96kqLOryPaSAt+rW/L0J3YajE2auqt1Wa42ybVJvqHnJaZZxBjhPASS4KT+55OlD9/w8QocOSqx
zA1gs036m+WPDfjR1oy/hCU7Xs1mNWxuARAJVN0z1YMe/S2sQjK6+rMKwdAByl6YTvbDJ9GfmnBC
iRgO6uXcORtPFsuyHdMCPcbi1BChYzY1JcbkqxQ96jwZc2qz5htb2JTJ7AZpzHZjBAqhBnutV2Yw
N9dcNJMM8BPFnOcDdTVXwEWv1he6/y49r0nlLItQxuQudOkkb1F2l56WGUVW2bkgpS8PrMNXpPeM
4PYDZVkj7livMUjgtcHdpQxeMehlW7y2UCnUyQeF2CaiNgtjS0Dsw7Mkn8ex0pmIXF5hD1GWnbhX
5w1icuSTndTr9oCzx4oCq7HcAmkLfT0WSJlJiYJoOAGtI5I/bQ1qDQGSktaiQLj3JXaZMqn2wbf3
FVTjVr1i/ENVjkBnNps6YegLs3seGGrFhKaIin7zGRjPOeRT/6IWMue3fOKcNqNX0L5Ma3hvv0Vx
E9Cvqo1M6h+fiiQn412ms1IpAkiGkT+iQIONq+Gnbd2BV2lUKwwfU4FgH8HFLZ7EWajgCoy1l0D0
eArRPOYpyRpB5tt25H6VgonhQy7QKBXCHTA3dYwYlV49t8r+8gEBFMPgBxhiW93jPxQjvQg9Epwv
YAnevpbv8coaxT00/OXbABfDkDRozT4FfkiLtFQoImysABexYe8TAyISttwATIreY7Dx7h3Djapq
MpOUVIeGHhIKGbyghSIFlkTt321cSBi/lNl/aEKKWMDjUU09ujD5qmiy6wUrU/18DujvfhWVA8JM
FK2kQP2y4GGUQcOrazHJW3xBjzOogoqYSBE+nTIub7U6nkCOYu1T/Yeq051GXWD4EoR41yKCXBZT
shm9YoZH2J9WXIF0jHNg1XTnrLIpK18Mkb/ThHQtqRbBbzlOEB4+XuCTknHn8t7MiK1ZkubM0bMg
KD4AHLmDhkOi8zBM0yWMC2CZgwiGtWypuM5NKfDVUItuAcOHvOgF3B8LSLoO4LJyV1ym/xtJA+Yq
f89hjZd2gr78Hz9q/Vjz8Bb3F1QsLZ5Bdh+hmusEVKaRICWcBj6U+tO/dThmg7y0WLn6LOgtX+Tm
wwMAv8czV7AMqf9raGmaG52ANEgzkgtUtydzVwFLKFvDhS9SMSQeKeOyowABgM5rt+cUo8ejkPQH
8mBF6V96ezUfHTlFvNSBV3Hf8B0jRfXEG9Y2IubzLY3/7Tk2rpScTX4EepwRvBjnYAqgSnkUumzC
cgUJ+EtY4KnSorurZGCTSSCjwCI1RsnHiHwlyEi5FZN7KXQ61NTXac73hVaPavE4j3kHtrr7EEXW
UyS3fNIYCjGmrKuQNSd19dbi3wTPDgWiIZjPbGoWKAgY6aNmeri+dCM45IfmCNOPV/wxEa8zNScL
cTfusYtHZ3tpotEphjxOOR+Q/3YvlkyRJmKlPYnBboSMcAQJhToVYJjUPuxRRz8potNsjzliW51E
xSTgr5f/I26K9H509V3BR8DND4Earu7KhiF3eGswvEklTxtmdNF4KImVEzwtoVxqWh1BUAeTpCje
qNew/Vta5Na8imBsky439n+SWiMwxk8eTgJbJ8ymfcKMK9o2FaTz6icOzNwfSrz9vPQ0COB5smnS
w59ZeaMyu06v2tjhAHQSWT/0Ase1iOJVPGNFWKhzgszvPam05SLWckln+p7mO8aOdx2BJf+c4e8N
p3V0V4aqvs1mMuKzy5D5MJRCeRwwtXX+B3uP6V8ViVLGlH8N6UV+RXDgJ4k5ovyyq0aSM7Qv883T
Q3+9UOtAgq2yAgpDRYZr710jeyNsMTuDhET8Eszo1M0zHhz219qAGHvggFuRspbmWkQTvsTYy6pp
gaJkufZgzf+x0D929rZ/aLhNKjpVdevb4mnErLN4/ETTgUgD3gB03pIQSTGDG1OAJrO6dArBfSUe
HP5GFXYyneMCujCcWZd3K5n837INt+B6GJDO+UdRHeJUIqyY9YGVeiyiUQcKkHQ4LnPDqn76kttE
5a9qty7ogYe6BpIjSNjucsON+9mr1YVzr0ya+i2Uow21Z2+pczgbKB3BXrsAPr3nc7IKwF/c5O7s
Nl/r15yWztz45G16ocr69X+Y8SQOWOveeq1H1nmsyAs+PBuDZGPt4o/qya3WeDdeXf/Tn2kIgyXa
fbGwZzZUAk2EgejDihPPR/7kfEdDXeM7c30fVTHa6x1brAZ3uVZAujV6WM4a8JM4AjCPCoRPI2uB
/ZKhN4fsgetTXJYeX7QOfa9HSSe0G9+mjOBHCVs5+r2KfVI6wmmg2e5txwQ/srPkjPUZVj/UDTqG
XewzTy7dejBmWpKQjKU6g71gmCN9zyVFUjA4475euqtLxZehjn4XG/Uw8Nh/pjFMYAtpN9brJaXu
tB+XEweDWnYDAeM+Ec7Lb7tq4ApXSfbraNfWyCiMvP5NQm7LP0HRqusplW+BXDVfujT79Ih2bKtI
jfSZ8z+bv/59XpNDN4VyrmyLLCBy2ZTsc1i1XzK/Pf26ElfI42E+P6JU633pFfHMam7Mv/oZHOAQ
h3mfF91HI6suAGMExLnf3oPqYnkUzjTOgRjT5ryVYpaKjRiig3ohwtkuh/gJagSg4zMAkNzw5iP3
nY7m/B7ukI4QI3DBylMJ61DS3+0vAyLdUe6ljWA4eloz2emuYzG7ikI5ZmuTWpXY7dUZzlWMDlCO
mOlR6wABYtUlSo7UK1PHePoU/pE1RB4BChxHmMjV0RZojMV1KnWOkM0+Xf8L3Lt3U55TLCz+cmVm
ECZbhK3hxAnbGkpj4/8gUpG1eTcyUKAmPcwGo1h2HDDfZJLFBHDOvKiMDdQkSUVz1eCIKosybsB+
a8L91MUKPibMvztY6EUkqo2GYtkv0jHlBSl7cqnzfeXxqrzczjFgG8friJTpuS3NXmzh3hpBWMNz
/zQai7HHzeRrT8jNpaF6eRTzbZgUBT/HXmPpIlzptfwKneLav+lwXrkkguPFipn22wQCIA/6bXnz
0KJ+DhUpefq+7xxnL8ssnKokmG+mPjH/yrWjuK5S/gO7EsjK8H2MwixxeIaP0vRZ+h/55VkxcUfN
Tj4hstgJ0LUhwJBLb4psf9nciWBEukIm6ixRZZd4WDIiZxp8cAff7gRD28zQzUNJSnTYC4PqiWbF
Ad6vcmWk+u8mtvbirb6oHVLN3OY1gts1gEAfUrufdGLhV1c+R+Pz50mOFroTLe5o8M4d7fvML0oF
CPAw+32FHmlwfeV3Lnd7Rd/e/NJGw0xekpI1pS1uEx76IzseMIabQ1hPy3ZrcFegrmkfRp8LyWM8
8ShXyNhT3oQJdiXuf54uct/pYrIbP/pRL0iSVh3sF5BYWD2kso46Wb4SZY+tQWWQSdggU0JbsSxp
dUOMIE0XNBn73bYTdzkc0JToq6aZRb8MtsrCpEIWlR4CmlyD8CBUL6WzO9e1jpjqGaUZSpO2WobV
hdmfah7z8tYTwSwwYlTNd+tGHFv9cpS98Z9kjpBTb8aZl0xRB89GyndfB+/xIbu0D0ULLI//M9fU
IUrutYnCaZ6OQHNTYSrxBkp64lkyxQdb1iL/JMe35s1v69fTCCV9L2zsfOQOuef6gJisJ30FxzfX
PbwJyfPj7b1gq/lkXNqdkQVjucpj3jSJoc/ey912IpLye4RoJ/apIdi+qlMXuuekfGeZXx8C42IY
BCZcRUmHV0ZExCtdO2KlZZGiNGaajfegoxPYyOuQM+U8HZPGVYLtQWVYAUK3ZXxMLimeAwxf+uWD
H92HOk+6IDbONITfBiC9YwfDJgCc6tF0T9ED3453Mo6AAnjXMco9NCIUnxLmDlGJmTIKJE2sy7cj
pJRve2HflSHHqInpWdtmfkic42D/t5BjkurV6CrXyrlLt20dLv+k3MKYmpseriaPeC11ZumRYpNW
QCPOgMoohtmD3DnLAggDNAJi8cYQ64JALG00BWCrNMpJF1wGpscC9sHUlFVf0v2FF+xvb1daviEq
2MhN9I5a2xcgdiCTzqv/VPWMye4vc5/8sodM2dbfeZUkH2MwvrGAoY/4fkPzjk2pFFDhATypNjh5
ptHrwKKten3g9Ligls1oHe1NrKHuBrvinlpRJuupSNcX5rbErlF0qwnRD2Hbzui2kQSBdtW7OSMX
m057ll+Bgef/PP3UuaT/SbZxIUKc/jUHgyxTydwT6WYFWsQ7eezlC+k0NbmiRFDklrfC4CMaG4hg
aDu915Ex0IbtJW7SdPUIhrZqeGu5UBgnGyF73fG2ee+z1IR+g36qyynem6j/dZ8unEmQtfdOHh7S
RzSXfNyIby1TIO8uV0Pu8s2AfhXdgpBrbeUOpL9MbbXFdro4AEFlZEJS2Tr03l1GoxbRQJ25RjeD
pp80T4hlYuT7JjNM8xmWhgwzYlOWjVNL0fRA+9aOnAbfff/D2W352HA6IEJBl7uLA42BC/AbtKie
OBsD2ggQHcyoHSLSFI+Rv8SOSTHPxyE0l/Qaco7JbIcxICjjT25yLi2Dx1gD3Di3O9Amh8A6sKue
gdP2L5i5Bmc0aoHh6cH+co/TCnQkPakZGUErzEGyUyivs1ThmriFjTkEyqb0LcdItukgiXtCttBW
fL/C/GMNl0FN8F3T19kCLotB6Pp7BDyHQ8nLFsfDBCgSHqFe1CjZfiZrixnnc2kvfUG1/07IkunX
V1H5/H+Y7AdEcfgoZMIP0qt4YHbMucQi5S4E9tB407WMFlQRkD76U+duk1BIZrB4Aquhd0H8LF0O
BqjHNzKVE+7Z6AlsWGvec96+TZYdCnyNY58zapHOvoFwGRfkzNwUc3iVHo4xLQhMJ+89//aqn1zv
S3hax/mwQD9wFFkZ7pFVpdKgtQC4z0l8V/SBVCxGGEtJBA6Ne4MF0gbtD75QdjAf4E08fEVHMAFO
ilMhMyBiRmmnNAFEdYMUOiro6UxfHsFj+OE9OJqESJZkYunqpuCYFZzNUFOy40q7etUBSz7LA5LA
OLFZEzMO6cVU5BQk2zcjqG2p5r7/Mcd4WUm4W4Xdp6Xf57Qw1LHXntdaq/I+BYpNf8Vx73upsvCb
XzXa+PVVZs2UOXDt62VrQ1UV2No3VQlyMuyRQWPEypZ405TCUuB52s0E5mawsn1i4OG2I6iJvmaW
3koc5eGSbsKp7P5kiROe9pXak1UM2CpJhEn/oRKiocX+zAxKRfW2GEJeDWcEu55RUO09pi+SXzEO
Z97GgYeJNPyzqqWdFkbAUx8LfqitNBqbXe7E5hkg1MtVXSqM/tHgfuaCNQGAVfcOgfVRkpE1s2Cg
Wx5qGHt2oBMDfSu9JatVgeTsTMV2sVAWjGDOKs2wVVNR+CCNHRAos9jT335JoxrVTFQ1QKPr/r1C
ty5HKNH/FAzwHKF/VEocKWdZqGehUJAH46sNa0ppI7uV28gTZZuOHF0aAD/6w/KpSCIBeDb88/un
T3ymtamwehe8Idd0hFypjeXyOvP3di2LnUQMUrLKVcgs0+7yy03DupqtOP/Ucl8+UDroQtW2ACaO
yX0LBm3Mv38pRIko5aptr4PdA+fx5sTug/6XSRmW67//2iU7w9PsB8A8qqwxwfGMjh2GBm+hwdPk
JlfDHE3bv5ha3Cpgv8F27RSdD+/Fivhnse9BS7T5sJPl7EsNtt+rcsHrHoqyTrjg8rWb5r0AKxrs
7Et7/SwU/Efw+0s/jRO37HDYFryymmJW8cWsI3yNyvHwgBOUNM9mLzTOqRcp04fRR6dHxpx+jUA1
2PK1qJyCiHfygrnbzrM2/agdRnGFlSjlYjV/IacqYWHyGso7xvPz3ipuPsCCkw+mSabYONXA6RVe
1MZ2x/4r8v2RYS1iJsY6EuXzkeNtz0AraHyMiYLwwnKvyC4UKDKfMFIymX6OP73HH/0YeVA9M90S
scl5NNRSZliRvHTQZYPr0zHRkM51snieGcfhW4Bb42GPPIM6dtH6V2cMEsO4y0BdX/R0mv6NnuiT
lCi0FKM2T8HS+wQZIMQ834Wz61+jjw6iRaj827Vx224/99vkMuN5unBejY71+BlHnOWfFGyjW1z3
gIKwU6kt+t9ji3L8pEG2L0xj2tTFCZhPeM1bPxdLVrUNORKR7xH+LltetWsHBwfGwF44fCr5yzne
kzcpDG0snL1dL0ugdSXHpEp2D9B/5j/cYm/DdUkDP/H20YRqMx6osoFbGq+OR3dmkk5t5G7Lk449
T1LbwV1gJvZgBCQyKCDS8JEcBCiBC7LY0UEUlnXTtWF9eHBee2Gpf2vGZgI/fdriK7LOgHEnZ+Du
S6SxjrwbkcTZanJ7Aw8JwcI8S69WcslO8OvrVUekL7/7krgw3i08F7OrfzL1AdlodTqI5/cr4LiR
9KbgOFQPxnYIcc/OnFDdURTR2E0OvrWhPX7tZClNRmuRZQCoat6Ts6j4qY/Dstn4/+IWCV75SHLI
dWgZhT0ctZ/2530OhOvbkgbt02IaPAdVIutf9dgpQC19rV97CxjB7aE3cM2SEb1Sg9zpTIUbGX6l
tvaRxYqD443ztiY0SyrVLGdhqhVxUq0eFdDeQM5Ef7tB9kSRnidqJWlWPO+nvtrD3iqsrKW8EG7I
BXjQRYeT/NqrXBttjAj7pVUZUnduPs+aKP/XjFyH9Xn0h3ILC8JUd2lf+V4X8QXoD+Wd6OIVBTnS
q56dYSx+7bSXhdpmAcFTBM8RaPhEL3k8XfkEIyBRCrwP6m6QDYJ6tyIva4MLnYQIvF+vpLXL/mKP
sD0RSAa+jdOnpbkPsmVe/hxs07qrwucEuTp+Z+3NVUf46R/vmjLf8Uy+wmZGz7d0jjjE7wUVUY/Q
DWpQDMGJQidJAn/P4oM/pEwKHaE6rOlxQqtYq9YcjzuCZzG+TDlNSR0+aJwlFj7nbg5FxEE2y8LW
n3cJ1bFkBB8kst2/uIZSAtfJWHu9ZdisdwbpNf6PpqoulASL4YLRqU+x/wPlRrMmcVa3DWG1pzmc
Upsg6NaSPQfd9I8Yvd2EXrUwjHrxgcc5z2px7F8WHtyavHyYfcYw48+mNVuiKCTQf3YGVLxQBQ3g
OE0Ux0KiiqNwcIY5pzY27uUrhLzpoRJ93tWLZ+SgG1pn0OD5umV7uAc94hVaiQSs59shitml47uI
2yBpx6ClrC412EmtiiFnHnf3pgUyLZAbu8zaal37wjOErkfmnnI0Wu9X/PQr3xr0AUSlqEDxGHkB
Kg9fp3hZaYixjYIuhgH0hLFUvEOh6TBuksONxOwKtRkA0Vw7Nx3To4uc9DiL6yDa1CyWf6KYYEuj
mr9xV2rM2Sm4h2VjE2JS7H3uXgPzB77GNIYgkhsDZ611fAarU+D6aV+HwvFeiASO7Mddl3LtcpQV
juHw6jCBusXlpoDydvkSpxuSb5ph6p96OK+YMRKsihbTouXVb7qYCXSjhHfpqAGcZ4/fqPhUX+wr
yhM1G7eRKulj2jR/ddxpO4LqB4IDhTIS9v2easBaXkVG+h4XqacCPWfe3KGCGGbL2z+Ze5ukCzyI
EHSDE+uzK7JfXpwg6LNv1k2QF+n7XNRcYHdqV298zHMTVKSsjyN0URCW1ST9pWRvWRCY6sDJ0ouX
15icdT/d3+elImfGrjmJ1s1lXTvkK+cIzirBkby3cTWSfcgKX11mk4Ep5eejmh+HG0b0qz5wzheR
wVlcgXkugt1WVjYYEwOziNALQW5QDBzh3V5CKPuaIg8loeukH/nnYCsv1OVqb2aqYHmW9ZXseTZT
/bfnWnJdduoyUgSYR2pukx1fgvd3G76ukP0Koik7XBkD2bJPpER02XWcVq1rrTz9lOjWcKx5pMNZ
o5GwBS4/DbRpDePaRaNWDGD3L6gPBtpDLhg/MeAKEW8mBKqYmi0HPJR2fFza6DyqssmE5POt9FR6
FLVX/btUkWeqbUaIQw5iCERYCi1+r+eWnLZAD+RhfD9fbrWJvCDqNN2oGI2XTFMlbcBb5u5661bF
OrH3pbgLjkHbwEE4iBWo+YI3jCDK4BKi1fasemUjUVEANNUDPBnOxb3CX+uSDUnlgicwuBM4SA+O
vlkZfcNItL+TwoF94KxysO6iTcsw4PW8pqqVMuKszLOpBp9TyTP+9RFhaLGu1a8xYmBju626aIvh
qGjS4NXneMUkTBTC5YWHCs1bKqSO4eT/8bFt/fLGqumRaRUEaI17xeSK3Jz/MdJFNfS2z7DpMpcm
Mu49bCWNpaZ3HfizHWmsF7+grCPeCHnwR+0BMh28buvGm9ZZCdYbmQOIGbQKewKKJDI4zdbCIO72
OmvAqypn+X7I+oXU6wcPRAmaaUULpg6HYf4lzuhbawZYMOKi7pqJ2ECuTVpJR+Gr7AokdoDmkVT0
Y3VnvUXfK6jE9U3XLBNUoEP2I4d+apsNqetcjMwCE8VOHqOcDhnOcOWqRRmkJjUvQChE94x4073Q
o3R42uyC4Aq6g9IE5YWmiOP3gJrTR/VyRm4sNRLjUQ37rOxFFBIrZd4d8lO0RZF9aFODLME1E5jM
OB38uqSzfpCD+Zh81bvQSIYL27kA6oG1hmm2ItBB66rc0aLnIFb/7qXixQa8LLYVgCp1TSnohvZr
Qut5NTJ3cEQuzzowtt3xoxo5rjIN4fbLY0nzWTXuhfqzHrRjmyV3+JncgSYoU9g5zyU3NR5CJpXu
3+EIIBGd283Q1WOMO9qabn0VHRCSFvpP1yZ4z3R5TBg/jvLBNb3/5HSdj/RgXCYGjL+Og8NOVYmF
e9G5YU1KQhBSQX7saqBZvW4kphJnQV40LkQ0/ipPczCF1JXxOTVBXyy9ioLqGvmjagkW4Rj6X9+C
pRHGTrsJOSc2LMb4Iy235AqlUGm8GYDasvUdkIgqYEsKIjlio8wRT8ErXH5oR+Isaqf0assQuj6H
TyG3BjWRzQY2fR85b3ISik7OTTQPRMtRnrP1VW7cqsqFLmeyyzgeC3CmsbYxZmxjtbVt0lvzRp2l
PYAtpPHjfeDxYiUr69RWSXTw/eff5a75Wm+aj5fmVWrIravw5TQyZUHQzL/JxCmcCpJ1htZfE6bB
8bm5KltaqZR5Pujkfevm7LtbYI/zndT1tGY6hwdVOpB3zDf9r151Iee+SaJNxQpfcKB88Bu7wmYy
PIHXSxY5l4ObtMHj4EdA4MR0XjbtqPLbifb9ytIrThcmjpmQ1kiysSCpYlcJCWf5Tz+jREJJMgt5
xJf/xqm9Zl7O3Ef72OTB4GsWj2+0nc0rPPg1C9WWZJXXdzOlVw+i9huY9xb3l72osvF+zaWQmmUl
bIMuPpvaKbggWDBuZzp5GQt2j34mHa/NLSQCPzvBjZScyNcgsmxFUvkltWzOQL4sp8VLFqM/8HWw
heWukgsB05jehiNerr1wxQ5Bbu6Qn2hFwLwiec0yV/f2a/YdWKQgNnCPoPQFUVmzvYs/Qh+swNN4
XuWQmYnI1ELoiM5Hp6S1VXKPAvL1OFuvIbeuovDHINcYTIKLFXp7xWhF9wPUSRGjssz9vTXZaIEJ
u8KwYGqQ/i7dTUjMwN0mYxqheknDukDoplVo7hFB31kwiHJzXBMcK/fWGMnUoMQbmfzVt9VYrflk
gMb7aW93GMFxa1YT3bObx0TiYDHTLWfOg03KMpRIN+dPlQA3OjXO1AkI5T98BsvPcKk+IVltJEMD
Y71N+ev6gCDTLkgONGq+z8cu+U0WYnvkXTh9Ie8kQrivmFV5vIESebvclzXp4hLTs0GoZV4Fi0pq
V7Hsna5v7bTz8Yn/KpKJHwgqTxvZNlT41p+jwaYPIb2b7yvX7QwcLRP4Go9/6EFCFqIfzal7sq19
jBjPXlkYfF53NWpQRBch1M9gag1+Y8rR4gsU8UupGzdFWctkISwf5B/7XTDNkAI8c2Ufuye/ldgb
KCqzTiUiufDe481jPy0XdErrEkQiXpTVSTliU9vSRuuqGO086Jcb0EaVoERDwLARYhSYknjNc3DR
b8MHdx7x2/d2pl3vT1SCLYXcGKYabePCkP+yCiBxA7/FYwuu/XRsYFCghGqcj/8IhgCkczlA0gK6
lPb8a2hG51VEH+yv6YPJtD/uRUQ1/cqHj/DWaRrWpk7bFSbnqve9/Nhq2Np7nfCv0vyfRr5+RKlF
cIvGyg8p5FFv1+gkFn9yXs8EPKz3J+JZks8GL4LeMUAbqsBAfXrw3JD2MXbNi5I/dEr4yti1CApS
/gLCYak/U1ZxewkDd6K6kWq+jHebougQnmK1PrpoiMqD+54jpU4XJxP2va+dWTceo7lHhtDlvwRl
sTZ9yhUqVkrnTR1e2qpvKthNprmI3Zh0+sxD6pYT3aYtA16x87TCNV3KgGx1NzH0oQGIqqZPKeMs
Pyrigs7I6M+b2TByS8c7frfnpdddy1cnNxq6YbLliVfsOn0uf24kspKguEywuSs95fFaqqmWXxvR
ildIBLnP2nnC4UaIjC8dgIBtD1NOW+4dYvtwchfIs4kmz3tfGXVz0ndRDDBfvdl0rAuoF5iZ7NE3
f540x7fy2r+ol9gXYgUholXZ44TsWhEzTf36+gybqKi973c/QXajZ3+qEFjJk6DxbLYDfoIHciHH
5GmlDD46SZea37pj7o9FL9w6e3eA3hYtG93syt9pX7X3KPibfi8qtDoPmxtOhZmK8z/Ux4W1m7hu
U3Iin0CYIqwhhtR6BtOK7P24jK9IQZmJllp+CbLYl1TB099t/sJasQD4SdpTQsowl0xYCBEHAHlD
zsJ0i4eW6kEtGt7NAPcX9E47mivQDAEvlu1IofRg9iHSrgQsLe73RIpJIACA2tMoRFnOnC1nfTyJ
eHICWDfv9Cuv58o7X00QKqpNaOZGnydvrm14SpPpbNq5tAuiLKFk5+Q+6fwEuovlBOY048JHpz14
G0cIVbhGx5wm+pVQvfAT/P9wL8FwG3eVEYT4XO0iWvlh1OBkizVxMSKw4gKBvUFpv0CtFgaUVTRD
apS60x2csKvYxsR5bLjl164QXH0SsAl2t/CchSFfkQVIUTqrV/JQlYOKmvJCaX1lJopGnVWBcak+
5WrYvcM10LHpnzRxEkf+Ku6z0TV1EHvSj024Q5mnwSGhcsRjqjpSuMofnuPsvgj2b4Mm4SRAADXu
FvPRiaihVjMFUxL2jJdkS5EmIhRiiEWgfCRTB5sHiFNB66i4rsucRlUVb902SjPlDp6/q7bfb0wR
ifOC7onG++esuVUibbOyA9bWViD9gptw03dUmvLnp2+5vNXpsIKK5FHB+tnlOpgRgT4RGZ2chExR
Pa/WEoSYJpcyCblTh9xumA4uD8CEpVAWPrwrHXsf0SJYq1v5DhP5uB0OgMtRYbekX3+CROzsWyS+
ZUcmaGl8AOtUNcDkHxqwBA0lC/kNWYT2rKip3r2dj8n3hNPJ8WufJfcWeW4Nk878/Ii1C/A5N7vF
WP+6hh40SRvCd1Plr46PRSHasvrSDcNin8UpWXMhaKjSLqp8rODA0+5AmYzfUYpUelUq09B5KGq3
ZAIUu7YWXvxMAwk1C2HIWq9A4LDIzNiC3QqsvY5Nfu7cXS62Qk0Z08qG6snKayqM8+/8M6rdRUI6
GU5+gm1eifUYc3zIgOUKD/jruJ7rlewarckJ7Ml5Q1pE4nveEOSNA7JRcEIsUPaLLUMC3beTDsQR
q53f4Oo2KCP4RtmGWdSnwkqyVGzECgeQUwycpylMdruv5km/FNCUFn++j7RqPaplVFURcmYxTrgs
2d4FISgLLiHVGpmPX3yfhyC1UfZxK4v5q7NK7F4XbiCKqFHNWl2ctBDrjFjx6A/gD0WTt5jV+0gF
s2yzvjUqnCNfrKZ7kCTVqOCCZdLHzYnTaZApySIfPDQp56dSz6MBFt+F983s4ci+m3x4QoSTwm+0
jTCM7gYwmKc4dbKCYl1SUJSL9N7fp8goCOXMtBQyonZF1wgKR26eDMWPGW3uaPCVitl6KkZo/dnC
RBr/iam3aH5UA4TcgozXY3V7PPUYfdEX/89BfUq5p3/Zk9W6wO8C0/jcC/mOXAlQKjs1Y5xz7I1q
D55Or8AFSQISfTSlT+JuXepibbR7ivi+6wMWLEQ5Jpvk1MdAGWwWkHwrN6J7OoUc5NwZVrG529qu
4sBTG+iNYEdzlWQLPLbb4bNdbqgC1GcpiCQTHtorep6BHOF4xC1s+cJrf9oMhz+OvNuHak3m29y7
BrpGBMapD3Z1IbymwtqoCcXxlL2dL/35IGOHvsPg+4i6u6LowVnUJJXBiYIQP/cUA2h70U9ZRa2w
mEU1By5sc3d2+pF4pNSR71RtrVEk+jXkz0RZC6w7mnKL/0nR+BKWZhDxihBfwl9Ywf3DnUiQ3VGl
7sxaLWJz6mWPRR9nn020qel+hObRfkAFRMTvEJ2BwBG8xlV5w025vMiLgsNVsQCWr/k4b/YwQyj9
jkM0UlDJ6ktGdd+2mUqgmq7+ADMPBFjU2tM3Hu8qRoRpWyc9hRv0RUOSvNju0SxRD2wYuimO9tAi
Mpg2bcyPqUy1xNccz/8749i2Hvdf1ll+QRNH7mkLgYClyyArmMk8DVPEpxn1fj//Z8pPKSNVsyMS
L5e4ergl7VyBO37wBwLYjc5wC/nsK0JyUlmhTLqUrPnNn9gs8Ue7C77oQErLh2gUHWI1MovMA0w2
O/LSeIBjZ5w3VDOsmxo4D7DEMepyOUr/13oor1vUUfPUB2uA2vxgtqbFdBatdrwWp8p8j5pXTyWw
ckkF8EPXAJ6zxMyZmIeeLNHflhHlmNDyhbnWs1ReJ6cxvE8OP1+7Spdwn7yaGAfbNKaopHzdujBq
ubP9Y/VczH6FtrTvkaqZxMlw3jqvB12yWPNQFdjQgyvB5Seu6+DU6nSytCMEirtMvz/bE4stRfWQ
4pGHxp5x25NH8n+40DOhOf/tcS1I8dQyFaqMFXY4inbgr1PCwOjS02A30WGu9H7UdGOz9xHx50Li
7hl1B/GgptqWKU0YwbFIQTx87HdjExMFrGBU77BJCoNcnz9/qnhccge0Zsgzv8DMPY/5b2wJ0St6
hNiFFQg89prUhmuqNP8xH1cKzrgwws3/Mso4E3c0EqWVi3pFepPdnu1jm0LtYxU8863bjwZ7Ksjm
Sfmf9DTWFaolOvO84PD+MScfWlNvG6xQkwXP/pRfkPOElgWq4gk8cHkh+4BlDPv+9uhPd6nkBLFU
Tz+J6TFdtjOBKl8oUcltH86rHErnd8x1ueCGPFi7kE9MnS7ZaDp9oGmyPKQYSPmiEH3jSlTh90l1
6MuzMdDVmvzL8Ywd9O8cSB9zPpTH4ap19JbALlHEtHx7WXkXGCa60ZVoeZUng8LgXe+VA+/WITqL
5A0fMy5wVxoZ44kPAbsJSwhWcZamVDjhS23wW8bcmRhXWdKVTf5AQvg0JjsIht/oevi/DeRW7gzk
hurLV7RPqilK54g4BLLi9ykAo+X8DVpU9g5Wwc5lyxnH1SQR0F+1gPEc+m8K4PwtT/H5YEMuVelw
N7xXau0vjYW4BRfUNzO27lWioN2IQ9PS5n8dMoiJDP7jvTwzQvE6G+vP4JtBG4Fv9egYYG1/Vc3R
X2f43NVDepijzvwbXKyrYFN/4/PE8sIlrdhYmGgT7jqtbPCx8JgHo7r3onZ95fB1SvjEqOKI3l51
dPIl55LiL735v4aomMqS01aS8CxPx/yAuJYw2emw36JODE24wLaTRG2Npsf9DpBxc4SQefFfuZ2Q
IZ1dE3ZU60OhD83NzHyIRRI8C07WgFeUqjyBtZXhjedd5S/krBGyVmgtf8IXO8phibCpNWD+mmK6
J9Ut4CAsz7X2LKN3jMXQ6LqFGzIlB3bZ5mMxaqOXTInpkP82REpMN6AXFyJZnErwP+arucfeduwJ
rHMAlRY8rguGbTOfaPpjJMAY9/V4+Vyad2I3kNBIyt7qvWDpC6ZzIJDm7buX0jJmHGZP+DOiQKyu
jw8OqNbNf0VO5oD5wIcGZ/vxiSOuNW2LGsLVteisW1ZmS9laJ+r7DOUxa4U9LPnatY63/Pe3Ffa3
aoaWqWmoIcjnkFxq27tUSYR3MdzwT9gasLzGOsOvzLX6nrn9Qdel/l0tux3Xy9i7spHGYQQstfvF
kNpu0G+58QWFefuWrZpIoqoDE13ii3v2dR3k2HwXqd05j/5FFowFvPB0ND4QaivAwcLGx7RqwR8h
fQH9iE+6HxO91Gq7VcAJKPDBWYXN6oAqU4RnpwcNbnQloGKkoaWMm+4wU15G0rzmIQXatX5+IPJ4
hWkcep4rqI4e5s0b6oBDpP1ibNdHJ8RDWHCx7WH10QiA18OsxciIQN4kKDRdMpUVT7GIqDsMxEvQ
E7faQk27HQGbJmrKo4YMMCaz58yTMPj+lzZt5GY65PNG8RPPjhmPPa6qsB3GjwGY4CXNw5xhLfe2
gFucBUVCPuxSqU747/BKhAqBza9edxbSKm5ViVim6AHNSAES6dsRrECBZKaloHS7utsIPsSH4K6Q
NO2wTWTfjkxXz0IW/Cd8mUl7heZcD/e0atk1placnVZ9Yn2CXvxN5o152LVwOaDcXE9geWMes2As
OJok/fyUsZBh8T5oLhkpQ043B2WZnhdPgV1uc/WWO8z5kzJDYMErgtAwcfyy3/fueGBy/bs0B6iu
1wdw42ZgTyls4SnKc31B+EIa1mH7OF2pfjs1liAwqAqpazk6xcYm7HTfazkEIya/NIy7UXf7WrAt
pKXPBxXGn5lh/kkA8ciC/CrKnPTdYZj+9CredBmmRA1JAwVuc6841nv/MOb6P1zeB+nhx7NWd6Sd
ZAEJuzt5Z7P8p6m687NnhiPr0v7KqIGsQrivDlwcBTbZ5UF7oRj7SwQvjDkjnVEz2edaEi5IMIMc
RJZgniLcNX3uzR9b43LLZt6hO40Y9Gyg9TvNtdT4Hn8lku6DkasP4ujFM2qBMUdAKiewYAgbWnw3
NPQEsCuYshQcN/KYokBBPp13zrVji7xLiuk7E6ePeEol3eGmsMwhVKZDBKz06l8Gs9kwfGicsah7
dFRQzqQYEbGvLJLC4tllyIMNBXzjpNvpPUAScKp1C+mkW13Xe+3gllMdnMwqY3qMA0leirhDicwz
lr5aihePs0HrObAQCH1TGM8p3YKZjRziPbkwXHbLgwZX3GblIAfDy6Imrea6vI1gqAyt8gTN4Vdd
iDduc+5sGQY2ep9ZUZ1VyzdLDPpSbh4Hd/83DMoWT+dGJYxmt3Ti5UISZWE8pdvf89L/EE6kzp4l
QOcHuwsexIkg66Iai2I5CSC0tlr1zrg6/Bng2bfrzBylwOYt6RU4bwNaXuDW03BPaRabplPkcH/A
Tkzyn59EfwXlKjVvG06l7d5bhWfFKAytwyJ21jsK5fuKnqaVJE7DYOCqSt/lfIeAjggfFQ0S8NTT
pVnLrdtaCpKe7M0KPjmc6khuQVfoy5gnG0rxr2Bo71XLVY2hwwN788W4PfCvWE8E5rmGDLom5hRz
/pZpbBBIYfhDbDXqookl8+5AObqBYcfZCIMgH21E/j2VDGQ0f3rReDCf4S+f85waMUAIKWzXz42V
kojM8X8jBX2OtdC4Zp2uCpOZpTl8DKQcTzdrfu6fMIT4Xd8WO3ZmuqLrcNS6QqqDnIX+IuZRDyyW
ev/9F32JkryvoIuRstniP+QO8K4pvkpIffKeQY9KTQPBdxEK9U7E+xNsGd1DdpsZ3XTMaWg0iaC8
D5EcGRVevEXmEMOROEKwjLFC5tUVqMyFGQIY3AbzH9QRjRfjp9EFuueS2ViLRxiCtejeC0r0xH+e
q4bPLx1GU2Yi0rxrc0SDZIYDTQTG1B9ust1VNKQVEgQiasvCa1RnYqU9k0WRy0lMJmWfXnJmxyS2
AxO/+lQRf9y/Mq8wRMwCOVI6/tbQ27i250oNkZE+krmwo2akV5BmrjFSaV5dDC2Lds4MTp7sz9eS
5IsablfmSuGeYuoC5Re7r9jDndNOmECmpF9rVrppHs53AaceM6aEkOImNL2aYbUvCHCud0LUsce+
d/OHKgG18rbE8S7XIBRi7tbGMSVVsAX2OeM9OZcel438a6WKovjeTMQsEzhA/1Mrn667KbueP13x
xxSMx/inW1afTWDM/6cTJLiqs0vQeG6qBTgHCz7kAYghBp1Bk8XnPwdqnv9C9qpFUS5tke8VX/Qa
Zty0iOyT/T5FrbQwZbyomvS2JtIN3DQbWQ+rCv1upeyW32FlLhHNdy+H/FMj6x5WVSFnkJoEx3XC
mYmPKrZLJ2wgw/0zjw5TCcAjr/BJ0UHAQ3DACh3mc+xJbyl6kgzJx04PZ2cL/tKUptz6nYfHSjf5
XCFQgLx8fg3wK5hw2zSgPVJtUuWXcsG34NSQIXHc5yNmUkge0XtIzIkqzRzem+594U3Cj1REagKA
Lrafj8MKcGIxSDgYSIgROuptN0JV4m4xaxUMwKtX48fs7dsmSJUB3eZrJVs5LhSjy7tLT/eYygfb
UtN9nxKyYqlDSYW1vtB1V/9SxUCwNag3WkCQQAwTNtxSVC9qEdg6NqGbCCTu0xp88Vw4fBnT7NMY
X1rw8edoOA8/B03LiESt3TKgtqtelZlyR991H05EGUo0B9GQd2lGJWgXFk81uDWRQnLivWp3TNsS
yhvmMMfbTnqoyhTZvsjXlosXEcaavLO5yBdtg0dvbFyRTcUdo2CDJs8LMwCRrgPBQvXoqh8dQ5oD
Y8OTZg3WKloQMbx7tF+X6pc7hIRgM0rN1bBMUIzQ51LHX5NEHXR2TIv/fzDuz7E8mO1Ph8khsbqI
v8Crtd8Uo1G/uI9DU5zoE4mOQbO771NYH4ymobmcdAD6tL0q/JAylIz/IxD3eczh7dA41uNq25dy
dVcSJ4vN1bBXSd8+aAjKaMkBSDKVMiGGB1L6qHgwu8h3HRK9iZC3TWaFdjc2gjF1DBvepQfB8017
d6AbyFMInx6987C7c/LDsmdR6YpLprS1JZHBEsXbMDrx3xsEDyjEv9bK6qGZ7zrsKOyjhAvFAnEX
lSYT7fMSm40L7Yd1nslbwBgE+8uFg+O1OpBH4AyQ9r7LotcgSmk+Becxcax6WKiOGpk+bbFpE693
p8mgxY2OphP4v+tAKa23Cj3UVEb1/BnhIFDDzGZ3p+B+Pq/5rZqgd9bcnQ7xSf/gWCnQY4H1A/37
m1Fl1oI6tG3dygS7gDYU7N9Il9hPvnDSKMF5rRiZ58N+tOabs9B3kVnAQYT9Y8Njm/qnIw7Ft06P
T6MYQGT/DnCM72ZXSdVdmwqi6VojkneJzts9lgenTzOx5JRU57hlF3a+Lz9ehVwHhor2wAcEvu+4
8hEj+UNVg1T0coeVgj+XP2Z9J3seGqxsJWbcM9JxoYSkTnMsX2dyMKoK4cD+eQ32ea385j/2Wciy
i2XUoRWz1kjv5P5EEKoqB4tscL6eFwNjedAqwaeq82GFrVFrkJHxOsFpXUAHJn5TfKkndGkqkean
XzclrDUV7REoOc0vG/IxvvAkH730DGo2X8u57MmuSFiCWrLDedtsoGdgAW961Tub5NKBbkZRN9U2
Yp1pyImYODcNz8/6LvhZgOGqzgiMVjz/pE8cWNWXVcniJe9jNi0eaKp4DWbGsmiNEVFsGjJYD+FT
TWVlS8BkT0XCNg7N4xj1EtrOzj6CSGf5V9SF8of0RmwNTE+UMtLG05WnLXhAzevsKplld9633jJZ
fl8d1yZ97HoYkEBLtME913+JEFcCo2fXwplLQSAh4Yc2XTXh8ZxwmZ3IYzKbkygIFw==
`protect end_protected

