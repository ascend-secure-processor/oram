

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g5OeUkgs5fKPqN+cBc8cyiee/OF3dPmQn+tPeV2m5UK2zlhgQ1Jxxy1JHLE1+K44sv/wK/zfnl6+
lEik6n4EkA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AHU2ZDUgfciZEJH1drHwAJyE0LrT/UobpRV5wEm0bSbkgQ684XVb5Y3svbwCqGDRzVFMenXdRAEz
Vi+A5fTunYqq0TRhD1qk+YmYyj8LUyTxVyLx5S/C8OGS3VGoN2BH+Aw1H5miInXAixSfnB9tch9l
vxRhTpqwYTUwEvVoNPg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jlV3gohz47Gonnat/jrwtrMN1XRzlpRcF7Z8RnmIRkiqhTEuNSWBYbfJsAyeBD7EmzG5JuMfD35p
56zdNebIykVBHIeKaY+z75375dRM6O4/ydNGqmjFBTICQgO06eyQN4fmgQHyC9fz+mS1M9dyhqXe
cwN3bQvOZDfzgCbJDh4+q0xL9fWP0OSM6VcBwnp/4c+KZSJTvyKLSfMaZi6Sd9EDM0zytbMjUJbz
lZpeUkJf21xk7ShuPpCl5Oyu7K1pM1SqL2HvEyRLRAnRfF/DRS1tHkt6FO//R9tvPN2ruYcmgM2H
+dj7W5C0qBcz3g2whND87NOQXYWPQO9mJhK1rg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
njzXAdIzTvpSV5NiuuiUdajadxDilXKaKR92syejhNZpaeImgNDLzcyjEN4OSc/5bsUGsG7WSwEO
LnmCEyj1rYeF6FkFnHbGOktq0b3kPal+V6Mkp2kITXMdm4zuzuFSwh1LvOD/cGfms5gjcl0MAqnK
7tjt3Ev/f5HeFURCQ8c=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hb/7/duNa1D27pJTf5EUHD2NyjjNn8lg37JfTGy5QkKnbGdtvC5JDcOeALohRg+UVom2rliLKbY0
Fs2yHDIjVL+RIumam2ravgCwhjP6TtfSPgdeKhm23h1kQT9MWUhz625q35W4XJvSRrnUUKIemLq1
cYiDAPa4Awq2YUNrkRbo64VsopYBcym3Nn2cy8++V4/uy40/3nzYbQ9Imnao6aj5gOZ9u3k7vLfw
LdzDgqlHbD8ugJJqN3NLntVMewCNIM+xM/Hvykq8cjd5Z6Y0bVWyTOLZfpK1s9oO76pJvSmk+PYG
PqFhaureSbQqqyMpkrIBB85wm7w5HoLgBRG4NQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21632)
`protect data_block
bAV50Gzshw2XSFJff8UnUXGe5hTMHMLSstu+gTKNQ6Cae0tAZuV+JnBy6H9OIHY0btZHYg6qxnS7
0MkANtaclIizJ17ckv9+gsqJscABfXqw7qlUJzAmAPypOi7njz1Yok71hbopJHLdvLFRTADJcaMF
Gm2dD1C37o6e/ZvOEFXGFsfc6MI1kFu13JaZpcrNuyhT+WKVoAmsRbqZNao7IPSx/yWvb4v/J6Nw
I/AQKUfocGJ7PXoA22xqKeWv29pm6czmn9+im/Xa0Ti0ktKRCYsawimaCrDVtPuVPTIkYn66MN3D
ZjMfuVnKyAo91cC/FHuwEfFh/dI4afFnDR0AF+0Y9ObFKeNBtvEmE2frJrf7v6kDN0yoZniYrt+5
xtKSvsFZI/yQCT5mb7YxRw0s3fD3beqV3zgx51TOaWiQCrbBvZn9rMyP7UyzbK134QU3EIymytWc
bZyLIsD5lX3oLq+3npJDSl0dv/wHTxs4dLqJdG3pyfDWhGpx8ya2qJQPMysJYzilxmFJjMbjkJmc
gWdl1WaMSaKhIiy0Or/dwl90Ii43+bPS3lMtNXEG+1SaostPKyIDA2hWzc12Ti00/tfMRedqeA1d
nj3FRBpHYLN/9CRWXD/jVjiTeMlz1Vxfszvn3Zi2RISmKa6qLJ9iDPAY0r/0cg5kCAJPlddIHR0V
aYDlNBHgbRiJKebRnoKd4Z7YYwYl49GyPI8BKbV+Eyp7lJe8uq3ScPP9KhFQJmYVmlQKIannQlIt
jlUogteRLsgj/tzkQy1jkrMnBWCucWMXxKoCcQTsW9SZBxzILhHVfF8wwwWhJIwhyZQ02s2IJjXi
vw0LOl/NGceMLopN+AgqLWeRqnB145CgGRoGjDdUvFow0pa/BU9Kz2bfD/DHFeDNFoz3fB5/GW/K
Gyg89UiR2y/o4vSGXvZM/5njFptGp79iuS+WpaEVh4D6kDBThxV84Fjhg5PvnYk4YfxzWfZFGJfb
NmPNXjFLJcWFmk5vivUUXlGupQukLMBfIwtMiXqWphdSiX3dXaJfnIi6gT8SGP7sJl25sK1iqWZX
ZlSKsijanprUIQaQ39iF6CfIJsV6h/uiazGfE5dveAaZQ7779XVen1s7PgQw+qmEm6N/3srVFuln
WuK68Nuhc0kE69ZAdQK9edD/5NxkVr8DyfCwRkqBKrNV5Bjby2p98EkAuEKK14eNlIlQzq1IOuF9
BSCzU+ordeSlxm0INBDSHKNP+QNjRDFchrt2Gw21seKHIa3/Ycub947a+mo2cxVoMuUxh67a8ItI
EDY14vZSlKalCuYpPqr2LHPZpl5ejDiz9ny8Zk1igGFXLmH7X/z8s66g2OC0v2VHd12ocTFR86pv
M9AQT5g8oe9xiWSv3+B6+oc6qjZgqPJI7v4+5LcUFKVJtor9L9q5sTfn9t7B9pmEzcLYYeddsEmd
fEdS3xt0jkh9xmE3oPoocEbtEs4vBSMbePOfUpvbHLf73GSc283pA3GE5azCml+JCbkY1jiOwtYg
1vKs0gdV2XjKYbdO4W/DME9yW8LqKd/xuxVUTvZiuFqHht8aNRHqGVSa+vlXOAvRJYAjivdj70Cs
Yw6PkfsvUZf2fipHMCtatPu8Vg7wmHoCj9934P82Z9sMUrDl8jLg/zOzX6h6H/5qAP8Xdx7DIJrp
z2r9g9sY2FnID8OPV9JVJZvFWEXRKPkvIL5KlRSw1m2jsIr5Kgeqgzc0G3KZF75Laq4YhTt51+vI
ZNoH7tTQm2j4ZPU98L0jqV+lwQE7iMm7GUy8/22toLZtYA92Jy4yRiL3Ka/VWw+7zXsfXsIJoZDe
0CoJEucRklSRgW1atIlJ8I1WVNo7LfPFUQmcRQgu8dOKrX7bO4xqsuAxI5eMFXx3BhXw2MTZTMWw
tBembdHWx1CAXgli78IfbB/yCmeGXfuKEDJa+ZRmpJmANsc4MaswzKCX3RRemAXEQMUOdMqx0mnD
oiPtVaDk/uhdNLxql77QEJqsRbZ/aYmUaCOytu6x1DOPj3X8QMnsIu8W3ihLxYEphYFQ0w/aMkZj
IXBW+h2rIP0NnDKC08KI6qHLiaoO/GvpVsOZuA6yV9TvKJwYAGDoE+Yec3wDFoCPgxqlxyk+fNxr
5jHtmBLDPd1kHJQuel/XcfMJcRHdB9kFIWRoC2KEOppVoD0iJFVSSTfgKLgRgmgqCpHKOH8YwshU
lsKtoXRt7pO3MiCom8lqggNp/IGEXEobg8PJJB5xI6LDbD7MQ6CsQfE3Z6UDJTO303wy2gbngai2
1kjvHdBafarg+RCDq7c2TgGWwZhwkvCHVdtV2DK912bunczLr1MzmQs46jSk+RqAKLerpIFaQTrp
eGYyw4loA4BL3vE/ehTqcLt71pnJztxjHRuXXEVelAClUrW5PPu5TIQ7meNuHLrA5tT0SJJo0xQ3
eDOmyzW8HE09RQ1xrAtFQ5EEI54jN3D1+8ZWsqFUH6DwamRRwvbfmda00S+h9qEov/8ys/pzbfj0
ClorTZETkBrTE2e0w35Xk1a5Asa4ZqmChH2bDn4OPhm24LqBXBBfpcoAsqCOBR32ilVuTBjsCAZA
aANxhlSIkX+0NNEXDlBGPO/ngQJveV53fIcv9jovT/SDhJQb11HGqLjYPHdHWStpU0L4vgsMAzEJ
ipTpehPFacmqPEDKEknnbpm5u3yCU3KwCs2pSdhEw4rZiVzScY6ctAS/o9yELHQ3Jwy2Zd76D+zG
gH3CxLGL26H2rsrlZVPuX/316OK0/FtZqn/hsgIB0JkpNrPXFoufuu5sPncJXqKS+DwWP7Yr/499
kjc96heL3o6ltirnf1SHfnyTDWyuyzmCA8W0OdokFWj0CpIN5rpdMnDESqmZy5w1mdfl0maH/lO0
AT4hvzJ7yv0Cj3Mh+jz2riwAJI78I22h0XVA5fNmlfn7lPfM4Gnhxc+Qw/uJ+3geStdQnCxQva+2
0Psgj06jVBpZKYZn09HnNnrSBdD3mRsRLCeAM5hx6+9lUwJevbB+EcoddXjVroH5bBa1qwdfak8m
QAf8BhBahzcw6Mbo0/AvHf0jdozCAL3NY0QHqt/nXimPQ4ZBISYUR+8IbeU4Zhm01YWZeOBDFN5C
oTItN+jyCSp6eBRrYXb1BmQxFyx7CJjj7AV+t4KcM1RVXlP8Me/k4/5w1tUiYj43FXeT9ILajCYO
7m7x+yQ1DRCpSRV1l0mCwcdk79bzSI7EKHx1XFxD0GKRuWydx5HTzHzqZgEotU+m/9ihzGKX7pTO
Cbek6cBwBrX+DumHgBcpWvd1/ovXGDiiBo8BiyqlMvknvFbr44dFSOffWmL6QWK+zuOu1JxkRdWK
yDWuhYFXNNUd0tueoffGpOlrZKr8bK3WZojdux6L0UV+B21CNqRORhrtJzFoBoHZ4xi8AvnyMHjE
1hI5sEjfqep91il8RtuAWg1DHboCyaFcnTCSiA8cxP/2Jw7ndsyW/+/xW7o/RfSJjkKd34I41F3W
boKxTFTkb0K5HPzu2XmGKWFLO22o9BYurmKbmttc8/8sA2h1Q0rwUNykZ2DPrl0uE2jJ4ID50EEK
Ol7rFueSA5FCwq52N4wzOv88mCzdT1fNe9pC3FaxEvmW60JGpyshlIny7lgn5n+NHZxp6uD5GvBD
F3LWbTDNJrPTnHrUI5yrzsV57ZkAKIByQAThDhavw2CVXcEUAxb1cElhdDJCsb/+r5mJRd26DGtq
jtL4fN6LAp0gcO02UqUbpA1W7HbkVNRkbLy2KxCl4nPeeV0v00zVgTw86LQzZdUC/EtKqWAphiH3
pGHqGuoA+QgxDUbkXWDimsxqjHeNWrbILtYcTEiGaB/5J3bOl401Y5YVBVoWhlVY+xbqYPa4wTOj
c7fbV6tjxC7fqJVc8u85Ok0i2DhZgkngguGQk7wbXQPal2j/XOqmPtQSxnkVEgh0M6NCWxgTE+Dj
C+3YDn6Wd3LNYHmwzUPUJY6xq08gwTj4OHUI4Tr6JEqo2RmP0RaVaMLLwm+gHd0PiBDD6+IKTLBS
qYiQRMfyyTf83TVY0bP0L9TFNl2kurnTlESo7XinCxBE6Sa1tpVLJoZPFG06B+dddiRD2zWtdinx
/F5FKKj3ajeyteUsVnd4cPreVcqZIt/S6FUI32vK9RlsVxXNWrWXGTGiuXv40bXEcH+/3+Mgxi7e
Ssn23aaybZhdtemEyDOGD740mEaeRd2EDhSBSYSvvR9opL/iOb0bRO+RT655zoUC057GKdAD9xDn
ax1DqGw6NggSqLefRf/sCS+YQRLMdVN7xGyKQu0DTghO/1oeXNuz8CDyTTZV1cmysDi2wdEbAYsA
nEP8XVP+HkVMaLKJyXUkKyhnowzXafiLkdNymx/BhnlFmxibglDh9m0oCSwdvMCfvW4Ezg9tSknT
RQYghQ2BFkaWOb9is0qHyau148sxGFwrPGu0QInzOA4+5djGZwX6KTnA/vIxkMTbH2p249k4BwXR
f3DPb9b2EF1qbPaDOrJMcxDc9kKRPW0pSKSS/CrwblQimtIHVJbxYW4OT8VrbfC32OKg77FkxA1L
XPb/l3Bbefcrnh1ZuEQSgAz/dmi1EPFwepWa24wygAVpH9HIQLte6LxgAON8vzYf5HFe4Ook0oha
s8TU4aszy1XCtEnbTLmyqxuIjD1BMj7w30WM8NkF4gmK4Yitw7/p1oxDg6D6p/0Jx0gpgU0nct8T
rqVJNss/rPs1zQJqygODS6fSEcrPpfo2wUNZLYbnkC0N5Cf6RtzvtrSG84d5PVAOCom856wZ1w25
oaqejZL5aPGuWbkk1RwYtdO8S3RKxl1Tz/Ek3XJjBkYZFGJmrLFCVCy95UPCfDYEiaU6GaEs5euY
sJECpyPRgbqQLGvhZth23hb7nKURd8z/KJHulBGm0XWlbNriNbkmPugYcr+xqVvIBFW1jdi6+N45
0cET30Ic0AjKF0kGNzmgyxepIMtejRIjUXaWqKP6uvNzbGBApbDwwtF5WyqD4KL9vrvqP+c0Lq5x
cGG+N7pjmEEluJG56NNNYbo8tYBd5qicd0CCFlBsFv3aZS3Bchv6CYCNcaIfsZoQNhwUoAWrht0L
b9MogemwBqBOt1rErxIpRF17LjYx3EtsKI2Yusc4S62rDLuP599EMUulUZSQWPZAio1bd8xbZMEP
JsOP9pwwXklvAuqjZDK+krOZWBk0zEjdacLB7VmqV8wTfuY9kJZT/oc1YeN/vV7QJTEm7kO9FkMJ
Rl9VDKm/UvpB9C0PYOW98UP/Gwr1uSIwe/9ztpi1Bx+IcZ7cPqo3Yb7i371Q2Vy/e1btzeBPjGw+
k9bVQqHj2c8joH0jcVbeZxw+eVs8XmiVW+sjBYMN9/gs0h8trqSDW3DxRm9tLZxO1/RCO7QPwJZz
5ZAreEOBXrxU9b5yZhMibqJDODhLRfcnzyVsDNBcU1B1pppMskrB9mJXIlOw1CVfHCwrL3syCi3L
oZU5Y+EwNRm/LVpG2A06MU1qy2niWlrbZwzyM7MUsuqKOE/2EEIIuOB8LccRQTGwy6MjuTUrfYqk
KaPE+dcKYueOr2F70ypdyDBsIglecfYOYcJbc83Ntya7NzFIYQQ+bAa0oPQkW/TOixvGmNHHq7Uc
15pbNabovRKHdqy9dioOQWd7LeOGuc3yaqqE01IZqXpl8aL6oQCe3Z1T8bgaalNEMD4tzrIZkNgw
VNktJsvuWZ+xoVWgjbSwD4lHqHlgZdixJAvUAesP+3sTJLalK2f25Cckdd1RGis5xlN1WYTxCZzE
gW4IIrW06i7vbbefsMg1PlPPEhNAGFv4d+P1WhUpA5w1Z92ZH6AV5cOpYhGgxmd++lLtK0GbmB5q
5EaJIZKw02QJHPbZuiS9IeQdlBvNoYBejIyRvZO7Kq2RGjDbtA4RKksTSrFsMqOUUaiiI/dYYgYg
aeM15Mmi70YIcVzdan6M0qiqRrak6XBX1rfMSWU9uAt2r1jjY2xG7JKcM/zGaZB/WP6IoaTAn5o1
c4CCmELR2pRWr9NjRS94Z/WG5t+12eWO0DnDw4/kuj7Ub//lQnEAoS7okXmSMwH/Dpf+sJCGt7WZ
iA6ySE73uBVJuEdLH4UYuPV45A54mf7dnb7GWwWchJ4al1Ropp/eDugeF1Fz2HAA9gtmY1kXixpb
Vd5coK/1ryk2XVnvBJnry7mpyAcKZrkXY8+0a6MqnWG5bxZxUL9lqyBS163s6/nVBxY51OChXzad
C7dTkT8JqL5jT7p6khKd7mnzykhP9SjgID1E+zZ7WEkhaG2AQNrD0+GPGgSE9rW8u1Ag8D3U3nJf
bPWolDI7hb0Voxs+oZ/6DbRqoovfBklGtQJoV530WP8BIXam2Vw26Kjw350Awec8uFrZTFLClW0g
Lp17RHy9JaAhSdG3s2M8kDsJrVrhNSMjFg8YuihrarMqxZDMfEeqsMBtA3tlp5T+S58/ZYaHRlr8
AeF+qcOVG+E9xnCOq2LZuXqHsuWke3AkfhD2CPPEL7iRxo1Og892E51t9WnaCuVF6qOx+U6yLx8W
KWJHPHGmdIA8x8GgSIipyCbHPJRnz69BBaGwQDwOy6OmHK6d2hV5EO031jXpeJAgPNOd3Na5+NbS
x6JHAS+3LeeZ/XrfmvW2fzsWBv2eVMQBc2Zf2HJiH/U1i04AUP8oBv9TA2VAqO+xR0hvcAVfeN2Z
sXoyrXdBL3EJTr6NyMpY2JjOQ0ppgCKH3LXJDEXHVkER+sAcYzVWALs92BGosvfaaI/UjVLTsany
SUaXqKIQ1E+slMO+XNM58kjtHDXxW/ixP/toBy74nVy1fGl8f3ApaiSfidm8c65j5wXmZeweg34n
yHAouiqr3kCo5kXtoMBdSs4zVV/pMCyaljURXGDTQM3uvEws0sU8gBrTdyIxf5/Gz8B/yybK+0KY
K5iyk4r69lx0kQORrmV8R9ql/31jpQKdxJvvFE3PhkH6aUlL3bDJscZuEKaBw1K/2RX5I3fgEv1d
kGGcVD5tGztPos0zWHvw12KWu+L6YBchBs5Qcx9nJIV8FkquTvSKpW/0wjqEZk5UT0oJHNPNt2kN
cDiXBpeXT1QmcRWc2Si3EHmBuDfH9vugNIvv8lNM0lOb8z4tR295PsY2tL8Kuk/bl5AOcak+bq9f
RXcXxM/800y6cRhwujnly6+qe3S/UXu0qmVc8cIT2RoIKsLrQnfUKvsS3d3cYr2q/I0HFe9DUaL0
8bWg3rB5nr6vnYxGk1vY5j72U0++VdfsnVjKqTw1ULTHkt9iszHGn2zuYJ5000sQJ1l4iB8MLT6c
O+gZNg+HSoNEPT1DC9bIno83O4yEfLgRFMf9aJPfaxOv9tAlPMa2HhD1ITvNtLLZlEjZD1xZZVxC
oAD3zRbN1KdXMZPiZPX99UcFsT2pPhwESbHbazyALM4yUZrPNSnqIb0G+FHCiBNzpp30f+5Ag8yQ
iv7TLHOZaujfJjfxxoS+dvnRuTsBrmDsPCDvVYfnQsF4od7Y2FaAGjj+XMvlzIq3dBZhjMvVVDYL
hyRFsbZyucexv2ebtvzOh7zkFvQlT2mkL0uQo1m7Yjo58y1xQMB14DmChYEjltIj/wHUqpWVnNyl
95ki7rE/Z/PI9e70nTbeKoW6TBbH8NX+/qLwFI03ILJzOAHVU22CjPAzSkxfSh8YlvdMLFvCwVC9
Uzm69sX2hdftWAw4SVnWzlnv9DQVy4sBc+DsA1C63MASb9g5kg5rB+3TFvtcvDXKRRE+kSMiorOm
Mioi3cBN4IyvNQMZVvtEBsIK9zpurbsa0DLv22kNSPCoohnZ25zAR4a+DgCekOHDn7wi5z4oeBj1
TU+1EKUkF86DtmBQYjhJfZ70jr0a+lXiRfHfwyi0owpL9iDLpksYZol+XFF3W4znHLQUPbrqt93a
wngn6XtPP/kCG0oRLjEugnrCMG9mYFfhft2w/bwvQCMGqQwHx8mCcqYMg9SheJARjZ7nAOpE6cMl
z9CUEpGmSHAURk3FZcSzBK5Zkn/qrrGPHYAb6LFojvDTRz+OV1g8dMtd4YiOqC5Xo4I64SxEDblN
h1vPSMfPzaz9vfr9hZCqKHvsyrttz0x8+Ezj3e07rrLWpCNpiLG0JCkVJ1jehkDYiW2ouIdBTYpe
pyUnoji7zhIOk9Lv2ZJVBwrMCzu4O/5n9IlOLEQnHcDdl5OsSH5LssKiAln9NWB+Wpuhjbf+ZYVX
aT0LGAmB0b6F3J5YQ4OKnal81HnO0by09Xp/W0tsaSU3XEVP3EZG7ksck+A168e72OxI+FYCA8pK
D8X1Q/giB/V92X7qCcArHsUARq3bOfg1RLDcMzE9l6n6s/HoO/2OBLPzCvPCad2cp+0rW0y3Udek
WPwApafacuLEFG013mwsZglvdo6iNV/xbk1g0ApbN1KmKafwR0z6zMVMvPHkNiuCkiLMFG5YgSWk
h3PymikcbgQXe9zHGOqA5cQ1L4INu0i+OwKaGFHLztyBwCoQBcOAH0pPr9mQwuMiABzYUp5xsil/
JMNbQ8nTIQ4KIFqN/a/XPvTs/GexFI4adE+HMF1LfQEx2RjjxLvqthUAA8ZRruXNxebh27ouXN4/
EnUOMoRllI8AdmFxn+AvPkGe5B1B05hNEhapBTK4v1vGWSACNKxlMdAD5HHWVKfE70AqvZyxxvBC
LiZwNjryS78Tmo/N5oVVyAz6h39ceb1jKbwxcZ9O4ws1llEHBeCKjkik/HCi3wftBV7vPuEGITbb
UvQc6eWBlaH7oIkmkL5bvfyrJWyl2+pUqcUtXPgBBZ8H0FbSAWihTKECdBapyeBw68LcmxO4MvIA
c1RJKsNij8zg3wkfqUMohSoYfYVlVi9AZETGHyh8I3x9bBTgc535ywQJioJlWzO9k8Ad0mJ1SmP1
tuznO1IxE61wLQowFxqQ6pql5sWHMJaTOTyIHZKO9oJkse2FhMcxv5A2loAm7a2JzlxX+1tw0Zys
Yvjc8PxGF0c+4Y2xJofBXhX/hqLUit0UCkVyYqPnADwtTfArFplsp2CCb6Lee6DGl+RlHdV5CIr9
cjjINv8LpKzKl6tLO82GtMGLXnjR0MYo8BjWioipVS6YDDH9/QhXuvoojOKVadKDxcH14+B+1C3H
efNJGvAQUXG9NqucYwfDkFDiBbJqvytBHiI2obAds1vlGJaxuqSmNIgKknLEclRFe0ouso3Wozt0
mD8gADPgwQs4jyh+Blrkp4ohnpN4L/MRyX543Eef3g7H+5F/T6X7mnn022gW1hBY+73Lkud1nikk
bOY1bx1H9BrzJI8eVOiGdlZCajWmxG4VohrUu7h+9KPy8+g6nQnItDjnsEJD6JGre35e8Ws/Riwn
3MQ3uCfPdj9F0gYdXFGkU1SIGNzkqfs4kFQokZ12ovb+bgUrMQ0AFcc5BAlidUKrRbPKD1X7/swt
/Apky9Kdh/yWTakwklnh0m7OHLlFuhWjJNeC+QT8G1RuSBja7Pu4GlRkWUPlQnTOfRsSR8pFSowV
92f3mbsiLdOT3Zprm6SUILgsLu62OA2tBAIQQOoSFGBr9KC0fFSud/36WXybxayw5s4vi2AJhSzK
AbT6S42h/AmBWsFL1Op5NWyAlCA3iktzrLTxugbqOUTvboYBLfHwEpUrtVNSMzNewITrZXOHrSWr
LpzXFx1X2cG9xACzoDkbDPZeU2qTE5wLjmOpZDj5ooxPtJzqyg5Qf7yIgaBuIPypKJoxL/TpIamA
WtABm4wCntNihnDnn3jzhuc1weab1Q9JCxEzghOuHzNtDeGnifUk1Glbrf/LhFP35PhSrPqcTa1O
BqYmVThqKB7UHa4iqtsWqrcMsK0c5ymVph5VuIJysQCARIJZtGU1ejLhq3tn2YNN8xTlxQ0HHOci
RjVwfzc3SFx2sWYtoOwHnrxTPo+Hjgm8XG0y1Kl2MgHffSHiPg2MTc3uo0WThGpuRHV9qJ9fU6ee
v48F642ArQ/A0eKO6fGtYCLRVQxrNkpD/+3Sp+QdCJrjMskOunA8C4gq8mjUHz/nHwWE7JB/8YmJ
fFew0awD7Iq31YEadesa92aPQxoqx++h8/kjxxVopYc8hLgq8Oo7p1BXqxzyI7z/3X7+rQA0EubX
M5gxiLxtiCx6UhJcgI3LigeEf4NhE3Fn/hlLxbIvtRZqnM64lYww0npME0W3KdZmIZULmCDc3F4a
VH5bJ69jVNAejIJcYEhFRiSFQS2GCEkg2uMz49Hud6DWUwoMLkGUuSbmr2+6jzT1CV1OKyUOi+8z
/F58j46wGDLaBuxDH7XZrEXuwfv62e8DGnVxkC3Y69FfgwO+/W0QSQ5cMUN/sUgfW+WZgMmdF50Y
rLO9uigFc2814WNx2PQayefaGE2/PROr/dKEJuABvx2iTyLfIJWFYjnDREeWmwbhR54w1mBdiB5o
gde4vNH/S4jnAqXYK3tr8lHCmUwD3fuX5gvJuVs2wr2jVvkA9uX6LksP3WZ7VJHE/nRciZr7EvmD
DCKTb3ywgBT8CFvFSuhjjxUQ6EaFX0xIXI3zFamSR5qRYxiZivaisT+IuAFNVlTnNk81IQzsX0AY
9LMiJZoNVFdHlWyf/DBhclHlFKgoVTzwVpLs1JCg1RIJHYDjqtPvgL88F8zGDK0BKxWDoawLzl5S
FIEZaCOOSxeAkcm4fMgPbwmmfMXigkSGEjNI9TylFUwjhruD/2imZGo+9d+q/XJfvq9MhfNadOf0
kfwSfsusyAV83Qg0RM/JyE+OSXRispuhTwuZt8ZZRM76Cq61mYDwVIZlXaWNLRCWWz3lqR8LMLHR
VAjCl05xZycKh40XvXs1DIZpRJya+PHJfcys0iHw/L2TV0K0guQLXCmPq41QAcupQmrAup39RnAZ
s9hWKtG+/6YerDMhUIGTVyNaWH6J+RhM8grnxwSxyIjSKqqX4jnGH6xHIrCSCRbm3k6n6HSrbX5j
9Uf2J0jLfudYlVu1GZHRD+fSDJkMGZiMm5R3+MES0vqE2g4PP9ucTNkVGJsG4IY6Rm785ukOnv0D
wdRA3hnqmwI+iAek6qY9rlyeTgYLAc4bnQl2PGF8SYH7Cfo22KcnDqBhFWy6eo+ZmcQ78hJ48eHD
win5PoYXZniF1fXmK9neUTJAv76HqTWsZcq0BcAi0wSwVuInfkG4uO88GhWUFM4Vz85aCPs/wW03
cC+0xPo0DU6g4PHSruJDtEPmKMvi481HMdFsq5T6OG+THYW6ALYgx0NN3c/ngP4BtbOulcfu+vPG
piQ0vwk+K7nbHuMQ1J2/QnXz19EIFoxzbJNAaI5n1ci89M9+oVTOEf9PvS+gLZ3YW1y74CWbtXp6
hfbOvldqLp472TjxmZvXWCEuY1neX2Y/2vC5WxGO08f9Vh3hyyHA03PtOCYfsDpburMVvzPhuRlf
XN46CY/83u1dbB6xnsXCaMrtFGGcE+WDhdJOQUajUh98MszVPPJTjD5eSwVwLt2HKeBhm/kXekBU
wBqVC/yhZwFSPqCl4AAYOeVeQ4v5IqBuNbdt9GL4OsIlpwnszN7EGx5UjXqbYdTl2iI33QHLSqYD
DKoOZMtokHFu7F2bRCddseTzJfFrkCA76OMZZu8lMMGO16mhfyA6E0oT8s+2ywsOUhnTEIIqbrHQ
AP8OJ02oQhPJ9ZDK3zFM2Nc0vFyiJ6ELRl4zmie2Xxe0piFUqTMK/0ltgeuRUX+3/xuInSPwyCTy
idUZe7esKhYLSB8iVdMyq5CXbY5zJrtPlFWmaNHYGrTA9BqW6ZzbbGu1NoSqI7j/lggbr3DovHEm
NXg4cDORCaEQQudLToVhkIFf+zafuwXHPqHVmoqRHCM8yhp5d1aPisEF3MUNP7VqzFiMBOVy26aU
zE92cYss0XAdwOF1QSN+iOsWak0I8B2WWEbwYPU31a9Frw3NGSFYjTZB0MygEraHvIpGzGECNSkg
67skv2MeMvvKxSW08Md+UYbt3ZNbZPQWn9X/N1OLPi/ipWIHk4hlkcUuUbFMtjlqbHSccK51jwdl
P4K8Pzth4y1tuzbvhHlkbl2+kcbiwwcR42sGTZm+tu8VYiqvdYJDhe3uX+a8c7FkeRXM5ORxjbV9
8I/6cj1IFQfY1bUwHAJDvAEXu18sQcv77kkSr8SDHub2cTgooOHSUBan6toX0wl1JsjFPI+kVhWt
Pq+bv3QS84QmCwI9RXH0ZFbBq0N7nJGlgbyqeMsH8ncV3QhVRxBmFevE+oh8W4esakaA+zfDAflB
mhNCf0vW5RMEI6kXUCuXupXfcuFWayVCYqv+Flf7koPE0MU0SmhRydy1kHXmOFktWiFjSvk+d65r
v9TVg9a/RsmhESxyuv2VC0+g/A7aEKgpwv2+UY1QxgUAbLJfPkNC9u1C6rI0w2JwT8uVVasr6hwm
w5qCnAjdKLQ2y1T0SJBQal+gb5qo07Lr7cMoxknO106i5raShsgUAuVtZCqjsjvV4wi8eVXuEGvK
HaZmWp8P7r3YKiyIY66RBERIdnOmDJxH5vxwZVeBWycxXv9/5aqtyc+bdYZZb7tpiXqWTtl//Nbv
oZVWTble/eoKnfFW+YbewrJEz/nekm3qmOXbEdhvwHrvETlITNBRW3oMg/O8PisZ/f5Q0Fa6lL0y
ZJazRiCTXTxCCaRWoyWQSKxzhObCO8L06J6Fq5AsIun7aiTDFdV6Qgqrd8A/186RO0TGo6bwThmx
dXLpnQ5ohaDSODZg+0QsFpPljv1JMAY6CQa2K033VuFnFhfpmDza2P/Hbr5SlYjQOEAfMgJYD3r8
+FcAlgClU49L/J0tfCgj8HPxWdYmOVrmIWZ9KfddH8WAG0O2kDT0uMMRv2//RQb4vlL5gsDpjUba
pjEaKrC//QW4CJ3OqwDEb+c28EgRMMe4IOJ3UhMzelUo63poS0nmRR3Gd4N3B5BozhmObQTvnKRl
gHPmyECIV7qfC1g7ukl4BHcaZDpImP5V/egGiJ3NwzwxNPWQiLE48QdhkORjV3TVM8BqBdO81453
97c2y+Sy8o7JqszDZFzcOo2PXCSWIm5z3+GGzw2Bxvep08s6Ykb0tZXQRRUB0tUZPmOmqn/PCDB6
S9FmjJ+XgjccSqP83SxzyR024wKC5k6lbUSYhYZlKAWA6JFV0QStXTqC6T1g+36+xYWkWYuwhh5v
OQn8uAR+VwTDk/FTZytxOokLLYB5/Kaya3DZPz+C0vZZBW2u80UlI19VPvE2u0Vols6Ow3WlNzdl
4HZuTszFB2PIV1Of0bMSECsYQAIqopjFmd16eLAes+pwjKiVzWeW4N1d8YBWCMvCvtzFRLP5VkC7
eszyz+ILYE43D8ZPrgkdKqH8Fi+MYaxuYmjgDu4K/+MneSuUqbioduCUK0qpexnnSazup8PRMkpu
2L8aIpFVby0AWe6IkGh7N5Gg5H6V8QahWlt/6vCtsydvJuebozt14CBYPWP1zaMTjBE9cyKqvAER
fDPJsMBp59VkoQJ9eDvQWG0Udin8dYeXrRRC6P2LJxov5kRcaAM/W4ehW07Z22oebw4pUKDteCIL
AP3XdUt4mQZ2VCfN/hibnkDLWjcx5QO80pHVPMOei1rD2ek22u/aRdc9VhBj7/+7JEJH3Mug1dLV
oTR7UQs8ejxyTts8MR3ZUzW8gXy8RFXouHwvGGyvvHzBSWsYCA4guWWb1f5kamlbgYyGso9zqyby
fEbaNnYs85NHcnNLisSq1v7VOVPhTdURJrDnbZJdlqB0by8anJXa2vl1tpAcZCv0NZptzfwVCxf4
EadNh0+e/Sl2rOXcJ2a8nvRrnkg/wxBtw6KyjpamIPBCAjg2hwSJs8Yx4AmZa+UdKXyFOvCj50p4
pYaudKeZbgm+qN1UljPK/pokSnoS+DyOx1tTcACJyAUXCzpeL58jFoeGPiw1dIkfX2Ll0Ofs250g
38MTcMc6X7vnsYKI1GO3KAXvnHar91iKMA5y5I+xSTdDv2UmM2lTRfFWP6DlRrahiN6ntNRLVgCC
XXZDZsx4+qYoetjuGhfHqtIYgqddwQPhX6fGSmMUc6UvL1YDPMfIwPh1mx5d5h0oml/MTa3GOplG
FlpO2ZLRJ9PZmPDbFqelY/f/HaNTwhNcRC9qeKB15QhQAZqcCTxb+yqqLECTsvxztCTbjGy2CWtp
OtDj8lsNIICsEvDktiDKwFCk1QKb+91xJzhx00FH6gq9MLc8nsw3tsOPDr5N3/o1WhTxDruyxJwR
mnJvaq08gLvrMddtKLt0tbhQOI/RWD4BfrRUzahRJT/VEd7VtF3sZL6kd87H+IoyQgFPROacKo1x
l7e/UWBNK3sP0R86MDdg7x5Tq0QcejvtFjIhtKRDHe/t3ELq2IbDo7fGuIsfwsndJHb797zEg4wL
/Kel9TXkH9cKoQQ9tJU02pFEQ+VAeKqdtBSWd9+cHHdn8XsaTyUJSi0DrGeUjBvEF+tlHRkXAAqo
GR8WSEPn6M9F6Qi/40CN9MpiLv5Imbyt+Nmn2QiB8gdwwABB4q3HgVbQVyhaNAxbgLEXqlP/AP/c
PBLH03TqDLVJPZCQEg6oFqyDoXBHBqys28vQFHz9doBRH9PROWeATfU51YtqSysMJvvHkxRkBXGx
WX044v3iTsQotB8oy/ommwMgzOz/GOGFTpqmJdfkBLpS47O5v7rBSrskvoOR1DWYc+jV4OqnduSj
KXPIjIhl0lOQa3TDotl8ASp4VyIiNKlOUBqCbslmPN4iNYHwydAnxzJ7Q/56crKh8LJnvnDa5GV5
SJxJQe3SCkPCczfiR9s15Lg63jKnZRunx0SjxBsMSriRbRJUBt0SXtOdfX9mQfVKX9/YXKroiHUj
2Wrpiht3NWRcqYFGKO4G29+r1WSbkbLLV/DHedGY6RqNaEK/8bAmLfAjA3lFAE+SuWYSgwljA+mR
fU1nqsUPNuM4mImz+o85U0/OfhMPx3u8LDGgUZJpRqVgZ9YfhNYHbc9AOq4HbltkCHRKX7lF4E1q
c5XaymjAshxRwxPYLrKheME4tMSu/QLC3wf37iLruPPwsCt3D9KtYNbqw/JcZ601qtDedAMfuvpm
HMUxo3+YTrB3I/wjVGCOSl9lZ8XAJvKn637n6zO/gkCL7OjanhBPdLI57fJhFRH8YiFDX9cf3lfS
M+au8h7Y08GqbDzYcHH11FM+GFpbOQ5B/PUA7DlOwpaWMnTt2bJF7ZfTYS8AGQWHDeXP3vFaDVMl
a/jIKTS9QoleLSjWGqSehVkY1ekoHRk2KFDfx8Da1PW6vtaXWL4SuWi3YfwYQq1CAiF6g1B7q6+v
lOh0EWrtz5hZOlPgNxV6DBQJr7eMINYOwYCeYQ5AZz5nReSiliOgley3N2YyYSCqXdedAUF6kiwG
SPWbHAQo/xsRPU1DcfTjGaxcCv+5lWSxC4a/Ng87yERJym8p7NmpM4wxOVhvBmTDioss5dwllAA5
kqaTIjz8+Jgm4JG4uFQwdfGZ1CiS+j+jCZMkrTRiCTm+ZGrMkvR3pFFIzwbHQkavlqVlEKGP2MFk
+goqhbAYVEAMdSMRYx8wAWrh5EFbiSHsDRXqGRtc0DvooZd/Cm3yk2aD3zdrZ6JPaCrX7tbRdWZt
r8mY2c3LanVagTioj/3CPyXdkP8W/YmfGCV9irwXUcns/2G8RNXaf67WQ4myr8QvW5HIwKOuBKZ2
mvJqWdbh8UOTGbBV867JFvu87DlzFnuWxzrVqq7XC1PM3SAqAnJX3NciXrQBquNX98oY2TrD93nS
SpI5kUvxouksYkoAFZEkOJsvf7tlsNu3wUNTIthx18UmqzNFCbIxjp5HeSY7hHghlubwaJTRlif6
+WPMWMBSJlVLD3xR9jWH8ZiDjOHC+e3Xaax5fZpAc+pAoAztkGAL33IAmyMf2Zrx1YXV9/Oq8sLl
x9cHgo4piGDICEotfdOAzIwmxYjaXCJfy99MO3msEl8cmgaHNBxGH9mQNiqy4iJ/1Edw/NweUC/v
nGoX8QylJ1/t40YOlLtDEUbyU5Zc2Md4fwUVqAmA4icezd4UE25Xzs71GzLBmWN6iLjsHFiqYzvZ
PRhn4L/GvCtnGAuEg4FBKWtfqxaZ5KtPmib3LXUsBadFaypkP4X9dssJ2njsLN0ydQ+uJXgdTpa9
0a3v5dLy1iKRpRTJTS1StMMONtV2iFYSGoepRtgomAn4DPt285NdQF8fBjVWci8oBVqUsUfpnZM5
kN1oRx/i7QKGf9+p1sZaWNgBsz2q/sH5M1QckKNa2Do0yst6Hn+Q4RVBvqKWEP120BWEc4/1xvLp
8OCM4l1JjptojgUahQTJEnbqHzo+dWf5ddd7iw8RE3jPgzQvHkqcZ8mYVr3Ld2Gk9c5qjXKEj/73
+aFjhELbthkdKiMooDSM80SxVJeAH76X9/aDJT1tI9BxaszAZ8x4blctzRgwhBbu2jlnfvuhS+V1
yjL7Zoe7XcY+oxzTpP0YkeN0EDBlXjPjs8CuTrBgjIfhgLFBLl1eFFidhEt9wH6v93FgfaP/WZ84
bG6Vly91ZNKLE6P6VOQp9Qc92wnoZosGW/3pgDOU7M6qwxiCip/IAiHuuHiY2A1ctVhfZtHdy9hn
HtApf2RPuUEaQQW3VyDpvGhpMpGcQzZodIsC4CudIuXmvdxyDz97EPBkmYYTo6GsP0rit5fwbQcM
kiLTMbXhSIIwp0ZNfttVYwUOpMy1/1WSiNXR65CR7l28g2Km6fyg7EjFVh6WmFRWmQulVdIm3y6m
wklHvWRKW9Y39mKgRJeMOnfOdrJDfMviHxh1kbbvcpVdvbH7SJ09gibgiOEsMarEzJKCtd8kYo9P
lv6AOr/0exOyB4DEa63UQN343A+QFA53KWnRBGE57XZzK20hHXRiDQQlJdnAR1oX9tNDqUBtAB7B
QDjwVpJvN3T6WuTRunpxuy+QCZ15KuVwWDHgNFg+HRcDWlZdDf2k7GVcQfYIPt+LlwL1Y3LgK75q
WWEl8KdDCSToYnpidtUen7ocS7XwyO+cQL1F392JVmCCBdMfJjd0MrA6qvKPiBJ2+NsSq4VsKgzi
FT5LZRFXpDuQ6OpV4asOiv6/DcDBllHNEHjt459sG7kdOClVZcM/x9b41JJ3Nsc7xymoj7KHAHlc
g1/qHH8Lf9+csJAB4ZMidxlB/s3Q92DKz4e7pU54xHM32Vk0vuZmt31EWmEfK0bc85gAipqKasis
7ILqFoSHodvr2mwZmnUs186iRCQScvFijE6yBcsvq0uyzueISfUlqzqGM0in8RQMkZq65XrzFUJw
y5CE4sKhSY78uqBKIV8VLcmb9B0hAlI6ICmGQBytXJwMiIED5QkWmxyUyibd3fa8sytrx37bjO6m
0Dc3QIClgM+xVTEfbsBhV7TDEZs97Q7ImY7qZxAOt6scectYq/AJ8vld+oo4FIik/tTKAmev3r/O
MkhN49fGOC982Z07ayzBED294FDqhZHhxCGrra/dGF4Q8Y+GPJyz7404KRSeyoGpMIAJu87u7S4Y
UYe6lBRPSPOseQb3vjKliROIsncmcaVL4sjxG+ZGrf3u6I44svlYQ1CdwNXC0nw1QPZR2bUSY9yH
up7AgMC7KlJ0BD5nfB76Dx+jq2/isFodAcjBxTB0oKkhHpeZKeYAz6naxtpZRU1diF+hgRGu2R76
ROiN+o/i+XB1wkst99pErwo7iThJ66wsNtFRqemuoowWIDTy7dlJQ9Dp/FhsOh9G+AQBg6bQLC7Z
XFsmbJ8c7dJkmatpPzh7fbRAEKwwiVSBMhW1CLOM6YLs+i785jxCrvuFYRrH216lPZJG3NYx7GrP
F6xKTIpI2HdJ1BcpOVFu1b9j1TSAn5NYDUzSzZe0nVoYOkv7gh6ct5rBCRppncaxvmtYn9V2WGLl
NVxh8YisY9fISJG0u2yiB5r45vpVlplg15Dgon3WGfZ8J00QkIOaypunCby1BqY6HkfqMxIUC4X/
zikfGzgMCDDZHC73i41aQFtcPVdUD77XtA16oFuqgQ5Nxn9dg+IVjwjNDNvqBpWx0S4Cui7jowzO
7iHLt2EIErrGbq0zsUFlzPVbnBTpKLd1R6IpJqQYsp/z7/2hcULxBC41kqB3WFgWYexmFMjHaF2h
s3cSMdIxFXLxke80wrgHdAQwEXIA9KX9YOjZ3jjbhurXK8rjtTzZeHOhajuu0GkW8BPbti7L4OK+
EDEPvygyKexwjrgRasVBn4yqP65V28zqNVy75Eq/aTrzO1vERD2xCBUGeLJiFNLhOj6CmtUMwhy1
fujcbHz+fcLiVeN7eYrnQBsg7Zo/1OGmGbX5eeG1T3WrSC60FgsVD11VsNPOaPnK9/9HjSZe/cjL
b8+aYs2KxwiugYKdu8RFBxZeD6BSSofXxgCBA/KmpMdds5h7sqKcw3NFHzZlheFkRee4YWYbBSpZ
JjneAwr35o+iuv7idyJpuLvAt30IIEyPeYOt8M0eluM7Mo3Nytp/r5GPic+wTguS18qJgtmdRWLu
Huo5S5tPB+r8dTReAyXok648MujH893Alqog+rHrBxG1e0KF6ig6ozEOT3fewexHRYDPXIwYun/w
tdLtUHA+Vdmuu4R1O0IWQSQTL7bvBEJplvGyvW7vlT1IP6BTV8UkokN4lD17QBjZAJo6pBVFIsSY
y8RJQAweLukWUI1IImn359cwgJ43eZG+GAxDAGnyLPle0zn+AQ6yYjK4krQ/EGIvJk6O9toHYjIo
UMvWLlLm6VpWssUWfXwnH3iubyjR42yLCnUxgdLXJj9j03TyD4g26FF4nSTiQ3RfKHkXcFO6pQZC
Kb3ctW0+eLxGw17Nvnb+1Pl0A01ZcGO1Sl1f2wozUl+oFLcPrsLYJoB9V4szhsWIPQD3mdaNUfKM
sxiJfTkbU+DdrlowhEDYuHiQBPhIPWrUmdcBJtNoLbBwfVGtnuYUXTAQh0Zx5iM3ZC0v7nfu9KjU
cqS10HEPwmaJ0ck8VbtZ+Bp2YJVkmoANIxy6Q2KWByq9WHVubqxxupk9VKxcBvHjsCWltpbiW41E
rxL6IqL8xiU27eKCwE/0dWOp9mE+ChcB63wxhLcj+PrlnawVeMzszeD4hJTe/olLALLW24g4ck10
7jpx8aPbdeeIjgPD0jFjatC52j6zwYOvKMGUSVmFQnuwc6UcD9/AGmRmWwo0bEdNUrozW43HC7xR
o8ZFcixkrB2+He75Polgz36T63nwZPaQ5dF8tSY+gZTRsfYGALad9DLShh0hGvIZDw5JEVI9zkbl
iuL6UsO8p66EmztM0qKChc0giYI0RGLsHe8yWEFbkwja6BnP/ZLELWW9cdqcq0qdJbZDYF7nNrTG
hVYQkToTDH/bMMKdiXREpt9XUGwJPaKbKeAtNcMLND8KdxlYST15qlHRaMfrH3FhxGIStq1cVh11
KgfwlWpqhmgwTwkGA7jG/bUnzQUaajqgp+qRksgjQGNicnxcof5I3cT7Vn5tN4FsLPl5Yb5VFOID
JkelB7GBhXg29iNEYo6Yjzv2bu/xWqZXzjAiwZE561wFmZP/Hj7GfEWxRbiYZc4GZFEPc2AQJ96x
SFr7Z0ne4TM/k5Oo/RbtVABLHFqJEuvn247QBICVlJJOXm9l6nBfg9IdpwFOEsKVsVgeNYwHmije
UnRR4+fkecxkE/qaeyxHvJ5T+PHsO6B6+9fjQ747dkRUfb1m14vDk1brPJBhAK/0WoYU1NBV1SAa
uLPNhPguc6QnFcNPQMRNJf0B/B+XYxh9vHcDoGK7xpIQhXpMS/eQEk/gP9mFUTbR2axB1Qr1kB78
IBFSkU6S851j9bAvWnbqmC0XmjzMAFS02mHpNbkyhfMsILHuC3Vh3nsKeNsdG8uUyc4G+27uVh9K
paUTpuhKBDjyMLtsbce/dYR9+xhz8ZphdoCJ0ZvtrSEa4ux5Y5dYv+wsQbl4f5leCD3X/uCtmpxT
CBtCGLkV83i1mQsqPj4tOLeY+b0iOpArYzZtxKk5v3HuDBaT7i7UtIZrStGna8+fAoUwpkLRTvVg
mX93J71vmZ0k2e9DxAKknfmSsM2Q7ZS9prFZzGoad/hFm+1drMT3Aw3a6UTBWcW5MPMBGx9IdOC/
cZo2u9L3gMcBmXZpG+IOlL5YUO5TTYcr23hs8oq8cPskOhUaPavIJygflX6vwTpFoGldC6Pruv8w
yLa0o8CnI+r7o9bF5wI+5CRAtDtjOR9GGYEULyvQEQxaFF1H5zlJBlAld1YhCHEfO4coGTXbsgry
hFS+rMWB7e30qoaJ9/ZmcZ5fWVNomnNwaQXWMaZ0W0Ni8Qk1DEILetiUbjVgLT/SlQ2gtLYxBOut
EEwXpneCN08Yiy9tEC6mTb7UDSeJANMiDiL+6nBJhkebJUiL8sF2Le1+nLWox14d6Z8iytb+Vlmt
/yftfUcKM+7vseGJHV2y5WVsG3QSuMRnKnaJkJhc5QMoaCeahKz3ywi9dE0NLtBMk9VAEzCuteDf
W8WwD1MG8Um6Y5ocirRTQC4LY6vcW+8u6UEKFQxyFaN4jRt9FqCRALy6dqPBWHIqpGONq0XdAHnj
+o6DqFfFVEdvdNSUerGQ8zC7hwrCTM7ZWakZIDToFuodk2kBynGhEJN5ZkAxNXFouJMP0egOepT6
U14PJfMDhrGTfFTWgJVgY0b5oSdK9OdvJRZcHTLvOo+wohYbxm59CUHQNQwo9+wJb6qW09zvW3Rp
K5dYSID+IsSOdh20YC7a+vQI393zcJ0/XWnJp3KIcchYtiWTdUIgMNtO9F8Ci2wlgkA7JHVSGiPg
Na1zsUhrxhqHqhGP+mj0z4veb0oiXkw6Dus0sJhkjDHF1RxPenOXoiYLcZyxQUjZWACLhMeOqRX5
n9HeCbnoWYnS/EekkebCaNJ2UsDJX6nUX2ZCObpPY0jf2/IQPwjG4jImkSmBGqbn5uGXV8Qjak92
bzMJyrksOQaA7L/AQuhDMh9cJvWSQIHNAFzqvSWRuXExDhC5gGYojEtqMglXNVY8/ni7wD9HQtC9
BB0gCC2hWbt+S5cV82G60tiOW8WWcmVmAcJaf0Oxk1daS5+PE2FWlittdsyk23Y+Lw+5zFoxoKJq
jZjVGggtGJN7SVMAqdW7L5af10zOFfbukND9u0ym7NNgQi3mk+UWv55DDOPY8Y4lteWS1P5ldOBm
Cqd2lSHwW9cer0gLyGlSnS7ru04ZI2tuqbhAG3Nm/sj2iwQ4dW/ZNxsWWtJDABPGF7WrpNfBKFEc
rs09670AbamPnSKYUD/TsuiS6ypEBXxQ0mxupOCeRhKbnEiFJgFrW1MWx+69sQXbpO0aGrby3xbf
/k165nZIsz1tLSDyCQ4pFCtn5nxb6wfwbtaHtbHGmjg9qq9+O25MKzb38vvkYoePLJIsGv30iGgq
jyCURDGxYZDVFYDUFDb/9q+MYMIKzOG/+npmLF3Xw0ePA30n8lxufHpZIBHNMPxbFb5FHpQ247Zx
uu0i/WVYdNhZRB2JBoL2I065+VmRZ4iD9qgcJdrJM/XNd1ce6uqoVBJ273JOA8Vfh0IpLQc3VNYg
Z3PrY/lMbWlRvFUuiQ9cXwDacQtnfby18rVyDRB+i+cG3PfGQu2dXbJJ8dDdqsGspq5Zwo+7w6m2
wlixAhTCPliqEt0raSuGuXNrdq+ot9OVErP8SDAnqhaEHi7H99FYfEwOjYYB9S306rzi7J6Jpz2P
sQGbV8nfixvZN4XEOoaQxNeDz0/Ia57L5uM4ywwvBjByiPnyZ7l6wDuaKb4IkjIrjnULuhj7KJ+f
MOSIu4yIe1CPBFAJ6Pnv20egafxwrLmpXlHe0MpEbmIaB1A7B2kell9bp7lDpLDMn8yvqlmT+qyv
PN8XEX6e82/Jv5VzYzQwB2ZJXJuasozbk1L5Q+FrvW4jnPPBxH1pxgbGl7/YBmSwoBr4p+LjSBHV
RGj1fN+x1LMkiAta4JvsrAvTFwzZwiV7I0QVX1AL7oRCpvbPVrYg4Y4MBDRx0/2oPBMNd8p7HicZ
mO+lwVBHCIdsPGZO6X2NJdVQstzHgFqZdTQ0RZGof5fp86o+hsyqau4qwrxMimuruSM8G9n1fT58
IZ/q0Wf0HJFzfVyGcOaQ/JBzetczJEtnMEKAQWw0jyRksSyVGRBb9p8m/atXuXKrAoOATX5nSTpj
Y61INZutfM60X9pvCUxS4TEOr/WwqkZ5WANaJ6e3JPgch3Cv23DDa0Nbm7ZudBFfwLjzivn141G9
46QxxSRjwy2skupg7jQACfDtA7dcD2CydYScTx5+l2vYA85E1rZNjC516eLPkBQxHY4O5Ss+gBc/
lIIbHvWVF7iVcTNgIr8gekBzt8uI37aZ1a2UsD4dztPlR5pHeaNy8F1sW2ERFL3aanZ99wJRrMHx
yhxZc9LRwAS/WlRAJJheFQpLEMJBowOLdc91HvqeJrQ1GWXufbN7hg2Yo8kCwrMWE1yJaBOt8Ewr
kMSepa+MSh8t6rV2v4L/ERkZ+3Qs9+D502nAXMWdGN4+/G4jN4P7fEJ880JF2lgTgD0L2MmhANwY
oo+1dCtb6GadDdlqOvIYZybJrDyTBJQrt6eA9E5CSjrZhUNSwjpOtXNpa0dd9PyutSxS7PtKZ3bz
TjnT1x2yjYrRJsbTVIrncL++ycnwgUxgnNDHk2S849diJlBZpR1Duu0HezMq17Sj7gVGygagccVL
HrLifnlX1P/8+iGwTIEBRlGIkD5xM/nouxFXsLmsMj75e6MXZdILsmK5lhkydNoODzaVabKvMSQM
u1aDG3sut/1it6lZIHey8L0VUu2p3tGjMJ7NcIhL/q4dc6Dtwmr2GeufJgmxA7AaQiU1bnWaXSh0
kV1XxJMjhYdYNB5Mp3lLPj1PX0GKHo1h2AmTAMxlhQYVP7Jrc/AwMVWkE3q3CTDKccDZKw5FkPmX
eqYhLAvmYfFGFoOo2WYdvdJHw58v32cdwbqc8JFbCbVlSlroaVjKRkCBsBVAHN7iPMUvb6qebt6W
5asOktEs2rh4nv+2SwO3eZABpRZOHVxpWlBKk26y8ILoZSjjIsaz0CXV/44y/E/kG9vktVrxf1dN
nPdsQ1lcUqiaFqLnsAhL4aH06AsEJ/j9vCDWWpnx+RD+rr7HVB28r0lzoMZEaMMvh5JBp4DkSMZs
k0h+OkoFoahRBGmE0zY/XO4U3JCwAeod3OAZTb1K4xEQgvoVzdvOZgsAGFdTggwayH81tpqfZraV
9bBYChaDPMFHBTAiW7IcHrUoRVmBhz/WQSkSJOvYacBD89OSb8xf5OzsW9SoLi7lZoloIhMK/v86
WAQDiWJg5vURLVJw7Xm65yL3lXWMOpk3HeA/T6XxJJsMJmSU5JJYNUAWMR+61pn/LB5T6nvcJd+p
M6LxNgS7iIQBAi7HHkehV6EJsRhdaTFDcWutMtRTl3F3fM4rbaSMAQkILrDaZziKx6b4w8pXKzdh
ljwSGxLO3MhViLqzVVX68PcoxDqqIRphGp1O3B7DP+PqlMTt8WFOwApQMF+tk4oZWORhlpByxt13
Y88P8cQOBL5Gfm1eMzYlvsgBJADthc8meQbpLFFkW/BH6IlUmDeXzshes3+U6b0ru5qYCAjvrP4Y
Esqxg+1PFwH4bAlKxWU1hSOzOsRLS/uhZu+zqGWztp/Xv7fa93a4tXcdXYB4wabPHBSWea9drs/F
tdCTLK83EC9uUqNs6/YGPzNYMk4KX7Pp/vKgRTVP9xCS/cWimEGABu2xsbDIBqwA1SSUrFNmlu9E
0zsV2lT5U0jA8HH8c5L7YBhgqODi1vqs8CM2xPEgk2hw1nOz6VVgYLXuRV0tyC/BFZsTzI4RUVXq
dKMlh9EZAemtAamlA8DqQzsh1TSnmUJ2LJl820PYYOT8zYsWG3RDTIYdHmBwJrnZuT7lAI0SO/JB
IpG5LUa68CoCJ3pCerhO5feRpUEaVhL6vo49rf/++PCP3Aw+cQ5lO+28Prc4cSweQjZ+y+3I/qqN
5y6SFcQTiQB0/AoTYiHE1hOWmlDA0dAZDVds/dkQi02SZ1JVRDUkmiq4Uqwqh2MHkMFFApZmmf8P
xVhQlZuidbofUeuHw/DdJ+eXL4z8KaG12kYlJqJup+HatX054tAj+YeXxUBhbfhZYIc68wKiijrE
/gnVH5TcAefJWKyBNUKkve8t0Ah56COnJjgnh/w88P1bvkWwznTFcavEMAcBx3DszocrXm6Mlp/t
a+IS3t0qne0yGigraVSE5094wt7RhSeIii1DMNAKKJ8TjDKkshBDMR87LSy5XDbCc2rTe2s9S3KR
u6laxCggH1tGJkuD5VRLLQKIaJOYRVUPAGf1+kRqLdT5s2gXy9Hu9Ol/zRYov36PIsZ72Pp8XO1W
shiD73s7JIueV459wt5qsWPz1wryEolvZY3Ij44Isu9GJj3mBM4E1pYlfitZv6NXMJuXE8bG/pWG
oMjisSaDDSMw7v57+840PELoFjFO61CF0rmASvlpmATgWVB+Jl+7+P5X7/FCNXfErBLIHLQ28vBE
xWJ1CsINxrl/Uo1DcietlI7Qxdm7LA1o19DFHlOuINJLmWYvjg7jDDWs6Lga23lf2z6tY6T4hlF6
IF+lY5dQ5xu0tbbcFpHV0jza8LGd5d5HBJZAO6GwFPk6K+IsrNs87f+2TA05HixeOJNtf4nIffEN
uJTS6N9nnVzlaN2cK1Ia1MwCQEQkEJ8webtfouWhkNw95Qff9iW9jQg5cSTUCzHvGgJIpU2wfosB
doPMD/9d3jnjqRPb4lzNIoEiFFU5kmfQhNa76FNmCbkM5mvsS12kDJ1nkVt10C6M99c8rVDNyobw
ikWqW9pedwaZaibqSxZl9ISPWhSsny+Gqs7zLejppSkHW9UbNHRec0k7qV7ywc2n2PDGZgzCjc+5
+9Sj1n3C08vun71ILa7kB0Kmn6b/RHYOhl9KqDGhZiayO9a5WA1FYQkEi6fsTZzEfiC+za9A4dSA
md3aAsADgkpLuQuj3rPhjORF44eI6bqmQkRtkjYjKLy1h9gTTDHfec7geAQPXqBsKlNpibwA3H4Q
Pib6xgx584/tsqfOn5/hD3e6QNdFMR0fe24FdRu4MYzb+RAc1b0mMqyb8naIwpyotqosy9KJWr5f
zRxqqbwzrYKTBoyQFROX433G4GFbAgTiX361G+5hTzRRUdyUsmxsSTwz7V9afmdDt3015GePtXRt
bVsuT+w6tiOgLJ9rgxvUFic2B21FGgCxNjDFWIdd8/dcP3S5Wtdn4WRe1ITHv6Z6XtaMAxxynWrL
EMeQA3ZM+iu64YUDc8koGGsH4LDspBFqGeGkmg1J4KSMAIj++wCrD8RIzvKLyTcz2hAi8oXjz2MI
8dYLa5vneuJeQ2TsI9efOaUTkOODjGkYtVD4ZBIpvFUvwdMnluaFrVIqyr4qcQawg7yNg4+2fB36
ia8qCOj+HrONvAJqCe8DZ6/FTaTNxypI5ptDnKeQTnMzIEMRfNq9JuGJvi78iJInWQp23A3TZ19j
3r3B7m4qoOGE+g1jZ21wCVaV5vgXSw/DsalBOj+98H/YAE5AllHeegAb+B/qd43JdrxkRbnokqBK
16nT5+J8Rooj7WWDfVUaJyFICbRhY7WwTsWaHkNOradhETazdjUxrkEaIwtuSLtM9BY9CNmWYZFj
m0eof8Oe0oOtCRqTxpXPdVI3iKmO6o8os6AjHXEN6L3yLSSmT879pqT/A/OmXXz1kNYtVMv2Dn/z
J3ODy18q1976O1ypykb0/k3PpxbM7ZGqicNieAvn+cAcu85WeJfCnWumEruqwDyk3jbfdXnY3L3/
z6wmbyIpLBxP978/5qrEAFnDgxk+MYJdzz7ncPF2Rs3XiA/FLpvs0nrWiAG9hDr2HfvwfHK9ERwG
zw2oxJJq7FFS875lpnX+mlcLTwME/bko6WNgXuaRMZtVglBZDXYdHhv0Jzyh4jMjptny7vXUclpU
V5CUQ50sIHW+qaguGTUSPgW3mZ9CRWS7C9CvtwrQC1uGRhwQbCEiJ91RskMeQJrgqHGASLzrQV9p
dicD4QxdIXmT2FUViDxxuVEHLcdkUEYRdXqPFKYRHus/MMPhbOwP4zjU/vs8bSI6lZHEeYVuionh
Fa2/B45Gpenmq7jFpVzILYnunL55Fl1SYRjG7SkYEQS3pyCziQGNCd2bi6aW2HC6fzkwqQbNqEZb
uQ/NP3Z9BuA33H8uwpoktQ4BsRi5/RDXETqLPRRT5KIAGafSrpOJFCoYw8zFXxRRPnhLaImaMH+U
Klsj22C/yft9Z/alSmArhEQ5aEbwRZaR+OG7MMxTWzn4P2DuG5/kSNZSwhY60A2XUf+FAxeq8odu
bNeKyOFAbZPCH0EvI0hEQpz3FRtokzKJC4w9EHSAjaAlGxDsxeRTK9ys0cUm16NjfnUoT7MIsUu/
hLQln/b/F55WiUZ+UD4So+gDF8h/L/vv5v1UiXIVS4ZIgfcI8UpfyvZXj1BuOe1+Oe2/MufFHdjP
scMxeLEs0PzrULE8iL3AZVBYPosilfs5xH/7JSuEVX50QLoFLcfF14HYCLI8y6iDAd9IQ6xMemSY
doMLuAVGiVYgcuTYYRhj0KVFeW7q7ckLG2xSM5k+I985TRQZJ5pPyEHdowwCpnlNRaI+nhGZYLja
CyA0STXDv0Q/ErRfuEU+/mAMQNUXmCRW0KeqhGOEdf1h9GB/6Ysajj5WqjJlkoRZwrtcN0R+vLTr
f+gXZaDmFOrZ5gC2SPqYwooFfzkE8HWKH1fNincVeKClBHFTdy64r+SNFRG3vI/FihdaeKxEhkP0
KzKsmvxwo0eVra90EO8H0/JPQcbjBQU+YH+7mG/XVJmh+e4ggB07pEEjTRF47ghb7H3A5ldYKrKK
D7866kWJgk2gwG8EpZsHrSFHI7QJTZaWnNbv/dPOucATM3bzaVMktiPMprIFljmOyW4IkiqJ00LX
/QEcLitXNRP96ataD3uX8PzOAdR8LH4bbe3EtwCT5/4LFUhjQS/QI0Rx+Vw5+xwS7mg+k6vviuKC
+W/+CTEzkPTdPLuA5stWDw/kmTaQnc6gQclsC4eMj3q+gXS6VIAtkl3f3Vgy1GvVajXnwMPm5uri
3cDrJgdcmjWCfyLKvxU817LXEntRdd5dlln34V4J6zjBGBFLIgy4hOdGtw+TEzWwGTIrVX7Ytm9r
uM5f6NTMbuYheM8EOWFCuV7idIjrDJiB9IfgeyEzzcWtEP3GTIpW4yEz3EVaYdQPQCQ5bEEQxz+F
kXDw1ebpKMLVFKIsYUE/VOOEy+LCPLDwuWWRnD8r1XLr7KdelsMuLgwSzQUVHlmBibufMNuOfaBe
wZTjRij1LJ/Zw94ImmCoqkQjchUgdsL0VJXzMAs/yHLMrsNFdzHkDp/Ugna5+MW7IOFCBShQyNB/
/5gFyCiNjKhGVI8PjqZnMw1WBldZlD1HyqTCo+eB6aDNpN0j+Mz8dBIFlWaBQMQHQV5vXNiQz+uY
IJ031bhIecWIW2tQvWJY9NrjbM0T1l5jvaPtASg8DULPH7yu284HvHhqNHQJ/2T2e/5SbkzR5NnZ
id54Ya8TpiB67drFMVwsu5q3o5y6XOjVI8OxsUWV8kgV66sYZ4a3rF7fp2HkX7wa98Mzpf+RJ9mp
iwhiL3kHqz4By7lQNQ4rdlUwGF3aFytEJRxHgMOr6RthtAD/L7WtQnfxeHQx84UKvp+OIfLcVAm3
rpjvGrGvrudrXskK2cgsnTBQNaatbT1QCmXb8/oKtezNgrMn9Bh3q7nQfcBwkBneAQhVFe4X1ASF
SE0e1D9PS6SAXJNHes7k2/XHqjysrbGvw6/HfSSyC7zIOPxfPr8eiylCEkjdt/Ebc18Hp5JAU/RH
nzgh06WG3v+7mAAru4ctcqHT2TcE3Jga+uHMkqNGwjLrHtVOwqZ457CkY+xxz5Dn/6Y4Xy1vGQxq
J358zEL733Xl6F8/hxJj+0hoPGrgkBmYoWqmGh9qEl+rtlbmyzWj6Ylf/UwBGtcnHbILWAZdmIVk
lJ1VebqsMyRCdgCsze2fzOlpolpxMEPIwT0J82tpgxt7xwRNI8j794O3wffw3lGGdKbc8C9QlXQo
kL+fDNqcOg53l3LOz2zf2zlnSPj2Mxsoc4WLUwMfyAGgxIszk3akl0O/o4WjJzDY3blBYQH0f/Vb
9xLRlDWqBoKcmZjn7byivWMl/U3WrktFLO9Ap05AVdalSwjJpP+v2fv47oWQ2HMjN9X2lQt3fumM
QN535QpZXlS9PmWgmAGzCglQyrzq5ON4ceeE0pwGy8cms0XP+TEQmS1I11EK/0VIaheLlqyLH8Wy
NBKGUak0vmeXvNIBznDo/UlSusMH1CDb4DwPPsg7kpA27P8iN54RGpKN0SqN6lT6Nv2YPKZpokXX
EdHqTORn5RkueFb8J+9pXqV+1+gO5KSk6nZF1xqXPW9tYpJoEWoqL7RIXjY5Uxsazlf+Sa0Hgt2S
qmtyF+381+5/2uaEVZBObWtYG7bFyxCG5XzHZzlTaU9MKgjT21oklMrb43CbFpq7AGUhnrUuOeLU
entOCbr/zfZu2W+QgRIIStX3BWiC4YWpJ03oqYBnqPDH7w1OXN9/xD717i2Z9ApOezXlp8P1tmAD
8fz51wNweaITUgQSXVZdJhP/1VJTo/oC24AVqH0i7R/9RNzlnfhujmBNvW0Gxy0DehRzoUceTbCW
LevF9vOF8Xr3wSK3vxtDc0vYqkswPNFQelKqtZIgq6p+KBFAptXrLfisMn8ZA8cGRVvwh3hgqBZd
H0Y2HDiT//fHNk+u2s+wNCBBC97ozQhrz9V1qj+qhajvflDDBFdbhkRPwKoRKpDNwT9+j0fzCXXe
3gjC6S/N25fQ2VP6IOYJbGLh/3degNaNB4rTDPw=
`protect end_protected

