

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VscJIfFTgZka3rw2Lfnx57r9iSPhRXi+kLnhdqz5EO/+OA8vdexQe6ce3UDnXG83BVOJdHtdZSuI
J91AsMTFXw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
db4dwZATkWURbjXQf/P3qPhf34lj53qLVmViVUVBS8BVdVAAny6oLUuA0/ARxZIkZFDW0nLTNAc3
iMNZJbDRMUgL42wDDdFSS0oTCLPLIfIjVZjD3q8kOVtOgpkQjAtZzHWdc+/y+cVnHMQ0BdzqR4XC
mD1cyMlG77UuQU4p+Lo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f07j+8ElH+sVCaM3Yoi7ry8dCLtvbd2nmyrK4ZSbRDrYOFSxnjql3oJk8G/IFhz96acf1qM/kinM
4DSg24V6d4iNF+Sc/WwnHHVdA/DQDGXwEsGvAxVjgEArzO/9ovaPy9zXCrxiRBslsn5sx3ofkmXP
r8Do1oTxPaq85CvX9w2/5w8r1SinpqLeUxXnosg1l6oQKNXnEDWv6S8+OzWcSZux0rh4et3+Qd4Q
vnNK6SIGpmlpWDDbUsOYL8An1ef7zNTEDVIWdCsTfYsl9bwkYAxxQ2Lkg2kESygxpths5CuDLxLM
M3annWfhnSarZkHVFU6wgl+uF97yURJ4ivAvqA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yGIEomvbV/vYOvjOV8UL/R6cepGB517KBp/ApWDS87JjbJ4Juk0Ygt1vk+okvNIg0yHv/44OpvyM
jmFTaFeB5R6Z32brqQgO3j0BP/DXa9ZjjU61Ec6EVTnuHwKX4Xr9osaMCcSMGmmr9jzFTwmx7CAX
5vZms49D9iKwWbO99kc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nB2fsdHzYNwhsF77awSz4nNul22cayQFlU46LO4sKhhVNnJQwNrg4Ji65F47QLz9crBwdwtrstYg
gMKq/9Eb+5eQ0D16BOx7Xzszn1GT3N/ZqAoaolBOvlKzK07++on+MIU18pqvHo1rjvKUGgimiIM5
0fUCAiml3CQQ3SVWdl5y+ovbhpdhjzmjD7YPlpSVFot7mVPcO7I2aCOSWVHir70XuPbF20cHRAZl
gLtBKStSr4oHAHAYT1h9naJsA7G2ZuRQO+G+72/Hn/od4gVX5tKZKLbga8w3D+ucChWWTLI/VAMc
0MRZyQD+9aE0bQkI7JDrGrtpCtyvAQffBkemcg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8336)
`protect data_block
rNLPaZ7yhzviBddUjvU/KkjzDdXTZQ5Nx+Pfsi+tFC6u2K0p19ivC75xBsByny0CL9ZbDEF0iB24
x+tgC8R0N7DA2j7+FD4Mn6nRKJ89t3PPyOIsFlO+zUbUfTOBtRB9zaoJ50xbX9LoAadIRLubt7mK
4+U0TvKWhaudgGbEmS7ZvS2HFveVSK3YMGIWc1mgp1xPAFcfECoKvey82S8/1s6ZfLMFZQdhsiSK
cX4xy3IVvcLqBKM9gBPBGXV7lix9RFRoqn2vvENEwk70RXQVov69jnxBNU3Gs2Ii33oXG06xfmsN
G1WrOaWifA1zeQJXWIso22FKSDD9hDxN8dn1MrkOEv78kZ0/WsKBF4s38Q3hZ8r1Vnd3QdRVLIW1
8Mu58UAIrsTgIJrDsRq/hfyubr9sAIZaE/Vbhc1AK6d9XWUu6Hr+Iu6QbiTlPC0KS1h0b3VaLs4s
8FxI7buX+7hYVouIlPOSx+zrh6Is/0vKLHgJ0JypG41oP73haRQyuxvRM60ZWPNaXQ5gPjoAfbLD
QKUHgYpitBJVBAZalGOztlgGGAxibMZXokZKxJrxlT49u2/AqANGDP7vlduuED9iwV8oyYf9mUY7
1xoaIELqCuI2b3BfxmDHW5zuClRN0VSAoHiHvmWB5jFOHAWQ3qagOTUF547Ri3K70wkWDLIJW9TL
OPQSQau5W84l9wRKMLgeh6n8X6iQCYNkdriBzDs3/fv1lqsE4aiEDMSkQW0ePzvpULJbpxdYwx/W
EaV9F5yIK7RoZB9tsgRU2RgltW21FjkM4mXzja5pm6yNy4Q/r2RYHHj5fz1DLDwSjSH9coiCzXve
JHRHoF38R3PiO/0mfld7i+SfmTLNr/KHy2kOd86C4HxTOnXAutV45QTNmpDDvS0eQPkdxdnr+Cjx
Q6FpuvlwLzQltzuUqgzHZypkbbEdwLQrsogO0Xb/H/zp0rBCoSFBKIyouqAag6Ne+pv7UCQRvUjd
RmJVIa1H8MqvwA5v2jbV0rrYgF7vqntnLAG/IS0W2VEeik+MXghHPk5u+fWSPMFrXEBvKcjMLzBK
43TdaXM4wgmvQJQlkQdVDyhQWb+MQcmS7zP6AgNwU4P2BOOoEmJQggLT5Qb1J6tu4Ei72+3YJDaZ
ccUDk7UtVOJynB2fBXwohmaY4+9FoHf2V18XvP7nOkGSCt5c+4yrfEYX6NizkPXugSPycrzklv6B
pvyeHZPZDtbjX/0ouf39BsDlEcdoaXvFySuCaMOofc9k/ZBqB8amm8GkzSds9J3/5hkmOCNKmViH
5wBxwajcKV+/7jkxMf8+3I5s9GvIZqULGGCMjidLRkSMNrT6ivwJC8T+bSCNjkN6K7CZuOgJtkW8
VADUypqXTgpzejP4f/WqsJOb2hpEg4ej0RJ6zzG6th8io6kN3O9KvDMZV7ey54TI584JW3TIVP+G
WI4bArE7ehC9BPemRYp8iSK7XpcYCIw01RTl6jLX8YcNxSoyLyRA8ydmxqZmVocnS7/2uyVxEgHQ
B9ppA6SLlSBK+0vMG+a1HtEnGSZ/hTCgUjJIhyABT2By46HJj9Ol2Hgp0TbmMc4WRBH0NAkgLLKt
q17keR3RL9+NXF8pqFNYEMrVh8VuHcdRAxF1+VsfNa0vCOHehulQhrEHH6bgPX6Xj9xBOhnKxmxe
McUHbxxlm7ycO0oUuGcmdwj/PzCEFeQ78OGsIbDzVkywIX/iPDorpJvTyPrgHiBiiLfs7BsuLvJK
ZxawFqNY/A5KLOF2/NFqRKbu5tCsNoGRGHryi1R9TvPX6uDFXvC5CbGVtBS9O2IboKP5yolbsLkU
Xc5P1zgle0mOHvXGn1Q9L73tCdPAVzOQghjQsrOWdsrfYM8mpWrkWNFatTYfE2PM3oB30restTIx
x0ajfxQ87E+b7erQg00ZaGirw0Ja+ZwGxtfoNeTTc+phijUIGjPVlqvs0TsF3FjqhvHv+1BxcQJy
p/D45hkXLnOk+5mMVZWemN+lBO08uXMSw70z3V3Sib1aELq+Wt2kLnkrigqOVBpAMrfMJXuJd+Xb
100PoFOhZojx3oCR4W72RAmjg/7pMDiUSIP4X9/bJtcjhAZlMHIggSsZ4ZYIZHNgi8U6JpKpdjLD
kTNkAP1+axSltdmvHri77Qz5zSaUyDiZnQ4iQeyygfMcx7DN45fXImto4Rrtjgg8qy84Scms5SkX
XhLVwTR0CPbXMTseICEV3S/7RKnfil3O2zR7MWpmyMJeJKJOKAJ3/RngF13musZ5c3vmFEdCOeXA
UXdOgVw1X8l/ueIscgMFTTiI+e7igGl4jtdcmO98uqHx3k9zTD/58vJXxCCkY42sbUsqDUOiIpOy
QP2XrO5za4CIxLfF4E1/IxiG0vaGFt70/w1FAwokXIWV0rROhGmyAXxDpAH/6K+a9+gq2ijh0LUt
JIRMWR2rtdnz35rhsJlqvacJEDyoAjVWZ1c52JNLOLv5Qscx3uATYPJalaMNDPxyb4+Lv/ujTpl5
uelBtGP7YI0pMWL79KDN78CN0a4329slBm0rqRvFbBWRWhnCJUz4vHKmBKr2P//siEO1nU78TBfk
fXTX48jEpRDvdH2edVZ33dx7h5CvoZfVQtcoxxBQhh/qUnFgZ0yPqD4N44+09ZsKPU53yPBILLB4
EWS0ih2qD8WRJNeTfTV5qzQo6NQX3Ai9uwdkxCaNNkE+kNBqwl7O9wfsxnrZWIFvaM30u5yZjTWZ
UIuXOSwB2p/jVZv8w626pzpdGyHUgK248KjCh293Cmx47oKMwWtrqsNZKS1rxmgs1FoNVzIE43uF
2YWYWZ+s/agMyeZwQS67OVoLETXHunWdqZUnVIuN6+v55M95krkGHVIJH0MB2xfUljI09k/V3scx
lWw7+foKgZoVK4KDGmeTlvSn92nkoCSEF45dkCHByCIC05IWGXibSBEGZYjg9VDvB9lJXpxckMk0
I/xDK041+ik0YOIhqr92k0zUY+fFLIzyvq7gBWorv948nXdJfoJpBLHEfOTOxkz+INt3xDhqDs1j
FBlMkb6Iso1x2wpwh6+ju05jmPMRzRqRVhKwX/JMz1Skj3tavO53cqoe/WgvobaufnClVEUcZ1mf
RdSt4HUt0vmEkUUknCNWwayMHNYqb3Z1eGG+fckLTE4ASk8ZGLxBEeg+3itl0qZvvADUYaCZrd6j
YHjI8tLyu/apUNSn0CJglYvklZUDVjJl+Ub+jRGR09+eT1KRevE2CyQjAEbP6TLe1SG0NqUYMet5
c8AtTCmVkwoLiY7OlOVB5fU3hFX0+ydsqxPR8ibAYmVKwng25Vu4p6O5m6EBicnvy5sE+M9qaNFP
2IDAoqdWXjFLoatWjioafxd60UGVmvHb6qJQ4BQhkZMLI0LE4E6MAmSauIgOXAv4PPTS1JG3G/Qe
bJcDN2dpZJQOhPeCAoF56M3k8El7QjuaKuIDFULpFFE+fO5ZVJ8rEnPArXBEbS3tTVhD21re7jgi
oO/nf9EPHgQm9cToRrjGoTYTxa5PqyvOzoPjBJ6g83VaVARyqOb8mbnhVhoN73vpkMN/z5hkxhNj
69/zNc4IGPx1PVDHOaalVVJCdBzHAgbKboaygd8utPdTuXv/n2YBMumohdc4ty2ysvDW+P33hl8y
Qu/RpwOj/aizMWmR6EEVHclIin1/+Pi/uorsc1u8sUd1CsZuGg5jET4F+RIjfaYrZfORJKHnNS0w
V029NN2Tef4Gl1ES1XYe5+U1J+Wz7VbwWBbYL8othvQnz2yMoFHVq3M4htJwH084qL2BvC57/lKs
slRJ3AHqDNuD1S/eFutvB9bBQ59J8P3AVyTkLM2r5GUYAQf9gUPd1qVPG+hqeSx7XhagbBC9LO67
g6ZkiRWh5RY+5GwgPIRnIDIzEw8GG38lBnRX6V4+LTRyHyCCWSdNRiGvi0sbKaxGnz5G1OY2gJmp
0hwBSF3XiTeI8gH+dKXZtpnaje4Jt2OdwzWr2j5y+dw7J9SL8zTw2mijMm6bu/tCvgN3jj9wwo03
qToRHskni+Hxu4IcEPXlEbLDt9AU8u9sSVAcs8k+MAxLFq+hciIYC/ZmQPWLJ0fMqkob4fBL78Lk
JQUCT9L70a3bg7FuFYznXJ5zVdZj0Xd7FQgap4kXp7MnwTg5J5J4khUJvzCCEI3TJmA6+OKBICvz
CKejAoLwmld6VNkYtrkmt40QX3nb8ZY/RlTt9jpVAV3TpnaIKY84FQzU9FtEuIbFdHFIlUWb0Ow8
ImHwRyVHY8d98+1evwiv3kfyKiwc0CRNGoh/uIRi0DPaSpLdiapSiaE1cD90X6cLE2SFQCuT2H2M
6Kux1eOc2hqy4UIKoBvMRX1q7/xGi48H9Xy0wDqY3ATRBPIv6b8eUYc3h7En+dWDf7wspcWlYlw8
a9svIYGgUe7gsXTNzJPPwJBnjEfWIoUMrOfX4/W9GryV5qwzyRr7TKZpkYfEyU8ZdAuUa5CrswyR
drirJgtWBQ4378YgoC0UY2/vEUSo07Jlmhue/oYTdwrGmM7Get5cDThGqteUiJxkvQlRo7GXyn3J
yqwriGoGqZrDgMvXVVFvDQgghDPd4o1Q0HYjO9kj0sd9QBRBNAXii24j1NMP52YkQqVTOw2YVEHU
V2pt3AvT13rarjLgQReYFc/RHDoVAvozBb4KukY4okKgunD8CNWmqMWMHjEJ+iAnLj3+5O2iRQiP
9fr+cVZ6QlLGu4/FCJSn3aq5SaLL/hKAujhqnH9nIdmdykoYsC+sTQYyHG28+MBNbscNjmmrp+6H
g0lb9lOER7Kl3HwiCWM/HZKAK/yvVFiI1/+WlboACmk4G8qdcT+ioOK9ztbTpDdnfmvgcUn2xig8
su7pA4sBqIC9307JK77b1GxGmNu6dD2LqaitYPOmC5FJ6Mgrtbmsv9DeoCDiAxCRTaXLPN9gqZ0d
l0JZ2kzuVRtMCEm28VyDBvJQsf92125fCVsbiey5rQOUHuYAdrE8uCiyaZjt1aLrOX200cC/8KIV
XHSgwItSfplpr10G9r1ZQuvuo1f+b2ZZUUpLwKI6CrU5/cxcO8bhOkDnSwGhkwuiRONZCmDzDLeg
JOMmvwlRZcBoofi4V4iGaGaoBRPFXrQIARP6NfjgvAldYXup/CdLDGiU8curdN6rRv9OCQ/qEYve
5YHcyNZjZWVXiBgJrPej1XkICFVesU0iLQu6Z/5hS9D2hbft7v75rF9YldAY9A4FNyf5NAIM89mO
wkgug8BNsiuBFd7X5BOpk0R3nH6pxoSISjHBq+7b+ReA3oGjzzuLNaXB94y2r9oI8cdvKoCfW+bb
hsX2K66JKVWZTwLXxFkugc6wzrFC5f6ZB2/PqyycHn9BozsfqJPvyqQczeChJQjHGHAfvO+5+X7K
IC/XXHpqDahttIrs+S8cofzWg5NnlVv8jvIXZJmJSIMRxMOfF1CuTboqoI6p6xBtEicqUal7k/Lq
Ek/B7B5QP3WdsFc+eqhuFdAxskJTPO+lb24GW8LYb3VcykLEdzRhC0ftkPHbO2+1vN2CzMbPn11/
Zz/LgCyYY7fV9i2LH55rI30FfCpFx8/MzuaaL5bav7VoB2ZyjWkPN4ML9Zc6GWSUsBTbJZ4PHkMO
6OPb+9CsNUtQNMO/EyAICbwAa+HsJJhJYyd1Q3Pkcw7uDpzq6A0np7CZn5xN6d3ziGMufv7nz9QD
7p6D6no6K70rUp7N1Z4Svg1eQQv0ljWbtPL5HnnXlgybvCYTbJzyshC5VlkpKKSamF6ZN+yEf6Un
heZiMuu6nYp+3kElymwtEaNwVWR5HG4CBG+QYTSOjFNUQVJokNv+DkAPMSdp/SxoUrj6QlnU6QoB
N+cpVkn9Pn7qcZDrkimiLOKxbUjW7GyL4LpMvCestXr6Yc0hxzJDYkzSuutngrewafUEPON7j1xl
89wETW1CwA9zLhiRKeeKbAIS5tFBFc6nIE2LSRepeAM2kCUVi6UwfuqVhsvZgYUHftvJiFX1wQih
yaGdiQAERY9VNt/69xbe3bBlivjWn1WvCIvHIpJePB48vpopzjBuo3sCAxgTIWWYlRzQXC09rlSp
grGRGe7IGvtR4zvleNpFpKL24IFou1ZtYo1T7qvmrUc1l3xQHzxi1AdWhTfBTtStLiqanZ3gWE80
tarD7rAeCgefHf4V/WagY3TmMCMzMYfB12IjjBxYvi56QRrkHWdNcWhtLdYISx7VIAO7Rvwo6aSd
bXZ5XegRGn4TicspLvwItTMz30zh7ASy+Hd+G+TlyxmQY3dqIs9SfExJXWnIwRMmmjJlprxkm8RP
65er8UnX1jfOxwOm277qY/eidjRznMdwhgyTcG67l7ssN29HJ1pqDBSWjdv5MpJ110L6uXiDYTYX
1+f5bQEYdQ43KuYeCb7ZRMFxm8kmx6TXEC5qrd4CM++dbZjEDRE/nHbRcSNVW+dxGIkzPYTk34Nh
cBeIYmy4qsfRhBIDsc0qVrbbxL1H05OyS5fqLIVCCdI5mMzDGHGyhDaiObABMARgNGvKRa9mKpvS
SSmO1Bemr85CnQBXA1jGsyMj5+YmQLPNuJT8UTuAtfjspA6Ta/9N0yf5nVUZXFdN4vEqUIfgUEwX
TVcTvgjqKhRzOYRNkOipzRdhcWYOL0B4qlHrsl+vCdk5xyyncWtDrcLdycg1/r+5UeiSZwWAr9bP
qs2UYcp4aW+juG5f/JsB0W7rZxCoWR7cA6sit3VuoeLA35TIUCuwQLUdvfrVNwAJEdYWTaq/zWbK
SiUs4iUa5cdyEs2h+KxiT+LoO7X+Lni3TH72PeCcMlnHbaqOuTEQrtri1rTJyA2oKeXopwHxFaiR
dgvzDnFUCPJdXsP/8zsvudcChbUCmO/G0rNOT6P7EI/29MfcLGwtiHFnCkH/iFbaenrYGXNnowqU
QizFxc0SktxlZn0sGW1CrTLXr9WzryO2sL1ECTbjl9pKx09e7+CpLYQ9fohaMPfuZgNr2RqOvKQj
0eiVt/oBHTBFEd530avGKmQtvo4snL2J7Uz55mbBSBDfN18u7nR2fWDgHJGX6Uojc4iRO/OTvJPi
+mLq4LNq4vkvtKUMXf362kpJZZt9NYmS9ZhJ9xOyP5GInLglYLWqa/YIlg9mGdPZPY4d/ONCN/1G
lNLARw5oPX++5gXBrwzp+txsRK6+xui230+HonGVGTNaGd3zOpRxdemEsiOMujAsbYT5uedFYA3q
ar9sEp+RU3pHVttsog0u/vxQ1oSKmZuod3STgbsTy8UnSIQ+IoYHMTG+/Qy4jPDKEMMhRmNM/3/t
U4NVlEyn1OBhWYbb5QuZSDh3OPAY+AA/CHfRFB0DevHtXnr4lFDzQqCe33m4DacKJ6TaM3NjOcN6
HBbv2Hv13c5NK9uQ6stifNk5CFxZKNA5OUOgO9EUIcaUaC3hOVKjAFLmwJ56YnsfXPXddDo7Shpq
EjN4fPxTwSPL8RlVlFtvHYqine0WnqFEPl4/+RxbZLL6enB+Z97GywqqsWnmtyRWMNNgmA5x2xuf
N2G4cXOQXakG/+mep7UynHM/6Xs2iDpm5tdk3BtPvozn7jnU7yJgFvhiC2xRJrs8AUmvpEs6JBY+
aCNJWvbqplGQRES8C8xsu3+/UXPr+XOcEEdkvpLXWtrt0uT0G/GCX1PG68fm/cXnnR9gUeR28DTB
p1TrSaqE3XKnq2sW3Bq09MqJtTJiJt0j2fZ8dRuZTWP6Zr0nTgjI9nw3gXNuEk/u9ey97mHcn1bF
ZzaKeVu8Yhxw/aI9YWackb/X1fua/LzhnEt51gdYEmbOrq10mVAGX+UNgpUGmZuSVwbPH3U9koDf
eZ330yE2wkbvQyQAV98XDarg+YHoatHXJrzP3TZexKmW2s+IQr9iEZ4484bPC44msCgYqIB5b/+f
3sKiyAnEEe4p7A9q+Hqkr2Q4CfgRU7M4eV3LK0nwKnlz7ESEVhkkhVBFJkpRgKN7tFi7kLJ59Z6D
Vo8DHq7e/c7kCH/aCXOLJyFLsUQC8mrzuwIZirig0LDR0dbjIXHgupSBV72F8E64qT6lX4ndIdPb
NEcdmlcZgyE+s6NDntAAq0KnuljfhYS/6u4DnWOAxiypTYIZvlSr2ID7xxjP4p2r1mTcIZ6mPpzt
vvDqIY6LrwByitCBtQixVF0ybwKwLFY0zNXg/df2jxnp22JraI77AGgN0HkjCet/I6jOJSrrG28a
YU79ABj/TFEtepeU8MYwg581UaDW13agzbYuI2tpkdl+yIWnEYOvqxm9rn8DEk4OJYDSVFTA4i1B
LiQCBBfXAgivYRE6vt/1F4UMy7SjUtVfVF4/UPcTXrLW11jrnZlI/evPY29XZDYJ7jfjngpaMp59
VnN/jGhkMvIGrAWLiK/acm53I7L4eEDq24u5HShQgXauLNN4KY1jn1g7q5VewKAYeyC9zjiLJWPW
GhR8Cu3HKnoPycKzp9/yt0LdkgCj6SN0vIx3KYwMWULvwzij/aJsU+B7Y9pkhRSXXHhh2lBQwwE/
jcuzq6xbva/weRv/tM9X/Q/vZynhT+LNfMaj6DepKTZ/3IBOBCNZwA3x0sSoST2ZPwrEQS24OjxQ
qDKSRSCq7Jev6afTVRAdKiJF//sFN6r6dvV3wKhAtWVk8C1poyT1+vOLGe4BvL9vTRJxZDFGOG/C
yjEG4q2rDQWa/K0cxt066lWmltXjUuNqTDfVqfQWFd5XtILIJFWgTDr3WzDgbUWjfTWIv2acNkzT
8rn30a5BxvGfuOpJZB7PDPV46zQftUVGdv833snpUS4reW1kueUum5lr3rhiandXd/axhecay/oA
GCLdfj1rGIprHzBJSi0R3ZKsvv+ru15JlzpasDlZzoR3Oz11Qr4ZuOHea5ADtfL7S7dVXCkQwz9V
psLpfvMWakTACu5QgJg//gSA5hc7hP3tjSalF3JInTOykQWO1QQRU4jy+VcI3gTl21tKfbVZ+dzE
Xy1/U2lbcOoqfHeYasfy86t3TU/LNDa2U5NEMrCmZj/IKPQQhK9lLILYbzmyGoqEbW/n1AUNvEh6
A2YepJN4gI9fYJOHxi+0Q4yDe+gG4+vm57nGEMGqGviRDwdgvwrdocKH+plxUs6xsc6XL0djFtC6
l4+r+vPuTwD9dKyonMo0mTMXl6ZOJx2P1JEVpp8BggzXbYZcvFQoDQC13V0LjA+DAuVIrnKusuNa
lD8Qed4ie8c5QXH3S7nxxAppdvjOnHPVZD0x7RfplPnHVlo0s8H/CCvyDir4ungAl6R/ttO4M3e+
iz1doM90sHkOMpBKafPEU4s8Fzazr5n630AKWOtMgtAJhcanOnSc75r//F6pK4/nJBL5jLKu0OIO
Wd5ANxxMm48MLjq2BeH+kn8uUVQM1ocdQZhSCNalj/VIEBL7WSIEdDEyXw3Hs+7A4GiEv6vfq0Dr
OKyxRIk7ZMz96f6tfOqp9Tl6f7BykaqUgbb4FIGJLWO4+ChfauGwxFFRzsA5ltKpQ8L1pzM84m1+
jo/0uFmXGGo0y8IBtGNxjgm5Bu21OkZH2nJkDFvXUtwD7OAWOy1aXDa+Vt0BIlX45lE8/dDRZ5np
51N/WZ0Ywq/HnrgA2fYORiPO+IGSb52SVZQtOW0Fcs7SQIdQqusYQ8Evd8v/ThjJH6kP1iPXJg0U
V5poD3jEJtOec/tAfTNVHMQ7Kep4xZKkWinUWa8gtkRGaQhxwKs79tPXnrSHadytjv+r13eFBmgb
ZpUaJ2DXAvltnfQS6QRbC1risWx0P8nX7PJrFIjWwlpDgWqY2/fxU9r636JFwKjXvxOv5Xu3JeR/
zBcQ2m0mjoBEwqduusfiQbj/dp9wrPITe6apT9zfzveVl4S5RchsR4i+/3QSVRhTGF/TLM1X+i8S
w9bnr4ciaoPPcPoE08NrpYAcpUG7741vcArDILdCzoaJRU9BGJGF6mbqILErFS/IMHE3VEkevmed
jwUO+qUz0mG5FyXKHo+l5kT1b6Ub8RsHc12Ie0N86VuVECiAx+QZdDpUvq1wsbMXKSU/VrNonTef
sA0v45N6v8EbiLUip5qfXAjbY2EayBH9ku9bRzqswscDNwVFCpowFSt2y0JY/8c/D+5e3Ol+pdq9
d2pRRzF7I35wXJC868YFgrJu9DQZSBO1+aecmEobUaa437rGIKWhj9wrydLmfiKdLidg2iZNOlJ1
MEf96OF6kUgAL5crT/YcZ3KO3g5EAQhHqnTUjupuQ1Z68GLX8BA8E7gi8WGaNHEbEZKIeJC/Vopq
dejdKE1XAFlUF4ejUfI1SGzBUBTiUnuEzRS1mgKtZlWh8+rNrTIl30xWPIsnULEI+MyxO650M0sb
yrlELUQCvdxujF471gprkj45MZ8COu1UCjpMEWeyqZAhhJzrHd9OinPliRCv5wK4Uce6J5fcTZvA
rdY8V5ZR1EqEPgqGna2sz3xhPTTSmagFLEuSYQEFcKH6kc6l7z11czjMlp5Mtlh56pi1dY2tcW0c
MfAEg4+1Az3kI0lMXN3yGeHuOu0YFmTMlwcZJR7eWZ2FlLKyg/THyeChm8iXJyEv/xgbn0WENp4z
wIAWlvzU/rAq/qLVPAHoYjLiy6yFUAlSAVEBTGS8jEMvJf8vNvYvlEhOPXsXyOACPZ0GnO8dwrAs
JxgLk2fuY9AOO88cDFxuI2qdDf1t03Yd6QLXQ26EgXUHiMDIVgK2c9LYB2HlaKDl+mbUk9HrHqgu
AsAsut/lXsuLWRnRpNv00gytLHH3CrUM+/2X3LZIXhhCVQe7Owrjps9Esy1uOSYZsa2vu+tuKD/l
dwMA6AiCaGfRnVKKNdazSqctjGTCT5s2DRTHldO17VWaTJm0FQYrOWsd7KNLM/CVYZwS0WbEjAoc
PaROGbvNRcBIQqoCEq0jD5LdM9kDE9X8zEMskjQtWllpw6nMM/pUqshnCv9qO8s/GfAg+EDNA1xC
1RZzXFoS052iKhX7faKCq26Ht5mnvw+dzStiLrRipyNeTUD73VwZy6NCOCfx9wMl6CK3ea2hQm0x
lUuTuk8o8Y34ddpW1VRYg3pds8a9M3bc1Xxt+aIfYiHWp3k7LhBgsmsu+yXm8EVqaw8M3/RnshLa
2EUovYbfHN5Nk9Z6T8k=
`protect end_protected

