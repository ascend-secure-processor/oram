

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g3LZfLDDC001qBFo29vLXmnGLSvYl9wHE2E0YdHKhBM+xkINtLSAJu5a2MNt2s3WGsZZq9QDz5mg
dPBOyLE7Ew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RAjpHemxT+gJFTGub6krRYsiNLQdxBz3GbtufV+ow7hOHViekS4XCPPlpZG1EJUke11uQu3yyXfm
e/0Do2I5k1I5yQCMCgK4Zll6QUSnREFtmmZz+WTszc3Hh8QrBzk0lu3eGdYIvtmtkdlr4AeiFqXS
7p31p+PUASHPLtI9nT0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
auDxpfxyU6ZzF1anxQlNNT+2qk5AdsC0BC5dfGvOdUsrNWyzC5kdQatuQxBuux4KrOIPTv5keT1b
c//+fFGWXZVDFeT/yJxeAY+06nJGgtNpQndqVEi+railp+/RtCAN+aiDCKyNMN0OOmkZ813Q3Gyb
AnSXG+R5vHOPDlsSsZ+ejjw92y/tunJP4MHVcB2wzrwVBlSN66wLUFnIHnYHlT8XB01G7cOuTqX+
JIWEVH3QFYJzvJ4PbA7ygqkcENPONtwO8wtghJFKwMpUeCbr080ZPaJWrsLVx6fo6wRwXNQo//bG
KuF0H4PHyRuHbmdSop2tc1Bxfz91bxwZswxnAg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j+ErPhn9TPYuMWsE+GEbemk+tQQUmHTKDzXAy3ZXauMv8GUC3PKQlFnFUtXsjT+aP49+zJgwd7Tb
4ezk/eJjCBmTMkGzkA4nGh9zS3pq8JnewBIY7HGOy5fadRdFFoZmVyqLQXRy7UgDoedS/WgGbbDQ
pV+QVKkOet2wciOxXvc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZFROGrleByVdYbylYilgLKOrOp2UdSsezhBLSUJ5Pq8aYPQLzlYuItK8n+xvexgw5U+GfDCakFFm
SwJjrRIlVNzfKHE3TIpmPjnpo5TXpmRgTcLt4H3b+UjwhPd+102kVn8cA7JBdDJNbqiYg7/76H2P
yPx0yyDytNnpYudkDNKWw3bw9AHn9r4GEjoVHjqx+FldUQZH2kAM/nkKcmBB6p4Tay5PQ8m1wchS
55a7PsELsdAVzphv1NFeMmeX54aEvMMBsjmkQheBTbIk9Kw2urhytx28LUGZiylyBpRLpOh7XOZ5
qrjKmP7hIoq49pKlxS9d0ULordZlfzeX01GKrw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5008)
`protect data_block
gzyg5JEDfzB8OT3AxE7fGs7Vmm9h6M93TEtzBfQTkrifyVyvSuDh/S/YJ9kY6WlJoDhrqIAhNP4R
3I7k4OYZkzZZ9W8yeCCkdSvzhGb1AQPpc7qvoXTNciZsy7QkfHhl55SeI2b6io1gXEezHysUlUR1
19lWG/JwW97jujRZywgGs66NAlP+YOgT5ZqvdQMFeFh/XlfYKLTni2qekoML4VVRPeGmD1Cum65T
43kNDjOppOZyHRU6zL5JWHWcXL0zcS7rvM4dQTOiSuVPje/QCNM8KZKbMeZVeweD3VvMnpQ0yLww
Had7EPNvRALQEnXn6AKI90l3+f4jfK5ZYrUr3fS2TQFVdVUMKJpJlo24cwKmZzSliJS2yg16ezhV
DgtZQ9kL5nzHFB1QFvpbefj13W6MaX+LHU3dMHOblYnE2OditsUuGUOVDjwGFxyKgZjkmkPjqsM2
7194hYxvxGd76DcRytyWfjqm0iLseUySTKuTlIw+R9HT6/cdJRjbb2fWUBWwiHetucB4yNg5z6jx
6f7glha7oUbAwew1VysJMVDKPwIs3Xu0LYfB6gt8eKidT9c+r/A3qWfPl6Q9Li99onRQMSiGKAwO
lcsbUA9XUc/pMfk8wpe96/MnJwrKzDMTmx4/qk2rhmILqPA/xy+1P7Sdg3xrewHZE8gUlHWpZ+LL
wqqgcA0h9sfhRLWjffrnZMmUttBgOHGSD07DpZttHJ5wklTbiifIsPYTG71B8jbzV+fVYq5kxGQJ
fijcqFepheos+ve3K7BGjEV1ZIYuBt3EUD4Ce8k0/balRsqL8LQjUrMVZM9o0qV+dsQ01aRIUI7o
ofpXSETjvyblaHXAKeAVMQH/0c4VdanNyttbxywaw7Ttl/cHyPajXn1tED+4yuTvogiFztbPb1p3
HBp1kctey15q/LrONDOp40UrXIDnDw3+5YNXypem11YvVXRTH0g4OsfXxivv4+xL3WX85Y5oWNlK
IHaQkTgnkcxyJ0xwJfmYOTgr+4quRFhDtrb8goVwfkkhWZ4qF2NLmGz5S/PLJjJnGNvQ00lDstcg
7FdEQbmB7EFAxeU0sdbC10xNFYoI4wIbEGd/oFcmlYK4b5gwjBFFMmbZ+grKxh8O4lZijMj1G3T8
1ffqeLd2KQd2jDk82onpVm5zR6R0YKq0PCMVUuRQXa5QQAwCeW1d2Zc4dEcV9dTKOhJWEqZzO1bE
dypfA3wIlFPGwQFCLhuVjW8Hh7BoS9t3upKcNtNWIEiGXiFyiNMUNFS9XcMvyk76CNQhXJEsXNI5
JUOmUomKjzA7vR0htUCntoEf8kQ4HeoK6UNFdqN7MtPe25Q7bc9uTjBqJqMudgw3O+eeERvoRsep
G/qvW689fWzS50Be95bsRqjV7HBCzov94k64Tc+qrDmBKWWpT7YhDNBxhCt1kb+9lxwnv+PAaccP
NHwBo7jX1rFwGEOuv9ryRz28zqlu02bMJYilmpt0Bw3t7uwm1VTok5b0zLVQrTaKApnPmzTM5YPz
l0Q0iKpZ+eA5LdotNg0ouLpci+ohQ6G9pHhXFEB+/3mQ/fN9dy5aGFyiQRsULATn0+72KrQYtCSs
6ef//mzsotPNPhxGxLHml1G3/6D/4b60Skxy5CF6PGN/USMlC7kcC9TSpxKLkEIugqs9E0k5MYPf
cbLNQO24dOHmwcknUe+ewaplKZkkUFVa86oUzpcbDwh5/QOThZ7k1pSd/bgFDS1LcAmobDrlnjcC
vdYFm0C9X4+aXdyRYVvY6OILO0TPwCgF5WWA8lNz4lp7yBRlB6cc6oaxWphBhcFut/3+eppaXBgJ
YyNks+GpAcARph1glF7/VmL0Dx61+yjnAkxVa+s4K+avnA3rtesihVEKloh26B7kePKvuspLx5Np
5GCOVbaZ/J3U3o0oImxqO+GmK2LZ7R/QmuOUpYrz8p68na0KQVPCB6Cj43LLK6Zrk9gmre1QouK4
YxuwGP6kmXbOSlLr+1qSPfQsC/z96ooviMdp3uSK3gsWnFKiLtVLYTyieBOOfcEb+lIF2ipx0P/s
GfRN2ie0PlN2POrsECSq1xbHPbzITiZ5GulZuqy/0UF0u+zsKainUgx8G43TW6lAAarwNmSGw/1G
gmEFoDfPIJc4r7rbvS2pFhnZwOEslkFyA8qSan5Wwlq9PhZF3n8+7dOrBs+RjtCXkAMTmfiAyiq6
fUqZEUs6yhUCm8IaC5T8qXk5YhaoNo0s7RpAgNySKTXwdSOLbhVwgt+Bvwn0iA0A97LjP0WgYyAZ
npQYx+rGkdYQ1EfgqtWJV3CCeZRvpF0mpITayZKHS+3bHTxsxXK+SqXik1zAfJWwivDS1ud5xE9u
52blxBha7l3ea4HA92vQmEa29DBNQMfqPExCAoRweSFPYVUI6zOIhxnNCQC/dswn8trejH9ndhJu
iqu0EZJ8uKzsxfYhbp8j7r+AyuH+dt4cn1VwCiYTeAC9KdogdMCThAsle8b6x1O69GH8LG42i3vb
upbtuST2YKZ41+AEbCCETt5WaWT3JoXxjejOrVB/6KI16ebVUP83ky7efTlsLccEROdeDfyNhuh7
F1DprvXEqLMNCv2ca3afAEA9rEfcDJqc7fxuT1z+gcrKaTor3AP/F5cBdm6+F8RSdueKM/JVWott
wqWKHoEPB0AWLPo7/zLqI0sgGHHXZ4ccr0w6/ZIPmSvWUwLSm9vj7CLxk8WNkV82WrLsYS/Z3suZ
P3bW6OVaFwWp6mMFcfVSbx8NjCTYVlrsNE3xe458e6OknoQ//N+b+zqrmG5DfPE3IKNJFfX4ERwh
LKYE3CODShBtc61OLuQ/sqkTJZoZPFXH5F2deEibWhRAHgs/RagiCLtdxcFP9Fb5uv57Cyjp3k8y
IfWDDh8BLc3A9Cwdbk88CkvpfddprCzi2a3I+dV+c9tDJNRR9gzQaTJcc7GF+Xb08J/FE4WvcUDl
LAr8wtGq5vG9VQtW4u6SmYPFT06cLObMZyMzk2rqrnxl+TFmGTLIdouCdsgKnrl7Fn/PEZR9J3Vl
rphFGgR35ZJZ67YYoEm+eW68LoVPRZUoP2RWa51Elz3iYrw80//ahmnphSJ+P7ddbLxyIOLbDNRJ
D+Hu5Cp0Kj/sTojjh8CpAHGaHWPN7G2qpuwlU029t2KAz/HOSAnlDpk7oiRjKaVvyskZmndFbqtb
X8Ho8yUbnXvUK50Ld5ThOOSs4wuVQZbGaLX4kv+PBHHIzIyXNv5ebV8137anAqU2ukUprIXFAj9e
o4OT6PQ0YC6UXZhwxKroEz5dwQ3e+Lo803s3UIzQYBCrx2doPgWF/fwKcNb55wl2Ns2cn1LbMFoM
UehcfsBqmjfltH4VtJcA/KOFoFLGT8+yRwyeXmYC4c4MocdsMtQjZ6XLk6GqhUKaaX3yhL4i22y7
/1z4TEkPUef5Nmi2WDeejus7SzI6e14iK5gkLs0lcOM7xonggO8D184wHGaaZdLBnszwyWLWDl6K
+fgydTnJtyZbFaloJPTfFRgSOSAJ+kX7szqf4kGXkXSRGjCRH9DDwEAnyw6o513v+hqUzFizjbCm
MKdfW/D3dWSYXzmRlVYI2fhisbugR2rKUJ90uKbLpNk3du3r6VupOo5TyBg0dp8YH1oTCHneu+Bj
kJsDGjwqNkgl1xI9ZSNbg10ljsidC0f3imWhaVmc10TsauFs79YvEBBO67GpYuk8Vewa12oN/aHE
2kVIExPaGAhCky5cBLH20mPeBlTr/AvppZ1SIBmw4X4+M1/s4zhuNKXu4LMJ0gQNSzTEyUfv/fWe
ESGaLh6kCaAhmBw6pJ7wGxQzi90RRUdy9i9HvHhbNhkEYL01bDAsExvUxjRQzYuns+ChYAuiMffi
5PbeM8pE0DGpn7RguIjLvbEFdnRcSEFSrfoyA3F2QxN31u2XayQzJEIUXVVHS9ixTLDRaFzO523F
4khLPvA77Oi5ypTWV7fIo+4n6fmyS2GsVo1h0HRFJROgN5+26JCa+376l40S4GGst0KjwipwnGvX
hZAnYVFOdv1Tm2xNf7NfFXtYBNb05kPl6yvl638p0VpP+zPwG3VLCP9p5IFPcENIpa5Xwg+83/US
COcqIMYyw3FkWKzHbOwMW3y8HWaOi01+g1nWk0F37U95FDqy+G7zVgzyRuekjbc6Zbbcfp8hQb/O
CU1ONYkDoPX2AUznem+KGAZ2HALapLqzjzssiLMJFrKby7gBUJJhN9r2IytVlQsrvQq9/xURQ1a8
+t0rYWL7Jillt0AQbi2z+amfOehjSRw5Q1c57cq7shDzNyRDY2o7j+oMR/1T4ncYkqPsGl9Mr5QV
UMbmPmVZRSnMcREww3pS4Tmo9wlFWnRfkApJKOPeON3kLwFh9iIenGwZgqXc/jdTdK1UcBJroLFB
5Hd5M8T8+iQzBBxwxJRIiRkMKpaFEpTUZzRgvyZFnb/LuxVksOGbMe6a1v56YFVxVK2sqCjJF7ae
yTS3Jfd7+uvoLvHYHiYLGowaACX7kFOqbbnHRJQQXJNg4ATvUB+btBhUs0TqoqLjCY+g/aMB4lp0
gM+PMgOK/1izSWaAviR601xqKGa9DDD2SzvEsYYA9WAj+ZqG/Z72hm9D9dvj9LFvZg5QQ2WrXioi
MfZPQpwOffoCXtPbBlC/TaxPtjCrbd66AXVlv3yb1uJFFNHK27zLkf1k5Ycbjk1Wv83qfdySKQ10
J+NE9FpDHTqFyoujppgJHuSudMQKOMjP2QNwI+XI9s1owo2ou0PF96ej0QZTZPazGCv4bwRV27qG
1PHayC8PyfW8YkUx/bfQHDbpzw6zlxqEDdyQJIevHdJWjdO7tdn/AQ94sqXyyxrULrrr6+a3m9LL
mXbhCEgvZq+G/j3EKYo3u0/HUMHUjNBPR0hNMHtFUIf0sxL9m3NAnwMrQm6J2XqugKmCcq9JOCDK
x6XMGmIdBtWUBSzfwNlXVxzHqBvUerERjSKyneN4SyeTjOoOI9aJMp4bgen+2DZs96X40IK0gVrP
iOITsO6mGKa9CWyIeRC6+BEdgfh7oQCG0um5o6CfkSwfH6ZZ9CxWWHwDTYFG6FaqcZgqGcxmPOWy
LJ28Djz17gHNHyYI7okOnVA7NuIHB6LAp82HauHZEgF9hplumGsJRwNB4ayu0RD6ExZLwdACHhmK
GxXHvVC9Pn2GpFjC8LxkxaDS+NDcf2fzSoMP0P7oN2grFPgxjkNbwcMX3/As2JSyCMPThBqCGwsQ
7ZQ9HhhP/5w9Ey5VbSuWvXk7bp+VDD1v/s54RwlAJXGbifoIU+3ReK4JBiwJSt82D0GosNHQMgSU
9v1bsV7jITlCH2mhOXnh4sTKHT5sh24ouGKK1kNPCZrYoiVpvj+aAF7C9MJ2sRm9VJiT4EweEDde
lol4h6kx5EQiezyqfZdNLwS0m5056+fJf04Ba+FR0dodOo9KB+ghqu5HIaQueGBqWJzt/ws0Iu9C
R1xC5bUNvaRvbtFkwD8Cy/6pZYpO+yjCds+aiDjL7z6c7XNWY0PDYSW/TeOxYVUrQtANFumzhxaf
VeN1uFqoE+/md2NlHxI4wmt6TL7R1FLN0XdpxOKjUgcrUwdHdvqBCshOAy91mTWoMqJujUaRnjQM
oDlOBCA0VrLtyWPWV2uqyXaoqr6GNnWdn5yVlFd95Qq4wXBzXSz/c9+Ywelx6leLRoe6Az47yt7h
eznjZ+Vy5p7jKXI94SjU36mnqiUNxccuhgoS7MPGBAVu9z8mCmZPUlHoBnooazxifw1gIPZRumD8
4xaB+g6o8vV7d7XUM64yAVtbjg7anm307V5U02Cz+XzmWk2sHYO/QHaDRXtwScmN34lytAO9/v3m
EI8SINja2NPKvhJec/QnK5wcAyAWFQTKWlhfmodFLj8FYwIk0NTgFBRU5XutnnQYDmWbCRsOMF3F
utAd02Ifbwa1OeVW7tMSP/fUCW3LPbAdyj9rZJacGmpm2MsdGNfVj68SwdM4z69xbHr7oOGpEmj5
DHYDXoc9KTdWU5l/vfSAyra8rYNN20DFMJl4+HK31anrrJexujpAwLP5r4al7cB/313sCA94XZ1t
+xlDTx4+MY3cYAeNyN9DfqmUjdczj3igCf419Qz9X5tuDD1TCcNNwXns26SKIOrXP0MuXUhTCQl0
SucWtLU2XYcxH9OZViNp64ODFay0D/x7SNxQKo4yELS2MClv9/yH59ZnMS2w6NGGKld+h7Pu+xfq
M3zZwhgERXQCFnygmUdas496XJw6PHWcUcyOZ2bmZ4Ac0soiOIHo1Cnt9A38AJJ/t1U8gWuAcQ97
4tC61onB4zZoUOGAbjY0czW8RsNUck1M4t84ZnC5ReDyDoemOB3oChsguX55SVed49eCxCEGHn6M
OarfBAVedyIU/sP8tntyDaiJYe+suwaAxWWXiWZu+J83DsgDeTOpJ/QKpghe7rAHhubEQX7289Nm
fL7saSI1GtRUiQjJeC2LdQjmSv8rNYcILXaFf/K50ZPoSzFiur/nGK16k0OcJnd6wkqEHxJa4Lzs
3uqhb8Rj7ohJ+eeVcNFal3OsC4OuXQK3bfWDAhoO2FQQ+AE1EoPoX39EwuARo3DDvUqUyA9UjJ5r
rofbi3uZPZ/0Eg2Zo9hDveFc89GVWg9muWck0056Rz2768KKv9nwEjgS7uZQIYRLAA==
`protect end_protected

