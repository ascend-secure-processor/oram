

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P3KUeoIXIK/J3wTz/ZCRx5eRtD5DhfNNXtHLoVtTodDCu/7pZVeUU1QLpES8rqBKiuBNt9hJbCje
6oWMMODr8g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PPo1YcMlwic8rtWpX7rBTRz3lAhEOHzwynxhGecVdaO1qnPsW7tizXYOFOwNpe8sL7qIGA+zbeJ5
WrSqlHThIMKrfi/0uTwJDmNOIDbb2WK7AZY246fodH9wuHvDTx1j1ZrMTqOerzY0NHa43bJU5uFb
kxCgtd9LsWkP68Ezz8E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dEoUTfnILuUdg6PdaR41SFSgPpxu8EdnniCcN0F5mRYX238GAJC3QLpSuOajuxNHmt58sBS6IqBf
DJtcmyqyTGjXBFXJZZXhpR/eabd+VEK5rHiqaB/9vYpGEdQ+xjbgTdzh+AcmtQ7NWvNFfbTA299N
niHN9k2+csx3TQ7Dh19KSY2T2/swsaXl6yxaSFJa/VMtUSbb1lpKPyxhQ3gpllkvN92C8oOgV0Co
q6ZKmNgDIhKgx/+mne45AQvCtlQrnZaRxLCDi1/VQD8L6dsRWWJzPgdnOrXX/bMIM1BPqiRMbICP
OU+AJX9n/46HgZNzggLtTbSMsVwYhM4lHCSbKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TGBjvkNTgy9rZxc8UcnovkLSrb/zttR8esIKPvvMU+LZ3hCkM1ToJz4n0Qm/xWO0pfPEy0N9KnKP
OX+47sOJmiVkmDc8kIROnCyJIff6AZ/LEktsQ4zxDhtOUpRl9MgnrV9Ih5Dz3V2RrfNDuXQVVmEi
M/dW9S6Fp+yVBa6h2pA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YA6mFVm8aq3plffXWE9/iFtoGeYFE5Bw/+h4QzP2+YOWoEfBuhvnyacmiWduwiLCFran2PYj0x6o
bwvWQdcIY9KXi66jnhK8zoo65HG2c0aEBDRmrerRrtK7Loo+vJlhQFLTdQSmC+VVKgTWGv9QHUfj
Tc48Kh1mTQtN9So8Oz6I/sTyuXohDdWZlDpWuZCHNEZgyyBq+dTtOawwLcyPjdF6roiEo5AeHQoC
ahOtWeXmfvKcCOOIXxc4Jar1BOzPGAjSU3r7hdEghc93LvYFuX1OEhJNnH71XIMh3XKuOBzIYKI4
NpPZnf/HDiosZ/1zkx2grc9oc+2vljzgMXhQwA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 158432)
`protect data_block
0Cx9ZLwgR+TObwG7D7xE5EOJiJA/NJP3+HnphYaBXYVBb3RRLaQM8ngK/98iz5qqTLA0ufl1Vkya
jK7dALelFOTTw5wxcJSI/58cyAl+khuP7JzcHAfauRi1UasphClMVVEBDDZlX5N/RYGYrYVVXVmk
e6SiPWEmi3N3feQ/0lAwejCQ72SvJeGJOwiUJuBod0EI89L4x2KzreiTPj+LmXVZ6eFK4wlRhhB7
EK/3t1vxoIOUgAOFH3vlBjDgyhaSkjyFFwazVKooISG6qd1R2f0JnSKnzncunhEWl+sM8+fuXKYm
+aCPcozc9GHIFrAX0ib+HUA5ZiaYxY4NthMhB5QmIutHxUScNOD4lLQkBydlRUmy3uEijie9V6hR
HRfX9u+N3uKWDXfLeCCnjF2jzD39x1+DrljnANp/VfcG35MSz3N09zrjZgT87iwOX4XoVHOa/VFJ
og83s2mgeYNZw7v01zDal0Tr1FYhDH6CsXSjgygC8MucUf20IFyove2qVwHv7e5OI4HVkvlMbKI/
7csJcRnqTj1hKX8n143n5Mg0ZlRxVsaPp8O6Fpcn3i5Wg1WWlrlhNxYgG6nP30TQUQvE4u5OxFL5
tUjZEJhjhH6O3HUxA1Bgfh3EFV5c718zxf5Vc0Z3g3PtedFN+Dy+15VtoOnkdtzQoHAIYz39z3NX
KRQL2f9FtbIm85f4x5DEC9GFq8k6X+nWV3YILAcQuHdVDppw2nlP/gdAvK1PGQES30gkvfrEkV1T
u9g6cwnQ9o+c5WtvxnZpJkJSkF8C5x3ujoieThFDKFChmj8RKCQADRL6e7h7ju7jI8YwFg9beBE8
zmnnTXnv+ujGfH3Y7oiAXSx2+blT/Tmh1CSZ8oaHFeCAAG/Z30/Sqx6mcHS1EWhUnLNq7Fbsdbp0
saxY+dPDayoBjcEp7mUICV7ES6sUQ6xlyLZuOKScnKSQA8/IJkAhlqURyeF7m1x/AFs9WGePnJdk
NKZsdlkPHsfzXyDzG7oMBgFQpiuUrhZ6ZgoRtzyNanBmi9QRr2MuBU3tNOrOsb4EcSri6Xlw5qev
X90AHedwo1kiDETxjJbbH+GfVh7YCC88OlqjkrnS4I/mi07YK3kjHoaZQX0YTCnro3dceIqYNtYp
eQsbj367rJtTH9meNiN+GgnEdQlHUdbXsgdCwlZ50I+tewqbcBKl31g4u/WGenUeOIP0wGXSeLmX
d3WnDf3P7ezP8B7oIji7lNuIpgedoWqNC5L3R4RgBtHBWFa8Mi/MEO7s5OeDL3dzYO6H4umS01zL
pIPNg03AnVOzoq1dvWXK5I4ebZWj+P+HpEMWylplJ74cVSK0wkKGAVHtwprAJ/UslA/QaAXwMtoo
wF1qNc9PPRjcsT1wCbD/qZXwIsE7Bmm0jCqU3rv0W82fKgzMlMd+y/PSP3J5BXxVpSDBeRA92Awv
GRr8oFYHtouvLLm9YVTVQhrRwusZi59IVzgtRZVN97s4mkpFwdZzlQp7Pe7oY5e+ISTX+XY8t80z
ne+CLwRwcze0KKtjs5UbdOg5KuL+JGUHzz5/vabn5CvW1+hVoGbIVvB5xYYO+doOrg5nhbLBFwKY
DF75iH+dl1xZY8WJpWwy59rGNYuwuZhm/CLT06hEaDmeGqx5tud5/ezocg0teDp0ACiI9oGg2lJT
+bj9IIxXeVEoWrkWJvhqJCku9O23Rt9vEZg+1H1M5W+hCnbXChJ6Jt0VK+I9aaH5jKXss+c+3XIT
583MLVaxsXVYe1G6qfPZ30E909z6vR2XN0PLUHEGJkLvz7mY/QBa6aiZkaG7iQ2tQL4hNRPKjbpr
DfitqNoQi3maMLVFjhcBRtqiOBJB+u9YJUf5xVS8YIyDNqlkNsyI61GdYidt6VA9AgeiiuTusLhw
9Tn/cSLZaWe9aXuTPtz8RMrM5pOg/VLczUKYzjpyuEy1e+VTPkvWMjhvWF8fhLjnhvRYilapTXY5
m7U3vKp/LIr+bpweX+ZulunYgXLfioLWn8sAKKXXK0lEY/unvqRjqiLo0s3Ppfwdc4aSOPbvmSSo
zG1NwTrSAP7BDG9AW9kimKUR0JwPgeKiSyil3ma6pTOSJFLpIe007k64sRNobs512Tx7kN1fLqDu
1Y698yCpGf/WbP9kqnQ/yk1O2X2OwzmDbYjB6C6X7UiQKc6H58ph+PJTd1bdy9ZUfIEXiTgNOxgM
dKzqpm1TJ+CsQPRA8f8Y+nf7RFa4tjfrKTCbdOub9V4jb2K2XDxlSEemeh5bp1/jhgynunS50qJ2
b0dKxtYhiIu6u71Rg4K0em17vrcsxCiPqixLsxUGXWkb0DMDDxxH6XvLiqctBaMeujd2tAVq+IHT
pT57o0sTgTJRXuKpYEDYQghvAB21142b1EK+REHQxwm3T6qLvcYzBgZDBvzG/WGRQQ4jbjai6Ban
eVIu2Ks6ovKAVN3ucw9oYz1aYImOBh2YFjQSmJSCVQnxrwIKnXjWoVX1A6cYLjFMq7TU44OxmMXt
l2whxtrYTbk1k0RsVtFm2biVcxNu//PexjN3T+BhSDYEepn/zsTnLR/5SlFm2tM9W5PTKx1YFGro
hYxysxtqP2W8OnjeJnPOiIXG25vxZz+/q7Y8hbADYpWH7nFG92E2WmFRsDYPSGImxebtcTlCeUh7
N4xN3Cuw9EgP5w9vqCc9S1bw34Zz1v8vXKKwvnO+z+UnkyqunDPJTYgqja/XwmCpunwJgnm6rxSL
KOWzLMYWl0ywnxkvCgcGhhFpaKmTJYXuEjy+nbBE+WME1aBux0eFqo6LsWRs9F976weHU1S8EbyD
49Fp6mwur4JeIRtksP2a6ijm4M2fUjt5PnjTCVMV3eImLOEdDpLij0DtvXmFPVkuUU/FTbecrz2s
YIGUFuJzRcCDYGfPZfFW2AC2YCC9ecyt038Po8OHKBQutNjY3lIyZOvOg0KSwatQq+pRuZ4gFqnS
4FZHT/JJtaqk1ncOBMF0/1h3ethva4O4ElpDmr7sfpqi3HL/A4wq58WWoCx9H3RvkUHP8N2ftehB
almS0H6GwoUs+QyfFjId839nJnc4v2uAMi7XkFJiMycBMg3+gLxKKMkO5HGvysdMeMnzGSc/BHe/
+2pIWe4cQEYlIWVTJchkQN+b+mR376EdMDUcbV5ylmqp5jZq9nrp+U9Sqo3lFe6EMkYdmZcjp1re
NxzZeyoWEnXEV04jGsygu8NrRk0EosgVjNIOxzWR+NwQW29bM3tPBN91dIlwZng4PiBvNASaBdmr
n43ViEFSuticU5VPrSoW2TdLhTtKOCgB5VVn73lEN6pxne1r3wOsUTDQAIHsZITtgw2yPz/KbXR7
HtByDm6YbAs1IjrtMSRWqLHlrmRr+qesKoxs3VTlRpq2fbmZ2JEO595LtidFq9J+bY9rTY+FkdIc
nguPad36X6xdm5C1FG2sJENCAPq022Oujmf+pWRquI6ENqOm7hw5VrAIb4Vfe8x5hNtqjR0pVymL
f4JrPVzW4XUMyD0UdxS26qoHMz3MDtbhlGpGloM3FaAdz9SPOGUsf56/QKd9Du5M3hYoSyUpLl+I
l8w5He0BTYYYVfJ1HKOvfwjh94lXH04aloNQaCr5NQhdtxd/ArMp0c2JLegkjW4Es48IU/fDK55O
p5qkYweuGpEsQwIG6CH2mIZ2WCKeNLAPeJ7Klbaw33FkfcbFduFuYSX1qEJFicSV3DkS1elKkUhx
T8sW2PqwTU35rfjqmxamgHfyJ9Mlx2p62u2YFkB6OX7ADwePNMtkEDr3Awf14wPQzL7dp1zh7Ak7
3S1fNxEOte72U2eK48SUbi6eFUZQVyOvbOTN5CuwQ8HWbdxG3uUXp5Ldrh+MOSCThamBnU7WVyof
BIIo/VT5E0RfyFxMyNXJS9JehAxK48aIvlsIg7OMyocW9JXMdA9Ipw96dPhjkPxHb8tSwPSxaPnb
HNb48h/qGLyGcKM6KRdrAXxecalant6qAoGVRCnJgkz2afG60qef0gw86LfcEvL2Z1Z7CbDeH7yq
t/eGMx5FhPOnK0kYC1+682SjRD+nJiHzzGpaI+aNTPi7IxVib7H33e1owqIJm2ZnhH01o65AhUzv
DuGEdSjBIXtXFUN32JrLn7j07TRZvLkoiKQr6uxZfU1TaW6Ey8jQrwMejj00R7uJh+HhuxSy/gkr
KQ2AbCCdfCvGasAmfy/gqpM4E8eRQ/OolTIRbhgDtPO5ckHoS3O2+rUI7sgKSWRf9RFSlyvRlhBv
MJOEtoK5fQpQoO6Qpo30VHQk0En06X/ynF0IGFJP2axOXBu39n16PnraVXGeE97t5hHSCci1Dfh6
6I+SOIOOKtpLcwogODxhD3SCjOsQlCAQHwMI7Af98oWTeCrCGvDycpa98zXtOp6pN8ow2aIRNJgT
N86JinNAVDZZH6pYAE3XZL95yT/tGCPjMBEQiXslJ47p3xCeGa17iNflA3scRbB47+zQ3Eaw7whj
NijpAtoITIlL45unqVyMxjHX24c6edTfBoxv0FXz/d0V4M8sIxsuJrZB177nGSeOcPcm+BM8DPad
e/mhyZ5Nm1fvLkp/ak9uQYYl7PJjSf2PDBLSqd9YKhH0pK9+47yO4ql2BDt1KWYhfJoLLwMrAZ1v
FsasmK5+kDg4HIr+xymiKFavYx6eDYKuUMHskiyf25w6Q7LgaklRNtZ2il/wMNXIWCfc4oUJ9IPs
Gn33fS20bCxjlNIC6o2x81cAEVcG3AMo3eO6vgFCZxqZ/XLbmyA3dl+Ryye3HfqILb9uWkuhmEhC
+3x/E4OZPj2h6dYwmLus/QRlQE/f2k4ZvwVdCsHUOqBtEf/slqVI3aNnUekUSAfQYksLtJx6VAvw
NJAQSwHPfqOyHcPJfrRuIFm3z/ZdAsMlF3rbKd5OWGljzOpTxLCzkE4BQdUJ+TYYTlLqg4LU7GuR
gRQGmQH5C/bectSe9FXKKyMJXI0oZvqesz06oVPqyBvOwY+e7vJRqaxF/ReGm7bMM5t8mQAilRVU
G4EnzpLlBuMO0HANw8Rvk22swxL2nexlizZC5SZNhrdOZOfqpBooPnTbxOnSrXkjYKXqtQxcn56/
DQzX1oKVDUTKXGqgj+0tSrhS4LPwKgiIK4uYRtHOtXXZPWzkvlAyeslRIxSFmCz5lQpdeMCSxCM3
u4grWhNdD7/2ld35L4XDToypiWHT6VNxb138wnMi7RE16IQn6JhkEtmM9yGso3b6ZNcPSu904LBP
YuwhXLzxGKHXuAkcvi2aCnXdXMOyd9O6TBXWn9wmclWDGrPSpCFiVCejnllyrNViyLpBU2Zl7Yct
VuPsLVdv+o8vHiwCO5cK0h9cln6AGfnWHvXAdRf/+kqqGoEJ4WyEjIPyGqUJ4Hwazt1wUxfWiYyw
h/soWt7X+U0Hg6SVdJqbGVnPKjn7703/qtAliPbQP0veS9cSwu1+2FdSePITcUy9Wj/9JQx9djJu
0NTbOjWuYA3qd1/+Ju7YCmQWklW85yxL55aAEj2vvsHzPVwKg6ltMKmwCsBjdaafeVSURdgldJtx
Q0FnK2mJtsodXgJdFIIlFXJgGtX+AnQE3RbDJspS7ossyom7y/kXNQ1s2BZ391bTodv/GTZZ7VTk
Vwg5xphnRaYb0eCE036Kz3wqd154jAHPSvtrjLz9aVTmmVqb/sYV+ml9b4IMnzS/ocqW134Y8DHH
ZbbGQzmH+WKRomfhoiSZ0Ak/9EVEASgMy2oeTr3TrHTOEX5JqFMog6PNsUpz6SBOF1DSBnjH8Ot7
kzjlFrzzngEC/f6DGP5hxs2QK2l/jPMgW7reTmHSaqqSWF6DX5lmX3XF9jLACc1DQdhk3cP+q4qM
QITYtgRd/hDdNPJ+DJkepAobiGuTHYERcJnT+PD515PBEBYgS+9owolFz8VzObQC7N6XnZiIeIGX
e8Ci9T1NwBxv9YPEVTagBVlKXDq2IOeOpjQsqohxO7WSoMfWTkViBZe5bYCYQs7IbZTAUQk31d01
yAataXDsb53hqMnkNfHzSGPZqI+AsA/HN1l036Bl8WJVt5x61vfZ8XZ86TgzflUDvYWaKfkLqibw
KCAZH16lxtOPwcWURu2/5w7P5+DE0fDn4XaWHELt74SkSSWN++D0i427S5PRQR65kYeB9agDAvAL
00QeYuwLWRBxWKgRsdFWawGFQ7U49D5ODTIYLko2hiu/0K4k2/L0dQKDjKFtW9XBt1z7AlNwQBRz
ZYit9hZKYU4oqCqPQm2qt6IkcKzm7G8EqAAQqSh2ROc8D2ofR6QMGU+xD5TqpSM7VoeTkJElXmWM
A+jl3LoWWvroUqTt6UhYT2pxgNsb5d3ZP5fm0Lo+nABRa1pmZd8jAGi3eis9ntojM+ao8k+JvCN/
5vn9o9NFNcGgoW87IH14KOc83Ic1nYLYsqvFCLu6KkqTV1m+mBVHPDE5bxqdfin4gtElFZIuDOV7
eZVfTtav9ZvZ/QEId2H2FKm2B1IZFD9wRREw8wnthWW4uL3PJZrelQC7V/n9NNI2sAaLWcWPDgce
rbZhs1ePEzTG+5TyWX187Vs2YfblfbxOHZA3+dwhxcYcOroAEJcTEdfEQ2FlRHfYLp0l/x+qxqej
cPs+bwYmr47bp6vD0Vb3kFeuYSiCut3jyigHHLaQzPCvBLYuCFBNYgz9c7jtbdRmWF+htC5+steM
x0Vq5+msF4JeLHfY4VfjAb5duk/Rb3ASp9CbZcvJ1v7BueXkRZ9avDrtCBD4UHy+t5hjk2GL5q6x
OgL7QQSs4+lSFjpKG6rZDgtfUKAadLL9g5NFmEr9T6exhh5ZE3yZ3nay1zuCj/F/1Kr1BibThhjL
wbbclOUKYVdM+iOtduW0uo5oNmlvNIvetkcVmKzPfUflUC7K3U/c4RZb8ulssGAOXICun56esE+E
qcHy0fk4vxFKWRMkQb/Z/jbBGpud29uumByVWIYElK2dZZ8e2JZM//txKuTauHm4ng0mq+N7DxUY
j8mZy8fCbWwsC774MakZsCXl7zYyMZ5koTy97VXD2e8WmFMNsVrxc2XqGYqEMiTNJoyFe/6wzwu5
HF5Yd3EK1kao+4yCWpN/DTGCvXWFa3i/LRcLyf6B6a4622PDj6bFyyL7dpbC36VCFoy+F/UNEOPF
j2e1shbMiLAvmrwnub+hQjfqeCuXvuAU3ORVsbFV0jrPsY8Bl+03hPyEM0+hchsB+yNl6NPGdDOQ
UbnDMTdQTS+tUull7UfydSkfN0EnBPlbtxX2s6Ds8vf4MOrlYCPkefrqlhzSH/sclOmKrYIiDX/N
sNGACvGTrjcqmnj3yDFRx9wUA9m8GJBZICgWN0Mv5Wxpvnja0IYNe2gdU3x4HtnZBd4jIDjaa2c9
t8vg1NuT4vdEC3sJwkpRFCFoomaD3ekHwnbNksExAxp25PuxTlbZGarFxafWJagk+4UO7WeUPv3g
ijbLPuMqfHIp9ZjlzVIRhSc0gwbYGi93sjU0H98zf4xk0wQFwkxnQwKWeS+E/9liqXwc4lxKjkSn
Gq3VKDprsWy6iJTZtV1MVWpOLjb3xLgLPYSVOcRfQJWtFMaZBPfy+2UyPIPkU6c3NncyOY4DKxo7
iwWv0zLGcMFdJPbsVtvdDiq//ZZcBziQR7766ddR70ryFHR2Sb6b4cFYdlhcr+6R6EI7eUSMhGPW
SY2d/hnH5zFT7yWnrSUHm11sS82pqq8QN2kH53ys24zZ4NE/L0JPUWjD9Jm4YGdiQxLZaCYPUuDl
zhp38pEtH7ZA3SrqI4+b+w+J7/+vTdvwgLlNpUyOdN18gj1VVi5gHlESEw+R8RvsD5VFDg7MsJci
ouvxb0MXwUra24yvpdsP3UTBflpZkYjCfSfbwLdlTYgcPO+V4VUpkKpPjBQYomCxxFdRDaO6yWWB
8IzrPZlVWZ2W5Dix8AfEkz986wzX4fXOfHXuSb0KhWNmX++nfzUUlDMjic6xT82X9ybvGNvgUkT9
CI7FmDDh37SINQKvYpyKw+yqpRr0L4/FoppYMyDIcWmhiOyxF1AUEVuVms9wCXC33VkFAUwNwU+G
9luKwRB1nBh9s+U2zrz0bJemUpO/qyWxbcM55pLZ8JlntTzGMQ2B1VBno22qWUiP48TJmbOxZPvY
HPvZ0SfK8fGs7GLBLiuZ4aYsiABQIUkvtDAxkooT9lvujX3LjaEq6IJdsngxxbZjDbeYMPxcljHc
X8uCSR0Jk44FJSvMvZEZLW1swOrgbCIXrXwPPNG2sNdlOjbGhd0lN0c0ZtsrDRig+p8dD2LLakZP
MtkNl85jmd4cqvbryOwZ+JKZzI/+GlH5+i8FkiaaA6WSqwN4ikAp3LH8UxYxNTpljGdsNBREKeCf
rDjS2sjpv4vEfFPQBFhl2gF1qLZt/tg1FDMTfTnoSnsYRTQ3zPnASO5GXzL4KVVa4L3533DlAeD4
3o/AQDpFQFN+ODZbDWang66vbEh+RzK9gavw3S3pq2diTD48OPSzj1fFfGiFoWzvJZpuVrOHDLBN
mtgpIj3xK9Wp8PTgf7VKau3iM9aB5byMkBrUbz9DX21Uq8Z4CE9XOXncwoVNzIynGh+MdUkPC7eW
weqC7m9qduNr7OvWve0C05eIrFqwiaSJSlzMYWpsJi0/ndkQ/sNmnvnCegYXOSR0EnT8dBXE00td
FknSYLcVvPxpfaW1Xp5gMD2yt10eNXhAnBtLIFzR/QvruE/WSnejbfwT2EWHjIRDB8CnSiMLfwRj
NG5eY3WvPssN/u8Sd4KfTWzjsIyqRtqTICZI2SFgQOrVfHix/BLBpCTROKGw1HpGCEo+SCw4v0PV
kVGqpa2FIfhjWhM8BOjIGVapoYZaUJTR45VnXViivKCZQKo8UQUEnDba3DxlLhgage/3UAHLTRhg
6hUBqMAo5BtPliDZmR6FLPawpH9wXbx3EBUql6tSHKetV+3XgEDCXyjTxohXnN6GmGr2DT+mVxti
cvR9bixR/Bxmk+pyyV0DP9O13WFHnqJEmkcibD0qCzgCJqBnrQtcKe9ZnTkvO1q9Wx3pvL/1AoWf
zMaZOOEVAf/xyfZQziay0BAWSOPK11O5wPUCXvech2HCCvWJw9VVYfRu2Q+UbbM20doftBIo1RjY
+9Tj+vo5KT7nqvfY0FBgfBfun7LcWNs3x70nGbYvPs6R6RDH+Vz8R2K/d4KUdFxGGUrep0Gz4XW3
eInWYmbUqYsRTqoNxOG8JTDSiVfFNlP0KU2QmAWamDxWTtrJfd9EAon2wrgEfuuRRmtYspaqOEcQ
mAjDVGvDAPevUzxjVWvVC2KIc1iU2fwWm/4+5uj8UDb+JR7da8Fc0etAYBVn234BxQ+Pp/8tLMyh
UWfPXoWk8QU0+i3AF3b3Y+ygHwtmTOxFqIcXf9M07HvaXn6Eqd9xfto43tnqkGNMQGhq2e0nJwpA
eRN6q3iWxvXXL2E8a/u/+QxM9M1CvCvxqRy0f1rCS1hBA+pF/2U5LZe/mlm7KkiSi4uUSQHiCdaF
DuixiPnEKWVXWytpSzRYjyOxVoUXhFq8ZKlPq/8Jqhaa/Ph0MuDpnRHFrkmi1BJNJzpuuoSlpUBp
MAP8TW7nQ4X3/caj5gofchqSwaowHn1QTB8hMi0grkrozrXlFTKuvTa3GZUQVpNmIw5LBz6pL6bs
V3dWH+W5yvFHHp9g9smR6WTc/O083e3hXdc2xRmgPor2dIBSPWgfm+g7a/i9C9j4Zi94hyH59hts
hx7JiFkOGtiDPJCgPqsfYG5Jqi9fbtuZLohus1XvnL9akSx6bILWFC2S3yueP7Py+rUgwOvY00TO
Lk3lA2bEftrXsXiPIqdsYd4BTD3+whfTucKvOfQQQQQxj8t7OhO7q6ZUBbpDIvi+WRnmOTuvGRjn
gWfWhvp++pJkwk2nV+03mxDWgZExak1w9Qm5+OduZKw2+4cXQLd4a5w6IYxzWEwCIOAzcxt2hHtM
WzluOOniyCx/CBXMBj+SgwSljgn8DXoMVDCBPUqhls++yeWnAUPiQPZnQ/5ftpKlYYs4LbHX3mD4
flGDySQRJ5gdAqVNT0uHADor/x6Hht713obFLbR2/36JTTFSS7IMyXrwGZK6pFb0rQWbvxKjOSyJ
Dkfd7W9viLV6Qxt9Zqons8FIULjugRF05+vdmgJBow/zTyuvUOeS+tZKt2GASluHt2WenQx8WGMz
zPtRp2AzjRnPthOkJOhHJEZBW0GbxpBUm7XcrpGDGGuGc55IEE9m9dFiviw9TIBIkzBU5X+Ng9s8
ZYYgZwcIkZWaV75Jsc1g0wqcDn7fUcyseNFWvZ4Ic6EFHwIpVR8Qj6tZIGKJ0/nK5mdPeX3w0M+n
srO/IZsp8G9VEsimswl+BPYka2MpmaHpROfqjSFmQikYPKhwZ0DvZWG8d/BTDWes5Ehtu4/dJqaP
BRY00cm+nJwHc1CA/3xHNzOmV6ml96PE14twuiOyx+51Ho+3G06NYMWYjslLV4IFZ1YwFJ5l56g4
cvVnE7EIo64xQ5Y0eVOf6+eWSE3qY7Ugp5n1vtCaqUPjvAZYPG7oaKmDZ+FaCmKiTxTxaDxCGrop
HO4QRncieVkPz0PeizzbL2vd2SlPovcm0EXIh/c9XMGVPCOlp5TbIb+uBioJYSmPM/oF7zKizEw1
/vMvqwc5oYWQ34WEJGU4p6OPo2hvET0u2xPbfxzdp7Pg1kVHV3PMt05NMN0vMsZaKzwPlt3VzJSu
BSbFkhKqsdD3TnqPpMYm+ksdMcEY9b3QX9ZQPwsxb9nvTnLHsoqvOpaf9/3IiIXQEWsB6HlCyzcK
laQnIAB32G/hOmKlMNo0szPpLN4OSIcyKWd5fO6Z9S5TcgaiMpDt1X65X3mQjb7eL101c+WNEBHl
etsvtEE/0U7AG/mKkY62nwrKTR9A8J3gaC8QwYsEr7nQ0igU/M0DqYYY3tvM+Xk7skMF+hFhwxu5
4lF74u8eEYhdITN55cvg/lAjFEjaRtE2nJRomp9P7fmx+6UqqwwUkRq94PlQPrv/Q+ut877n/tf+
cGIh6Z0qNTtu4Bz70k8a/NgK0Im96KQ/k7vs2lmsKkOzLdMPfveWthoLtGDpyfCCY/S2bEwCF7fE
oZ7YdHq/S8/EuTcEuOUj5um6hWtXUofGjBcIkSCiUnKP00wShNwGUFk3Xs6Q6D7HN6xA5XQD5mCF
FW7yYCCIu2EU7nWuBQg85kcs+KFPnNUjjMXmnsls+iWcoXuDJYdeXriLw/53R4XnpSJeaFjOIMaa
4qtQ3aJz2SxfKFzfRPBj6yHRHC02tcJvIZppfb2dvgt0obp7Id/oxxOquO6SvYnrbanm43NPIjUT
yxr4p0TUHD6MIpqBHj0AZB8tRBiLSv+AqzJ0DBqSIe3HAYN5Tae/ciJfHzsS2xBlF+3608gnJv/T
yurIu6kip/pqB4yviAM3u6o+NXMTkSb6Y3Ar6mPmqRiPwlW1pgDNYDVswvR3CaLwjWTdEbXbkaZB
mhS0aj35lA3+ZDnNONSuPUw4z5z68rL8ejtlyajkHFj5pV3+lKSsUfstpy/Ns0BiCBhLmxqK2wSC
NojOTm4PNN1bxDw3hOjRM4yti0d17uIf74ZNuqolyglh/JacJXRp0vvJCQoVdTOetNvop+zHOOok
7/zNr+cKGc/pJFGBbIa/yUMSk+PL776uzz5BOnrtcWPDF8YGaChwdLz1IGk9fft0mv/rSj3O7Bpc
zVAE8nZ1h1eGBgFZH/al8yfX46gN+hzarK362W1pc2l/aixZUwDbccU4YFPIWCijMGpuPzCt12kL
HGkDPRDW1UsviMd4CT3aogva4R01o3oHxls4cQInH9QgXZ5Ri2sK86dRAVrVMjdUTzffau4+g8GG
6v7Dpbw2o2pT1X4cHfBUeAnbBycn3jJ4OOcMRfrtkBez+hb0h6kdhxjyY9ejMQv+VTZjqdLzv7in
TsIRot6ej4WdWuYK/PZq2oE3Io/sE/kmmYh7KgXwYn8oAiK3m6Er32exmZADwlQipfRsM6jWCiKe
dO/3k4+0d40r/eYiupqNlTWcgTwvoKBSbo/wxc5oKrNDkgIlEVi0UrKIBLejn+daRGWlc2R9IptT
4gCNMoUuv7n8PDF8b+C1/9wo1AvUG90q/n04c8Vjbcfs9+eNE1EodQqUOqHN9E8oCp3S+SoJjNJ7
ANPb50z9jEOSI33wXl2fRoK3LXSjUTj+fPDv32u6cvUSoAqrrfefxL1Bjw4gHFhEcZkujylzQKBK
7ZsphQ7/74ZLagQDGfGkzOlFVLQ2pfKvK0sEyHKuhTaaMOLXNSg9fiId5GDfotl2EjFFAEbXsza3
rC6eRHYPoYB2Pj4ZVHirtuzj/8J+rsA+Y7I8aFdjg0fHel77hG3O8nFTWrcHCPpdIebnqNFU07po
2GD3sIoy8gYkSDtAZ/AXsxKbebxgK28zBaMM8FQ8xNFbWv4Gb2aRDs5gWWsk4DKdTJyU+VmEpOR2
CLszMeODKpRjvsuMDYSi478hLmYAFfnbHaCiIx0Wr5PCQ83GPy3pSjspHzLdyfZEYlVzzZNJmnRS
cKlCE0lEFr3KKWLBxqGSOdqDqrlXSD3ibbIhV3xWSdgWOkz9xWqLEKDvTzcy7naDXHY+qE+SvGmb
FkPANFQXvsPTrG/D1HwirBwDVLJZlCV0XaQv89Cm/5K0ZWWlf0WBVfEHRfsCVWqqKZSla/Doa6/D
ghLNcaEZjPPLA9pUFB5YAexjmH0+UyPyBJsPOFg8kalxQX77nOztx51jGRdLAo7MXplbcZayZvK5
UBCfuilxDShnR88nED5PPbouMfYv77bggNn1VqnNz7/kfAonOgyisPMEnyIWvU6vS29Hu6g0o5v/
QBun0xlcUQekatTZnIuRX7JXEb0fHjkcc+8wcHYbP/112QXFI98MDcihvqEM1YQOahW4QMZK3T38
pDp/Z+et41YiXaa5SBPbOd7J/j6gFhn5Oakg1bt9A8otfT+SVUX0CUpLxlVgiojib/PPuNAJ1tCZ
G+hKhS+sbp+DY1rhlokDrPfu23jXI1XYZM36QC2PllOh1daBHW51/1ann+5rUbXlan+b2bhEnJZt
9J4Am2CkIZuvcNdko1VDQsK9l+OV7qowe7BpbY6+nypU0/kGqqcy5jN3wbmDZs4k8JB3EatYNBCT
IzRPIxnePToMq08cXny2CcEmZsZLGzqjVOJSoXlVAFwO1FN0EgDxFna4HQasImFybIEUZfPKV9jC
21zP/UGWyLoE4Wini2+NqTQPZFG5gHYLEixQoD5wmZuMZDwHq0QuCvYCdP975y0NuRiHxOlkDN2n
AGimQK+WFkIYKxqyOt8SNUpQNAPpYIgNL1ijfvShIdeu0ZKsdqZYPxZ0VTkKr0cwtNV/E15ml9+B
9/bmx1k8e7BU5tJ58yL7qW4aN9JAUC1a5O/Ru7iZkgxTtJ8xL727Ih2IdQlFsqdwuas/j1zzVPxW
UicZV+0HuRDSs2nNQeJM6s3dpk79yWk9xrmgkCE40/NK2J5AOz5fcoCMOgPjs3lNJ+eLKFgVOm1r
f15FPWchsUPE2VbtPrqOOEeYa27PoPy6EHQrP9lVkChMFvDgQ34QTpBC8YCf7nR6+MHij0jaNIqh
JrcykvTf+vAW2u+upNAx5N9PckWoANn5jCBfAKwhGLL96wktI3pV7E2JRIy3VgfdNYx+HOvz6yhc
3wiqW0ZMi/Y37mE8FqlLB31PF0iHeTO9bd0lrvWqXNHYAfw9aUXAyEqA34UeI+Z8LUSeS4radfgT
EeSYz2m640+YULZyQYFsTSJCWlSdZFRY9jA7QcNytwEAQzaZbvjSE+3gqSnRF/yJWjAHRgioBAIP
plHKQvPP55/+FAsbZDM87CsnU1W8ZiYSPrPDLlZ+8aPT7DooglG5E+wi/H6SOdrp7LYMSItE/uUq
eLxid1tzZMp7SPcNV2bKINOqaS9w6wAB2P5XPM/g9CfuKJUf8OXEeso9NxEiP2dEwVshoXZ6n9Op
bd+4oOoPX5VTJpDZ5GGYgYujWBRNFW09OD6xooNACbTCheoFDkwnAC00wwm6NM9QL38NANF9JXAN
R8aYbwBFnSwNeAgk2iH+ZVhUIx7D9Z9B/B73041wk65cXtfXg42xFcjwCbRWofZt7R51wGSYdhNS
TuEPzV/d+kIRHPukLQY9BgSPahejSvoHwPAQDhj+9y85tvJkbuefphTb2NaQjW9WT6sSm/sWpM4Y
9QDTBZnrh4JBi7ySWzUygauc3Lt4veuCHGh9V7kpi2qZDk7Qd8nXBYfk5k6btSZ7SSDGqAxis2vG
DnmYyi8GjiYEpAXRqaL03DjYVu2smCRchcrh8l0pECwPwJbEK1AWCOfeh6819FIcfEG3ZFfEhm3w
MktrjkOpaGNnuDCnqolpVmK8sAdWiPUW3M9cYfeuWCdJcuoAMOZfD/ggoJdaEw6ct5g/wq0SfWni
+d0Haj+uf7/uwIInpxVLMnnJkuS37/20uObmGNGhKtesaLVJo/ffMpW6x/L0SRIPrjTU24J6/9Dy
xlqnKR9//mZxNzPtnaKVTG+d3OKOehquUOWqMTdmDMe9Qu2UmslKw+KrKaNyjQZQb9PBIzgmvbv3
qws/LgW0C0L1sDb1DsEhMZnnQw81Kn4Qa35SFyFb2yeZNWUDKWGam6Of0vBK/MUIyyTdJGmf0H5q
6ZImZ2mZrXDpZw7bW0gjCBPyfDuRQ6arvQrB/uHRpjlgu+MqsUBrs3uH7cr7c/utlNAIcJbjCsn4
6in3qUgAaSjyr0w7j0kNbDLqKlwrpF/2cly5pNRHiK4VFVyG6xCTbDDU+CVylgjHJ8mBBNRlD05Z
mJdgd6pVKiLOcThYbrsscyWbtrs9soQ8JIa/zjyEdKGKP1Msq9/HIMeOxmt+Yk6AVFEFugIEwQw9
sWMlgSSkheQb4JhJqaE6VRIURoiXhWJZ3u1dt7OvEfB1AceXrhqP4EEGiW1FCPh/MtihRWABzLX5
O3gGAMJGaTm6AfuxoxDFkASLR8PsXdPvAIYhgOTDQ2I7cZUgIdPlsxW2nn3eshN4XpJnDh+H9xOO
Xqs4HiQJPb+LbISp5JgtPAIuvrAdLFwSpJawN9aAMlkpxooNc8xadzPeACohokrk0hd7psSfgtqj
HJUy1ri0ypAz4il5tt9yPWO/sY2GEmV+7EW4qGzm2cqkQYUHh7lACmGXw5YPfhhz+IVPDaycKqDN
siHOIphV4g7O/8fjy0tdsaTkOqCGiQRpWhM9qEpMsefKV97Acl/zzaegxwwipVXWZ4y39OGy+xfD
iqv6Wv6YUXMIj9fNISYOq8tbh42e/q3J5vAVfVbHl1tUxn9qV8nUwH8qb4Won2X4evZX1N+knBCJ
m2j+vqCFZoIVGRZPDOvEhe/Z1xe08FhJox6fRqDmyObu/6BNZ8lY351jNlE+k5hAhia/KsuLED93
QsMhkm2v3hEC8JWi+qjHo3W8RzREkkmt/AUzFM5ZXbGt7AUfX4i8RozhvqJaBwWaqHfheJ7B9QHE
mNcRVUO7zqtHeREhR3abjA+3kuPNbpYHzOJveLMu3kar1oo9LAjoe7sAEcBwvIwtpj/jtrtGijLW
CQaeSzMcIohl60Jsoh7aL4tNvANBXP+SxqrJvSHgb3pKcvfbDILgL5Az0PCPg/EE0/V7Z1aKqI1J
ojplTEyKCo95hsuYShxPesqiM6pBDjY19rKoR1j0YitJbucb0eeDr71RCJt0X1VEA8nUk1ysYbU0
aMeYk2H7X/IOeRvQXpvF2RRg+jfzNFHmfkUhE30kaBtyKNidrLO1L7GoZDq84HhplSDgi9RNSW6A
c7yCwoPvUMXWclSGv8cmU/QDzHg6xLh+/JJzj7r72Yq+3zBriuLfcECDzY8B3f0XmghcGtfnoik+
PQya+4lxNpi8zS5AR3XIW+JVLX1ZWuxO8uEJg2JYxlHdACIj1Lid3Lffs/OB8Xxzo4tTpbvukY0+
Zu/BqZh7R3LOSCzV6wzsRDlVP2YR820aP2KHCBJnxVsBa9lMu6D1GrjzGoHtyfkYcYp2aGn56Qqh
T5u9YNkwJsN+zxYQ4Tonc3tDAVjbUepevsTPzeUIV3MmLz06BMXPJA0JX4l7UQKJGpCZc2CZIKJY
16RXzumGlGG0STkzcg58I5eeiRMdWHbq9GbR9vgFQeUQ4Grssr71EgpsYyO9rD3hUE1TU8FHWKD/
JCI3w2XqdxsHcj+96JuP08FbNCtDLxxNVyOUUAiwbPO9hmC8DvwEsF2Ka9XTr2tM1JnSDX2sGYfT
7RPQxp1W6wmyecxodEsgHh1C6SBlVAC6Pg07fR6Uu06O7RgAuPwF2TcugYQjxpa/biHjvzTbgfhq
UkG7ZoHVTM7St3KvOBUatfoAFC85Rx/80mtVkTVNILlIU6/8jgSeB+tMaQO3CG0Gh0CzzT2ZM7ac
i9JW7eYcl68ov2bw/qQSs0GBp4yGc2ITaUL6I78x6Al/+FdHrSoAKJByeRQcY88TIzWGU3jM5BVT
QX8B6FA76Q69mjBmGshqKc3/PfwE+2/ndr9spcGoUmObPD2qkysL6o9+bNKTM8mbFhD5Qja2DFhu
FZMN5C9pF3T+7N2UHJkVT0qs5SAh+q6SbmtuFQ1H5aJ66jhq5Bd7TfTnl9XdIYTuvAXbZK0ccmqA
rTO2cFD5Vt86VIgZvxKuRvwFoFFShJoiFGNm680xk4VW9W1mnP+2Dn6KtwQvAIaOphqSTY06oyv2
SaRV3EV7Y6/0tBPvbhyU8KLLy1BEJWeNyeFgjPvvM+02y8JyNSXs6495keFddfQJ34quLObLUHVb
5PnCI7Ch/PvDdEStpLnz8YbiiCdD3X7c7Y6ww2sOrCy+xFPUg9tR060AJ5PZuPpDjvEifTM4SVg+
NH5fJptDti+OgMMiQrJl4gUnvzfrYIToFjEk3yrLJ6zo5wCYCmkHt9EgTrwLxF1LivZRsAknQtFc
AMaFw7deXog1dUrG8j1xLrLkNRbj6g2X+8eS40xCrSF+AV+Wf0omPAxUwlllQHIWVZlNcDWjEiV+
+p1Qns+z1uoi7Dx4fXkEf+b+K5Z+KR6veCqCHR0o/iCgmNJVDeq9fBgMHszbdy6/zNKx4qevefgs
3++140Z21nb1fEX6LFMmYGRGady/CE6CmEGMcGiC9q4JWH6sfre+68IY0c2Aveuue413PrejEwmR
eE9AJpK/VK5kANk2iiOmnvzS+v+y37/Mo6gHifo/u1c5gQE4cVhIg0BxX1caWSlzDGXn/UHRQ2eC
kLbduzesJ7HnXElgQ+snIdBed7uG8fF8j70arKAAEDF54biXSuULVzsrTIXaXI8Gksc0+eyLf5VI
EIq99fDj2LvkjxIpfH14EH3ILOpvaX6x3mR5pwi927ahgnTt7avK+Jeib0TIx8B9NB9lId1BEzvH
5qHD1le+ngGoCKDQ0GHu/zERhzR+oQxIgo9txdFR5qI6VHVmYwA+xvW+Q9CzRltKxnMZhwg6SG2U
gvMumEiyAIbu1ns0Shf55h5dFex3p3obZ/0gmhwRwSUaCq3RvAreWFyuAKJwzD72DAQhCTZtyN4f
WeJsOD8xlcIGDaN5HWI1wDHm4orOlwVS3XRI8Y9Y6c6n6ySSQhPcptCui+NHjFTKpODeBw0M3gdL
2iMXvpcP/A6uD6F+uE/r23uZKu7clJO74Gkd0+Mxg9d11ObNsd/MAI8FRHteuBfgJspEPjZY2l4t
1LkH4IZ00Y1WHJnUj66jesQapp+8uR2MDOvUHEE+ukI5F+QaDzskH8U5Tdnh+N6vEvyk0WbChIS3
m/cVBEApj1LE0QmllPoT0GWEo4SwzydCpGKvLc6G3Mgm6a3w6jVQdMsNvCwRuoxKkItQzB3suCZR
pH9wKKzROOsH6f2UpCejWIMxUlAPpzCiVslrWtdNFwBcsz+OqEEAnl82FPRONfVKfKQqrxjjielv
jl57Srt7X0OJ6jA2yhh3j7Owj+UoFiMgaouYMaX0vlzKgnXapTuyyChgKEptAcLG1QU2WDr6YU39
1U6luzuRqWtd7LhsD8/ycp6/tB0PYhXUoDHuxxgUXJzmX0nPyBHLYH0pJqa+lXRq/pPIL6xrl62y
Rdt1J6ZduUH8PoCWNhlVxdsuwOSG4vDqrnUW5RVbz9UM1fqbhMfhcYMfVjLcl34BjgG5bUea7Giz
e1RvjU3xB7P7SmQqx2u31bJtMdi309pis7m/wDOKbtdgjdaqXGyARZLP1DGwabwzmprWGw8uF/y7
fh4btxClx8ijs67bKvgRRhhhJATBy+pgD+QosAM8AotmRMamdVNUdKY1TcuqZ+Z+NyRQaW0/eZX4
WMmgHX0AYT9g//cvLesxxOlVdIXumtYoDBrCLQ2/E8lhpNhVSWzVi88YQAmLrl26Q8NgHpAdbsKV
5FYQmsFzjMVm90qqcanJKRKQZJnPfvionxf2EgWnhiq+BJmGMUn0EE7RkpB2PouFGjmstTYjyKnI
kUL1onrXgYSNPhed0dpt0G9QMw1BYAJSRN5AOKXq4JNkpjAkTYG0MTBZD5KOXfbR4Mp2XxQ3SkGl
b+dAk4WuXisbBo4I2WLP3ana4amwKWttwh9ySDYGCMvPSUo6tsQE0zNNG4j+SlpBuDJtfm95MFqi
i0TZWtrOh+GOIRAv/vBRpy//dSpBzETrKfpd+AfW42jW7VaRFwdMVYK9V55lbwcaYpZDM9uRzbwI
LsyfH0kO+VYOuaQeUt6citI12ykclGSzHZ5Y0G35rnezllXMrlBxu18le7dg4fnhL+VvQ6AnQ2C2
7Q2qTlmPwzEhaiIWOn1bF5EG+G3UoEAjZOrt1BSyUXWf7iAkYnco0EihJocTVdnyXW+yMaJcmYMz
KR8hGScmqOyINM9GRofZ2jespWJN4BId6vGZWscNdxFjM7AJKAjuqYTzkegeFmgeN/+aL/Cin+7x
d2fnBPFVuEk2T4LywgpvyKI2dG1SSwvmLR5tCVG8rsKaviwNT8UuZvRO+N+kzD8C5kbKnXzywJUJ
JnQ2qoi9pXtLBXF5zTPAcas1U0T4XX7q8vyZagiGnuhhsZVCTkBHJXcZdb/FvXv6filB4hhbhR5t
/kuwUlpQHclvkXfEtdgmOZ0q2Rj73Z6ie4LYlKW/P11WPxDwwBMj6IbW18WvzgJP3zUhu7L7qWv6
Kvg2Tw/E96e54/I4ZETkcYTCZlM5CYNoEzlXTNu4KTBHeQlD6nK0Tt1j1hNFSngawPBf8h+YMAHz
z5r1c8FTRmvFY2Ey5TEjaBnijTvxoPSSc/DVcUWsnOn2QPu+A+ZCKqLGXNSKhVpSFAAQ4CBqpdnB
Kmovg63onYj6tNnaqqDj9y6g1wcdeIQPG9ZqkWZf/+Wz0igqBDqKomTEefPXpsVl8eoXQKfTi3gE
TepLKPbLzeHBhFM0RZf3BuVvxHbEYZeG3Sf14mWCwCWQ2N5oOujuN3eXdZTXDpM5+2EJZ5thQvef
k4OyFmEee2XzLs1NZXubIN9bK+j6EP3EoHYJB5xTvSr4XZaZJXUMAiLUBlD64JpirJ5CVpAxMJmp
hv+8uUIK8l1b7hjELs4T9O0DK5GPkG6cIXbOYKWdo9vwRG6djp1qT3wE6yMrYjeoLm3QDDBxSGgP
vbWiqK6TnwrEMLMQsSdsSRbY/kcqNhLIxOnsHhcNAA+ydAVvzlpVLvjbhGUU7N/hWhK49RW5ahy+
Cc8tjzfbVHMy7eZXPRey42aEDhlSCEq9Xrni6VnW5dcR+/GLOtqNh3UdE/T6A7vA7Zqvj3Ta13gA
m7h1HX/PvXQrWGF8l1ibx+mTFk74FgHrM3yvT01OjLLj1yyfshnMVdz6pdG/gAV8Te+mtlM569xK
ui64Cux7Q5NHX1aT40EO0zOgcWmVNRYkvMEDt1FUTieIDegI2hUwAOprxrkbNgb8ac0dQ/Jpt70E
cElaoEcH8v6k62DqAh4FgNtKhCbsiB17jdum5k8DnTzcKoCLJTNPXBs5ieM4eZHGnRtUl5RVTYCz
AYnpkaJ6KrHz1mxPxON8mdUaJ1zh8VWRK5O5OC0lgKSxmVi0SkndYFmi0NzxLNjijgjamm8+RtQM
H1K1PHjIibK8l7//0kVl71WLmR3ruNMpwtg92Q49wZFm8q9vRnqZPAX2zxK9+/o33hdURzCxw4AZ
HN+p9i1ER1/+0/evvIpRejw2kRwGxutNeaxhYsWJPrtcI9yUj9fBry9M7Y+cVh7bSsOsx4Go6uS8
JbNIhmgwIjAlCqa+PPqu1yNcOL4M6o+pMavqtl4Uka2lku9BbzhBIpajmS1IZl5RkgmCWCBLiCQk
LkxUCOYpwxkRypKPMXUxr21q7qhRO/zLhCJLCudLqM4R2oI1KDCvF+9QD8pcwRS7/AEauC49Qt3w
HwkYeKp6O9bAa11j8vNy+38t7KjZBgKXDaREuuf0qmh2t9u4s95ef32lJ2r/ASs5dZrC7vX/w6N5
jmTWPHgapnhs0Fq1wYUqaOeGK4uQKGmCjYlYW7TBE1o31zRXsbWZZ35y/IRol/a++axlvaWk7Ou1
5MabZAYirP4Itd1HcyTKOSF/Pu6+4KJHp7xuLDBufNt7t/vDN7lHvUvvxrbArs33pM/p9+5KEOuy
5uHVgH0xo8btQqcc1Pq72fLP/WkJ6l4L1dHNGhdwpRV3zw/eZ8jOS8rXiO3h3WU+Npo+NC2fW/yV
DLOQhCn6/5jrxfsDCAXNCMabDkQPLhdnebegCbTN3lS9Q9jhJTFwxtHrmoGI5YDAXy/kYQqeGtg1
wPsjy1i+WBfgUZthw/TvdHU0jaKbd5vG3r0OAXCYX/31iQBpn9qWe6G3ggdBPqCtFV2d6aesSDRO
yGne/Z+tCOZUWQKieCjwTTYDvnupotkStBydcE6FMQQDvQxc7IqrobMzoEfu5jOuTaMCbHfRQkKQ
b+/i2WUqdH0mThDvHpGlDQmrYJMWIT92kIKpbEuFtf6Qh43ETwHGcuoVtF/C3RgqfH9C89hkvLbD
hV5o4WZ+uVSt5xChhKD/lys2SJXU1KI8ER5h+QReqHQdo19eF5nIsPwfVa0XNcW/aQeYMF14XNUZ
KcePZAyq7TMHAgw/tuZd/HLD/OFjsLsp1gVXBnIxkhQlsO9f4egDQKHOXw9tQz7TDu0GyX9i9KXs
ZcQpwRCQNjrz2TVyZoZ0VAfhZEse4pTZLeUbszxY6bwH3vo5NarlGukX+GCO8pmQm05KFGm5NFb4
LMxzF1PmmhX8nif9rQBdGVsrDqB08RuH3G8dw88ERkV783rL0rgfIQnljw9mf9YU+si+HVtfHJHf
M84KJyGXwMjR230Bzq4MPhncUnkm6T4FjQ2EkliQ9B6HDi3ak/KIj0vFHVXswyH4yNZmOJ2ZZ3uA
Bq27SiSpTMvd1zm+pFEFSac3Gl/gdvAqMvbbc2Qt8dtdAj3wjkTzXIXVWjp5H3hc6oIrHvKRK58t
GBC6GM245vm0E8GmAXexbokr2kkeXs3D+4+wZPov87Ogn9wm7rJqzO6MLlWORmYAZRdBPiyeT1VJ
xsFRffb56+SucArWpwGiudLIFO0nMnWqw95svBZ3TNtTJcmwJN7EHSNy+qbit/A9PUPFTfad3BnM
p0a6kCOTOZ5KhufbTwTZHiYyp9LQi9VJ5EgZfg2+D79iJBx+mm3esm8mQyXk/e1cZdvduTrWBm0z
52CZgvU0RqfxaOSOfPaAe0505eKZNZtPRFT9fNt/HDT69XDtl1P6NE/osB+pMoTHREQLfbeq+qQ1
HE2Pwvkxs8cVRno9CNEfbOppQRQ3n+Nl/AwjceGbNfSZeKv3/xjqEB2gDjoHzmVfuELkuSFfimMF
Ul0hRJLB6/rQm8ZGO18wx1W5Xl98xA1oUjpH/QlyCqQayZAuzu6vHXX+EYGOeV5eX5sAwEAaN4jr
a1yUIaXYnpaTgVUh54OWOCrWsHhNusGAFjarY14927hinpZZCyZGfbUlCM9YieONH69z2d/w/mS3
2qVuAatiPM1qkOY8NcP58/DrpnEICQVMymai5d9eyxaF1i9IpaY+KSxFdtkk8+JY3meZWaJvaC+w
Xxdu+7ifNfc4JgPP4FpCjWhiuKyhg5x1iDbAJt1aGLFLdL4FI3x6r+RtDsFeXmaxsDHDI5rR4xdB
Kz7MQYC8xOrq/O84u/l2tlI0uKy321pxrswq6MbSPVzuCVWUZkAKXI9bU0ReppbaPULuMv+6wyiT
4Z0yfLVxoJzn/rDpcr/kl56EUvQFDzZDvyiSPa3KCRgW/CO1yiIDO1dsz1a2i1xVK//Y1EAzjZoI
qMIkb3vw0DhXm2g1DokiR3AIw1Wvu1o3ruAMw6Xu7ae2iVhPkSp+vcJK+ZeHNlWaw7Evj/uTTZQs
cBSdXS3x6elEkoMfWSiPhwH29SfLGqfqqJRoLIjw3g8K/x17apcWfXcUj4DWE5k1bApUhd+Klt8h
bvCSeMS5AGbsaThhJo46srpmYxF8As6L2wwiwwaSUys1mYn2kWFKb0V/bGS10/hgHuOviHpkmOG7
hl6TDDZfUNU9k2iufhmgGNqjJCBA0bKabZN4m37pBhqEdXmaalM4/eztoEqIiPVLKl8kg2pQ3x7g
Sab7isFVcJy+axlP/ER00/dy+HjqNg9sbwchDYGuxySQHnioeJiWcSm8ExMQjMp0CZuV+JzgZVBq
EkYx/7Kq/rFrfuI46eT0H1GOiU4MfR0tLNNWd6IYovS/GNcJtglPsVimhPfqv5C/VxmxDgNlXPbN
qkAsAOrICIfX0kMf2RUxrJOBEMFqDr8vgx8NuuH6FOCcHmI5TWY/roNacvD6ukwG30F33lqLRERK
cz9kOutpjqitGxv2vsd2vsUcVrUVhm438tz30iURRXYW3qKDw7Zx0E+7DxbqDldbaRw+kDRnLSby
1j3Y/OZLhBEb6XpuIFxuoqaWZ76fLQ7W4cG69P+lQkPfj02csIwP2iZmIdZ3NfwFAfe2mBF0flqZ
Or/euwgx5sJFmVmCSY4Ire5ZdRu2tLRHc1jzkhEXbCWamwnNejBc0HWt5cl1ewco1koNxpqORaIU
zCSRn/DqeMJJAr/8/hFPNlssJY4N9/WB52kkYL5nOhNPqUsR52f2WB/n82CvSvYSbILY8sMhY2NJ
rJczvGTHLUIruLOp7XycgnyRsO9FoKtTbEflX9ixRqtExnahQQBtpegG6/1FgkLhIKzlVPE75wl1
jiMCd9g6qlFEZUcUqCKlJE0J6lUhVyFrb1eN/sZd49wUzc2HnhE1QCmGJIwajyQvot9XByj7MuS1
cj5NBvhEaK3BQV5xbJV52qFeTlDM18pNQReEBqKuKarFa2dcHwZgdVd5C9M22XEeahGw72nQ6CZI
mf4z6r6r3ZCZEXfAS7F4tmLuF743FWlb4FsS4Ohc9OL9Gkq3e2U9oPf3GPSb3MBp2ayW5c1TTeTN
EsolAgJ6vmi7rQXE2TxsAEqWAoacSjDhvsCeb8pH93NVFrzk0A1/YMEUoYqXQHOCYZpsI2VWM+ZG
Ga2z9ajKhFh/qPAl9B1KFnlx3sQJ0ezA6n6gJaxqxSGfAO03UjMFHdCqPUzxmjJaa96UeERq5wfG
IcWCgpPXSCa8pp17fiLXcS9kZO/lu2/SHZTSd4HJMtj6TSZexX8JAKUJITr006/8pQqiNxZfXQag
U/PPwofN2F7DdDSelUuWIvTjT2/LmZo67NZc12GT7DRnHvDqvdPdQ0FnZeFb1gjk9X+uOsrsq/gs
Hm5VJWvG/fJRJenRakxpai7/MHp9HrGr+jYsdENeT00Abhqw2drNprAqz3f4ySYFuOEpAtDnYTR/
Ft5NASxPLxMdrdl14Jn5131BDyK3o+EKR+OupZZlqE2zccPWIxgUwCib0RjO3WHTp7uJbi5jvOT5
h3/q1+gzMd9nwQ1mfCiETliiZlMbDi9//u0HIMGeSFi/w9H8Q2xQ/YOd/QbXxDw/lfdsappf9k88
UrFJ0uOvCKrQ6OWzHq0d4DgrSNpOX2TErzxdjtojyv++i7C93F84/6lWGqWPJyRZLfHL5phwdWSu
EKY6ZyQ7elzgeB+dIbfeUe+BdRYQmJqwi8RRAShMjPpVtCwkDrzGOButfaufAybtKPQjshzBnAX5
AtZsCvG0CM9l2zZtZSgHQOfpf2Hg7+r5FxLq0mWAhj0Aj+aKzMDPRDKUKIauHyNVzXmFtwMZcMis
BbCElvHg/NyC3sOoh+N7LEn7/UVdg2lDZSKJcRhVPFHn4QXfoluR1zjEJpzqT2bTp0yEltT/p4ad
Ox4GhPkrXgWqLdetNXSShtkiK7FMPPnGADMV+nNg4yIYaKqKbTVBG11+H0RqOQWuVPssZQ2VM9IT
yAd0YhlnbkjPBLmiZGWaWchEfgtMwBiuCZSV5PziNtlzjcZ2C/qhQZk/WmoQWf5dk2WpUEKtBDzv
c1BpWndSOlnfx8RQTTIrRSRI9jlV3y/zkmUjVGHuuGAIjzAYLJrRqeNa355hi4vaTuIXrIHFu+qn
DFRdi2seNb7cvt0bsgA5rcF2L/c4nNPRMHf9LFHNMe/LIMEtlTI5R16C9mq/i8U2u6hH2XeW5Pbl
AgQ1IaflPvWmhjeTcrNDRzf7qUhMCuh7VpneYw5w2UmyvCMc0mJGjKdwQvtime2OWcXx7UtZ4mca
++feR+MCteFihJHknCzFsFiUDj65dPP3cuCCF+8HYFUlyy7r3MyE8V9RSCvgRkfOZO6//M6eJ4JP
PzN/XJRqIMsLwE0KRj3ClNyOKmDhwTf1pruhbDB3OOvYB52qFNBku8TuwXo0PGwVm9YSlSL2U0S4
sZ7WRa/SzG4r7D2WCbT6RmY9aUuVVEHJ7AXhR116CSHQICn4GXt1kHmHQ9/mmGWtPyRHn1rv3S3B
VxO7hAFfB0ktqavd/x/KfCithWSz98K2uM6eZ+xIcYdLpFrkG35W0HNAzJlciwDDK942jSA/jjsO
xEnnPrDYNG5LIumLO2GkQLHk/PdU1CyCfLsoEx/P+gAJyoPj64rjdbSanSIm12tOZcJGJDgJGX1C
andYpljCTARGOOQnAeyoSm4oe0iJ0+PCqJd0MtZtAIEcfAsBntUXZYiqwxn95r09gRJ1Z9Hx7DeU
xIB6DMqmcyf7M7hA+tcc/bCostPrLCqsF8/toqdeXnQ0yWmPu7e1DJMO9fTlZR0Mge9KfTo5hD1K
P9N5xxUSZfqX5fqebH8LBQol6VCKjFLuafy5GPK4hpwlcqL2L3dDCkGAJlLOT86cni9PTukNyqbK
HjshR/mi5VYj3fc5tSaru8NvLzCd2AjGQt5+4sCFcwwPEWkA/D+qaYsTUL0wUTj7zpJBsBKUmTSB
u4quvtZ6yY3EpXdsWyTa90u6FGzaCQ6Mn6JOuIDjQza9EqaRe+gJSLjL36j+jMvU5LBSoj86a7QY
0Cm0Cp8/OZ0IiKLC5qYstc/1g0uEzAp7Vc2zY/8zQoUsigUjv72Ha85qQn2KqPe820qy5eXg/nGc
aJhH/0lLrdB7QYxLEe+qwRAvk1bZTSJS7cZ5FsS79e/mcBQH1LqWR0mtWd6oPEvcpNW2wKQe2KAB
3BjMMdFvmL6UTI2iHoIy3jOb3LIGn2CpoSQRHCtZJ8VXKu+bMuCISDhTIynkVEIafKI1GROl5Z4h
Q3zIRIXMwcREy8d77Iqj6csY5J7dpL4oZQfsrq8D1BrZvSMVYhhpJOu5Q7zvpKWNNoS12wqNZ7ks
4KUKRwbZi7ms7htFe8aCIrPUyWvM84DVrto60HB/qsbtWDPfwnuZ4IWJYh5XB/QBFsM1fcyhGmbz
kk+AEGvSw0wNgzJLZpYBV2mQ05kDE607FZm0w3NPI+fRcfJfFQtFDfl3MokpD56RmFFiJskhDWzV
bPbifJnk1saMmER5oRrrriofD6oAGNn5Xo09Yf6nLUAWMluE04h0FC/KMwFsPec7Tx6kncwJWZ0k
bWb6nKjfUOg1GqcnQy2kz0W/rVoZk3Gfv81e+X7ZJXPC4p5eRwfMxn0BZl2vIm4L1SCz4zX8swoE
0+OjRiU9MihZ8r8aVY/CRaf+AXJMBgwym/A1HuhzQxB91HSlmTu308nfY5JkHXBTzfDoCtvni+11
Q7cBB/ZrSy4Z2TuDYKRjL02n7Tvh4v+Y6tshMJjFYEp5aSR26duGZIOUbx8hZAp6LYJBpiRD+jhB
43W5zS5IDi9CXQz88xTHWLpLbC6o/BxwgHFnI4ts+GnsE+JVCWNhHjKKjnpcCb1tiM08lYEMA3K3
QdgvTT74cPN645zJ5QhNUbIAPlkKeb2ziZyvyjlsGJEmxIULmYQnUWACDFuc88j+z46XGJ9eKBv/
hiXN3Wdf6Jfy/ekaZCbE/Ru7R/O+h3exuSQ720jLN5/nbpybW+q2j/IKoLtoNKpP7UgXYsPPe3X2
wqmvTW0Hh0jm+sGEmc22qQAchynwHmTcqi2tDy/jN0rgy9N7xUo8YMOGDmfc60W+gHT9Ab/K69Ku
eAspVVjnEku0EcLunS9LxzDwO1Hrd2qJQiQLH/SlYSr7ZKQxgJD4BVpOTHZpu1mhRbwplk5JBiId
3qpFULwxqec5Le8MIq9wr7aAkdBA1cWZozIBbe5s0HE6kvhv1yor2mGmlRoSMJMK6SAfrQHiGUOY
SmtSOhtgwKNvq3fqAVacdf9vagQJU6kWzbcT5/qo3P08VEAewIrUH73sStGYRkNCmqpl4EcuYq+w
9ULt7kVdogIm2Gv4BMIytMC3cUB2zPptn0Q2P+RS8E+WO1Y+OahuWsRtMYRtu0QxS8DCk1d2gnT5
KV5/JPrkZ6ouJAnA7n3cSIQbmxRckBOce6Cr3vuxTboYSXrZLqCr+OO9/ENtZURIOnh2tyXPQwMO
ccjGEYPcXAsRN/8u2Uut2p/+3CCAxxs7LMNXv6dK0HbyMXL8rmRJPHdQxy6wvvxYXfPHClEgSfTS
RaOcn97jfh8+YrR16poShz8JvVt4hKcwhENqfgpuMIcATEGmLuVYAP8ZASGhEWCVxfdjz2h+qBrr
HTkzQXcxQV++CtoDl54asM4nE3e3fZrwFZmQ/SF5Un+RzN3I4b/XANyQL+8uC0YXygTY26Jko47A
jyRUtgdRGfmseNHm6KTc1vzxR5/7pNDeP0pnLuqhYGxTs+tq6zT64Zsk/b0zgqlC31o7l+icAVOm
AsnFOtKrgfY598psQyWYDafN2dzY7tU5oTxUAXorcEtp6oWOIRRts4P6YJnFlc5d0i/jVfqOr9QV
YPlrK12hbmpc35VQxY4SNENrbtzZ9IWdrOnwcO1a2lVgOXOmcWGAxHMP0WrzvmnUKEoMjjU7VCJM
yffh21F6hkcYjwOatdXscTKCYu6l6jEw3+yqj3V5TGXHBQ9IqnSaSjM9mJXulmSkwUMwELeIW/Hw
E8I7evaCTOWhzR93DzpWRXVo1kDSTuMwrlHybavsJyxewuiCfNb1cAJRFdErrdkyaBXk1YblJN6i
zUN1G0qXEeE6CtynAyp//prVfhhTZyPKGcKnPFHYd0f9TQHAQhbLxQH50F8dkRLSET68phE2leqS
nncU5RPsRxtinrAOBTkoBBrMEW5zgmg0hwqE10I/t6t1VtSeFaUw+XEa6wMtOOrvJ+V1MFtIgR1K
oze69kDx4wyUEyENG3FkUPoUVD9InHbyBWU7rKND3NNBSeM8fDp/VPY24+dfP6+5s1Xvf60yt7D6
vzRR1mEaO0oaoojOP0fvYX1Oc+6mDvBjasb5sUfqcpNSBeuWHAt6gW2IWlOUXsGHV/BA3O0ANSwf
+ZWT3oCBLisZ5NhW+ojbut6jPq2ypvTQREGaFMYBniAsgp649xFAI7vsMupH06d8atsNGugysN6D
n93QjYX1sZYw7MVYkfs4JCJ4MCpFGsP7NC31WyGUOVDcZoa2Ys88r+l8N38FnDf+PTohYVFkZmYi
FmCMWzrCOuG02I0vlHs/LfNKlNjYHLqhQbuiaVgsj84wnkT6fnMmmOeD1KQUCrPXg5iEqfb/wV6R
7kvvOefMjYHCVTcctemwjxM2IIFaZk1NbSGFjIfelunqf1r+4DdKE9alcaPqzV6hlbLzR6xUiXkI
IEk+Dgy7weCELLILrNwg0AkWKtyCS5Az8FaHb8ynFn48jNSukY3gdvSumuX3Np3aEyDxS/8WUm2p
tcVeftJHrx0hBzxI7/LXdaQ2b5VLAxS1wkmLSKspP12czwRXVjcjkHWg9WFFiNFXEsG3IYM9S+Qb
E7eUM0Vjs65tDqCHijhJKCdXmU9NiwGoo2aAhf4j+ZcpJcxGI7IvoSKfrIIuhQgHFX78e/4JgRTF
G/eyMjAZmJksvG6Tys+s3DWydGHdxjqE3OR43LPaNlX6NJZiDx3JXBpPDj7Og0Zvf99ezlppmp59
ghIpWfi5yAkdpVYgK4oBERbd+qw2gTbcsAUbEP/iFmEwnnrINESYQhg6un2Kdkse+ho4oF4qu+vK
uGl118vDAgXeGaUZ2d1F2qfjWzKtjxi1imd60hJy8NTOYUV3QxCN8c0tKn566wRvKw24UQHkdIt2
gJq/FJlQx3Ak8mC5PpxWGiYyAngpuOAS6RK+5ipSsjGaYFISMPdIVj4ZZEgsxvxwr53MYzS78bjf
LEYMwPfxYEjjkXiBikGTi2suVFW6Zl0Azlk4sZqvir2PbDpHMF79JsERSoJU1CgljurebSbQiFqN
JYH0QzQ3nul5aOJ3O5e4OmKSEazk5OzA5aHAz6b5smP0BJhHMQveByvvKcpuTaPb0esq5ix+O/i0
V6PX691+/VFMSisluwrLxwceX2tEIVtLP7QKwZmYJlxnHk5aydiHfQT3MJHNueQtsbZTRmCmWaHU
sKKFOudUWui/lzLudh+1MJtjWGKJkTgeDFBi2wKJYs06kyZFQz8BuLVXXhNnVSe2VyzHJuETVk9U
e8gDFCMHVlhro1r/rgfLS0RhP9dRHg+NTCkhBmxHHc4SLi6R703rMlGtv27x4C9A62rLb8WcTEhf
7csI6Qrni0ncjw4LjBG/I0tNrL05jU7+zQD4wQ9pwBUvf4mwXsqBD88/ZuYo6SZXd55mkD8avg69
C7/3kiz0g2elyto9SQZdcrGbIM6ehFt/0PBPc5Ir5lpDvAQ3BX52WaKp/MWm877uU4UE730j5CjR
cS2RC6EdaDYBASOqaWLJyoM3Wbn71F0cF+OQm6lIo0aOYCzFZOU/yWxnJPi5jH9Pax/wQCBiXCDM
4N8dXOOrXZmEw5EjLXeOi4C29Klb8UmbdkJmsIyO+pSOqRFON2frxP0LzcTNxI00YpI6ozx3gEvl
DSs50kfpkC861HoUS/S43cXDiIdJO1YzTc2ZjY+xNkg3OYxL5jpgyNeCgqxLEMdImG7ICH3CrLJ8
MGBHd/yr87mNyqzJqvN18D1QRxL+Fzhs0LKsNe4LQeELKGd2eS5dhBtv3Hnf1qvKzi4xZZChIVgm
HN6Gg+NQwF5EIolDYMkNae6mwVZlewHtt/FQshgmryCvbfST4UnAJ0l2KinU8Ewx7q7s3H696u3U
nU8dQK5Xe6A4IPlXVprtFRQg8qhMEngC3unMUbQXU8Cqa9ywxtOQt3twgzGmkTY/obhsfBXRVwcU
OOAp3E1tdECaamlUV/tM4vA/LaTrG/Z3lSMZrJSc8GEuAv+Nspw1HVHxY0rPbcK4CaIXjUSOtDwh
s2boTEiThZECQhLvXZxNHXpnRcbIVKC2a4PcjHyHdzP1hgPjshfxTdMRqtiwB2s6DdOsbwq8qr3g
cl9WYjpSTBUIIEua+raVNiyB+bM3f3N21Zj9SYcnEJfroCaXF6pJbxs2kpXtCXCfa1lN9w8OTA6v
9roOSKCqXwy13zD+EiSmS+3D91jwyERppE/KBBZLRqucLtFFyZlJhxbF0bcce9am1RdXSK4B1p/p
tLznjAvMkUboy4Gakj7mAT3wGEvjNX8QirT4krlR7QTpxszQCxgnvmEOe3FNi3nGATHzib3Z4Y3e
K+1lKlH4T3CaHbpA6N+08pWeiNpSWFyNZ6SRtTpwacq23vG/i5jHWCMRjnwvo7Zg7ZG8EhiqNIPU
pUHPNyhMGONjyNExUz+BfTD/URQVkR/UZBAbyQlvFpTXYP+OS/xIkZ9zR2UTAk+k91sBcCro146b
I/uqBWqsEBRmvkEZgZD2ILVrSi4DEBhhlQ8cA/APOEFTv+Um+OfSljq5J/r5RQXGBtnu7geGOCEx
Mhgp79Ztyd/6oKUyVLcZh4Tuud/m4VTxc5dRYqDaiMxjk6SyTNj5AGMcgFXRCauYOTj8yC6CyRZ1
BV03waPKT+DfCrf8QfacNiGSA1ICdJMitzB0ZiG6qSPTYTTujoSsWTeXQ7lKSFzkHEq7kGNJG5/D
24s3Lr613vsBuoIgnfsGEavZjTjKDRe+VZqsTT87cjGjVETDkaRV+D5BJsyuDVUJ3dntvBtMTSKP
BLNszKMdXPzVl1h9fXPMv49oXGvC8g/FIHA9xUXL1RTDzvzrH2sEKnBH3gkgzCwZyZ+OIny4a0lZ
EO88ErP7JkY6F8mtKXaagsd3k4pBAdD0xdblz4vvn+33CjKHVJB5O0v++sPBJtXvz3/MG11fv+O0
cRmcWebPnTQzkro2xQXv7NnXmYqMDAChY7+USbf02wE5HMeEV7rARJlMSbBOxZYzEyGDW30JCxU8
kfHOvKhbRRdTBAegvrQFmgCv89eQK/grfoNMlawxN7j2casXR5T2/9o3i7jQUU7qnMo5fh+n8MMN
A1NyRrp/Iflf3zGnaD6/uADVb++JNuBYJM8ECzxunB3d1DZNEnKp+u6wGkvBaM7xpO8gKnzc0c6Q
/MG/covteODMBNx/Kch3AvENfd2PI/HawNYXQGRFdV1a9CRin1METDFh/Eh/IeIGesBTFOsN9uEf
g6VJhWlrlaoeIaRHfsyhk7eMYgpkWN87hYM7z/DnJKBn2qbgoDYrR7/6OMnbsVhSlTES22UICA+D
NmsD+8BAt4qwkWuSOzf6Qcd3uqRcLjUiMeAIPtTriNJBQP8uyc/i7OFTvzvKL83bsMxbWP7d5LX/
iAVNsikkpDdhDmnauatyza4BmKtYMbU6rxTqm4AGtmnDyS5lT3H+tTSkGUcVZSf3PAFYKpGoltub
77RBiXQTRHAXlExd+hzIYX8xYdAWcfx0Rv2DLDJJEuZn+m1iLHYFAFALRAohisnOHQqbqq+Haq4w
EcyMbY4CYbwvqkCjXhXzX3mB5j7kZfvI2K+d+yd0ukHmMA7hBdfexbap41yoy4cs3yqvTNKfc0PU
Yfx8Dtr5z0EYpvrQ1kuQrPShyqV9nUgBbWPZOuBx0k4yMGhde93HAILleu7pMBlf/nKRFGO1SZ2j
WkrLs+ChGmvFEQGC43KeEfn9GLz3hosvoxFpHilkR2MeZO8Tj87ME5CUvL7mIuNLfLDz/4BP9+lo
+o322/gk+mI7BV2yWCmKThIkaz5wG9bCAY7RC+BPOMaABlwXrOUSCRCGxRVofasXM2YjAXun0V1I
WR96W/UBXgzweOc2Pch2BqrOtWp6T6JDrWlHx49WTKQkLbkOG5ykHcQxWiPYUKVMiR0bLSoIDbpu
TrWBKW1BYes9cDJ7GU/WsS6e8I09nFzkJp/cBXk2KJmhfPLVBZSHuNVVUicemQ+UVOlGh9yzdPiR
z69pwaTglrJZnFTQUBWmfs3bdrB9Js3VVxSPkBN+DpwVFKWdkL0oEkjIs/84QL9vvfofu04PMwaZ
v45/AIMc6mWfzJCDZ83vzti3OpnzzLnK+QJrl2zNaMVKEypbHltbVLoz5nkgPDU1rjh4iIWfqNFi
bo2EXyR3xp6EekqBslbPoAx/SQraHnn+HnWHWhzC8o0O+KkLpfxzK4ZN5FYJpjUT+60Zfv60zakv
iYDuW4K2XgV9WAkiTde4wsfI2zxEAOiDKOjJd/M4lWe7Dkz7ghRjzOKSgNjXmSBnyyhPFm0Q5d4L
AmwsO0GzsrcIl9yhxvtMO/nZ2xuNgSgquaVQJqHHO/yKbhtIx7o/iF4RO89aYrZLGlatqLn6iveK
kIZ9+XgTxHyEHrA4fRMDrvKZ+5vjJSz59BfJXRC9m8Z+nHuobtfNxvMcjdCR7C+xt8suEMBP5laV
EPDARphQj6cYnB5nLYLOWpQDOzhz2ymyKdhDL6O3mEJJO0QXQvVpRsdHVbEj6onmxPxDSw5BLyyg
zDM/6iJAvfq0YYs49LgOTecdDMg0U8qIDLJCc8qnRrzQvY7TgwqdMe7QV4VyLqe0g9xUDcs4FllT
XE1HxEzPJw+CK2ypaL8p1p75KXGdla6ScibySMvJPk+I12Z1kl9mQ1M4xiMIu2NSg0egkyFSQSEd
yy0Mntclu9HdXc5w7+mAiXa9Z4Sk/+t/ajOKThJq4tfkS2+DNF4QKb7GHMOtKaZvfHmDV8AeOIWo
Ey7/ezG9QL5u9JRECH1EMGS2VbAY/sJgAOE8/TFx0pi57z8RFRhBgfw3ryvPM03LxPI1TKIG2uU5
cUuABU6XwoeD9rOqLKCeogIjZzDi7O/PtgzaAyGc1mNUvo8LESmGmkpL9wI66l8LmeGahN6nb4De
YTZ2Ux1Mf65d7KgGO2IPbnNfpzrgR2mjjunz8ZCCqryxAr+8GWsd4QQ5yzFMRbDqmz1vu5xaMdxB
Htkw+gWS95XEEZf47AiEcWhZCxesyViLmiCKpX0wNbC74+2/XC5vKJCNDk93BD5tO6UrVzb7ti9c
tEiVnMwIZfgq1vRWv5IdtKpDny+s0Wqqt368akRZjK4CEqPY4GPhr8YxybEUplN/dPjY3sHkfWN0
hT0FnKsE1A+s6mdT86TjTAaA4Co0jNUaK5kxGhxvgSmnSb2iDnemruk29Xd8KItTwQ53+HcJYYNt
/vQBIiAoqwDfRidNtotkFaRXthbPCrqHwyH5exKVjSVfkBopOSU1xJnZ1w1Q+Zfn+6Lqv1W2ANrm
u8rx2eNjKk5bi5XiL76XH7yOhyKgwCeMu+bq4QSengmLiicHQfivHopzAHmkcKR38dYXVX/rWd22
ZY/xhvLjRN4zdze0gLOh7HiXakfn1pC9g8tIOmpte1Jtjn+hKr6WQ7gj8gOMGgvjdyyPwa7LTFJx
RQV8v+yRGLdDjmqEHXLhPzNLskx6gFTRatNyvC+zWvjOTo2dCQ8F1ZQzr+Y1KZJMGKIx92fs+wa6
cEAUjfVYB4YobP1ak6CP8RIxuLZFfZkQFQUfiB/0EeHiuSNcirusN0ft2dwphkfVcXmzpxH6zhgM
vXQEBBLrt1yMc5w59T3XIHWQg0DZsdrD7GhW4xuQkT5QsQqM4pZLhSUmGevSJHk2MNZBFoyeOKAQ
D5eZNwlIpXBNrEHKsehSQFhYchkCFSUP9TX4CclIlKTqbAyD8hcPskatHxZk3qJ2JQf71cahwjEU
+WVvHOa2zjv31Qwvl0rsZ1sV8ZYAso1n58xzbs46pKyGalY6Vc5AD4rklpG3f1FsFu4ftpI7LTzr
BKObi0C2uMScWfV4gDFi1JR0dQFmzS0rUzEZUo0g9sQflCBkws8Du0Bq9wWM4nEdYVXqfBJi39bQ
NdsKWCB4Z+7mUBGa7V7EkG+04j6Y8LuIVfaxILouc7L8WNzWbuzOzLJ+uYTiKLppgapCBJdbgNRi
sVgP6xY8kZczexkyXc9mD375raiW7TPpmLdKICRyV4RO7tHwsj2yFeV0ZXC+hUvGOo5IMFLzzKtw
/zpc0pcxt386vvRUySuCQHAsivj7YMH3Wch4NF+d7fMein4htrrkYCmtTUdbpL7RS/9dCHp1R9eP
M3mAslzLCmxgZ0JEhTADBM0isrROikzTkmqfQ8bELhuYnM/mfFMs2s6ovKaQ7NElXlceZILVtCJK
2w+WjBSJTPmn6Zy0UOfAvCj55tAw2WRtR0SsfBuGI6nPIr/u944P5jsiQVpevzwAukzXPWkycAI0
bwxnG7nDtfselZlwyaLRazrw8Kwbhg4upC7R3dt5V0Zu3C4NC/1q7m1mSSzkdVBM7a/TJE3c6ebk
x0g523ZXWfoQlX14CucXTddR9qxuF1606qequ2bp32VLD8rjvuYyJOTYYnllHUtug1InJWZX54Yk
drxPW8AcWgHwoRQyLF/HVSUN2FUEBbbIVUZ5gOmLICXRPfl+UJa3AQNZQTcGuHh0nTP50MQLgf+v
O4ZRXOnOHLfe7G7DZFsv4rBuYzVW/VbbMSVTjO41XdsHyCQqj12uIsRFH5eU05xgE2nP/Lmui5A2
Kg8bY5yAbcW+HlP6WUPqvMjoCAjX1sGrj0mUZt9zP8/se8rr3m3SgPudWNwI/4Ma3IOJrtTUIsI5
NFDseGilBrUVijMxyIZrfmNa3G4Gqq7yS6gd8HBvDkb0i9ovZUQc97RMAMwYA4Us2bVCrcO5qOU2
RVLLeFBcpDz228cGnsgE6Cy3EQOhFzHth55iR+fkl/2mSuEVT+0gxUpWHw2m8VHkaB5dDkEh1FZa
T8Li1nu1o7nWaYOET9CK+h8ePTmEZeEAUnkHC2P33lqx8JTExleIu7wVBPKxX7w7xIukMEQPrwiI
GuCReR2c1aT3aS8oM2o2i2g6y4sUOE9er0C/BGpISQTEjM0Pe88u7/hpKMa4u+fvu3GkxvVnZj7a
A0fyR6TaC0/eJCraVoSm3yvNo7xo1XAaYyzktBtis04R9QQDxRVUoBe4xb+4Xw0pqTTNfHuM1l+8
zERAxCf+uCBf7q8T/YOuG567VeXavQPsI1USASxGa2efMx3MCZUqZm3VtGFsiT1SHKh/jsQ7O1nN
1nmVHuxo+yj/FtMDiuFNFbG4SAI5a16zKZCyautKlOhpOJ7enCa6bs2mSb+t5YUUy3pi8x6mR87v
vYbYLGPUZcGxbZC6cTLq+HVz3+tDwflldB1tUsVybYz0lk5wqYnzO9E0LYYgJrtPI0YDst/Z5CA0
N9FHOfIdi9ZJHhJTbj7QQrr4AphagohgpFLdF8O5ztkBBipUCccBg21nNlKIZi7OrVxrYwJBQf5d
a0JzF7rWC8rMcLUUH44Kg7MWZwN+PqxZ1sIirDmuKQnEl5A4m9zyjthqIM00xzEvKY7G8woXPfGx
xVxRFb/RnwdbBjmlIB3a5Hh5qaQy3UvtD1xdRUMs0OXYgGBNFYRimrvCLBDgddyHKem71AAtoda4
pUFbpYoAXh22rBd9Xs2N8IUj6qSjr1nUoc8a+Z0kwUW7NKvALMbUycZMMnYM/5d42QP863c78ttJ
0YqGlKtPgPFZHDAcs2jl2p9alSTlwwtYNjE2LOTye3KUtTQuwUvUXX3VhUQPgV9rTARC5GMdcp2p
mYzf9WcWojtYOF0GVmE5Q9jvl5xDnzl0VBEg0kZrVdjZwYt1PuSkjcCdkK6ITx0oq1W/hvim1atX
qtQ5WQkClKNtEdXDyUZ9EtXc83tvy+JOQyMCJKcQXDsRU3M2zow4lXexLkIfG9QyR93P2IhvpUkM
4H2ThMJX7i1zgJRHW+BvC5F/oR03DKFuHq2QsZjihbptoy2If3jRgp3X/Eubfbk7/CU8wAgKhRpX
NgtDppQknw53r/gatZJKzB62qkxxm40AYL9/nSwNOjL0l6oxxt4K8w7VzHgeUJistWwUQzpBr087
VYpWKyg9qBNK9G0iEDjsgMN98+DQjY6aA3ERuvAXgwuH1BoYGHFUUgPpuKy/1Iyc9wXrbjMwkkTn
1sryN51J1xYmjHkSSZ9IT8gMMY1pOpsP+mg6C2UCLK4PR5HXeuPy6d+WWjr9SBRje3RJ28YcIwbp
Mh8EnpBl3WK1a7ajP6OgunXv3dMh+06/7VNFLNXVp1TawmxkZ3p5JfCjalrRljAaMlFZHbKHLTtG
9A8V8BFSeIWxDLZgJ+fkKCT18y7o+6NAf3AN+qz0fi6x3dEINGVNuYW98zj/5A3SXAW70x1fGHPd
aB3KPX8kZYeJPWAi41OGLyA0l88XA9C3gzBiQZUKZE1XNJRfTB/7n6pQGuR6dDQ2YMaNiu/l+2/v
glIhFTxDUKd+z3p6Kl8xtXYyHKUCXyvZ32XyWmuS+L15kYlIE8gVl0mi2l/APNLAJImUgEVV+kxO
3JLljepyOT7qgbrDRhJIK33XmFSgbbR3Cg075PyFE90zB9VROCZic+YT4gkiRwhFvbY8UmGXcCmU
Tnr4Qh34l7T1KSp6gUaDXX6bxoCvFgfWw1b/IylApzsrdQFxDBNxslPVa4cIVz+xAwTf45nrQ0mZ
1rsYZNizYZKgIw4kTZTO0n+wiZdte6U7YOXTkiyWirJqjT9aO8EwxyeMb1mLcXdv7OipiLUn4DQw
ymxJoKQBWTAIsDZvyDYb0Btmbd198XGllu7CGhV7qCcuEjk69GaERaGH0LMV0BV2HGt0wtkX1zuL
EvS9MWEaE02dzs7q3ckUWrJrWX1wULimmbJnYXuw6cOrvSrpvg6cZCiY2D7f0vtD5V3loEvrFjFD
YSbbuKu4yo622ctDeXnQVj44Imn9sPxJ6j+zryCWRxQ7rea3ntG/CMQzHT6+dZzODQgVo5topF6Q
igCP/ujYLOnCxkiJvxuAoHvhX513wYKWi4TxJV+CInfJRE3uel43cxUJ3ZcjVhCgtvF2umRJkxH/
WtPThEszyg773aSLU3a2A5cGF8QdO2CPpxdFWtTTLaBvQQw2V+Th5Luiq/fJaC6rQj1iZ7H6eDR0
Wjj1w6qmkrWNOS33PHAM/NS9DnmuoI4bOcpHzWTNxV2Hx2AwTddNPmjGVG0WR0plPsmnn0Z6kYAw
BDCR9uvsW1QnPDeX2J/1ZsaZPV7rJ7Rx8U05prkZ1OTqt+J547cZ5n5sUgNLS4KE3uY8E3Vj0j67
O6+xGf/jukdlaxW8Ixj6/+L+pCGG4J9YDTyB1qT7JNUnlQJQcIx1yFGCzwCzBTvPvvEG68JRbH69
RiTbIJlIUqG0YiBzbYQTZ2DfH/G1awlsAg5TQIc2r5nJWWXPYx2h+ljv3+DIm3Kg5oza4sQpxlOp
erhh6JkXLyOo+PnlUt8ch6cXEYQvOI98MwSFDdd2QQLCdfsN/r6DkRFyuxmBG21iENEQ832derTv
V8mqA1Hmi6Qwp6FK0PfUj/DmmvodFP/JUDPx5Ro0qrBx3cvjelGyPxgORINbXkwGyo6zpFoiMQdW
G11bbENAKWc0AflflAznFDYRYm1TOwT72iK4B46iJ+VswlTgjgCkliWJUylWwdRosCcHca7vQ+Nt
C96VqcS123fBAcDUDboPIUigXf3QyWkoYYDCqraXhY+Em8g12DLAh3CZeAGxnVC8YoMrPgZpgyi/
cJJgkGuXwT+gVCvkdJxPDSt1/LWPmBzPf8EkU+NNnVafgNAoaYK/ZkzPkbYlZjKYxOaih73DKDZU
73a0minXZ44avQOSe0VvfZHieGqCNrkMNNHUzEpqs4GKncmZhsRO5joSedVm6/0CsUpD7J4e2E8r
spHdjZZe3C+tKVcxv+2KiAXg0rYrmdScImtnqKMdpQ59QDQEw52hsEBLKMkrylGL/O/6BsaYFYoH
hnvocYItsNXijyQWr3QP7SPBI9B3P5CmYvqd5U0C7+x73Le+E+kocu/lE/xRf2nH6gSluJEtE/2R
nodPlwANpsugXS4f0U9MoxTWWufHXK/Qepksc0CCYCfn7wERbNxbe4EHAYKFhtxjxM0dAmiknTbC
+TTbnhrK+v2IDnmjlHrK8vjwxk3jxtnfTlnvcrG5/wApKIusNJF9J/JFFvmuErl0LxxryENIICNM
rb6HWyfrz6pUf74+eo0lCK7korT29FyjB7qPIUGccuylzkOFQi9I0uQd1uk06/2MY57ojP8wUOMX
BNyDDZusxNT3jztmdvnEB5xYLli+8tqA5cBOMFdvaYxfI/ln/BiFo5+PvXv3LO0XRPEqjtwuDv1a
W6T7pGvgxbigO1Cdb2x6+dfjeqkZMsQCwF4qR16htt6QugdAenmlOOvnGTQcahoFiS11HhV4vpNX
HuRBDzbcBLzwIvqZVZHv23nakEnK7Rx/1WtoPLe3ldkrv0fLIym5lMLwX/hCUhm+ohao5OEZdQnL
I1EeWv9H6MnXfYvGZpC/Wn6MmchJIm8O5VnvL83a+QcAprnMKU1E9vZqTNA9QNypHe7yo/zakqlW
5ckXw32QdMA8CFPs07m/lxxU3B57JcG3jCg4eG5SnKCa7Yqyqz+Y2SU6lZ4/hzfV2Pvy62wQOUEB
xYaOd9iLIN7NxGAxNXFlf7PpOUxTq/zTsii97CDRRvyg+KzwFWc98dwtgUmje8B9+aCuNcLjKO0g
9PWiRJ9ue/o7Y2wycoDKIWqL1R6qiWwLyio2RUIFYlICPbBGng8Fh2TfMI7E4yuYOcGjJ0Zrdcrv
W+ZJBxdnOHFzoSnJYRc75KVH8JZ1hZzn+czcG2YMcnqIdV/PhiNn7fLdL1qJ2RjXGsGCpmg0vxwk
OUDtLILPeAEOGYR7CN2eQfY9NzbRlyWlewEGP36SGQobFda94u6S4A0LE4l62aXhoKK1FShpbLMp
uF2ZjvDA7xJ6jA5mu/Cm/bmhHDQBa57FRnntY+s67hac9nJrvhwigxSj9z5Uaa8Dg4i60mRHJ62G
kt2R+nUGtLStQH5mRYZMuRZwlXzytD7eiFUirc7j0IOCkUmEMa6sgrxWTdQ+UzPRFI3wn2lxMhfS
CpcprnwZkSiUFFvpOjLwt7lmOS8uX1g6lWka4mNBsvBqvFxyXL/epeiQQKj7AAcVTBku8Nu3nU7G
5GnYRQcHDeCtwytthwHu6NNHF/CLM+txwbxteGjdk/vKU5PgImzw7S0Wq31c8iw6qwBY0dmhABxX
qFulbJIfNnbuVnLTTorKfi6wBdxuio5d7PUt2o4j2f4vY8agv0vty+2DXqz5fCyazwNBf/MJAihc
hpPDPCYBO0jlWetiVplREu8zkryDCFeY/YMnp5txVz2igQakHV9ObUnqnM0KknA+x2VyCAF1gyzt
6f4MglO1YnaDwrbqWZsCgpvBUOV5WfIMc+V12rqgx/FvbO1vn8ocnWxWOhCJSaCQtb/MZuPb1bL4
R4NekBBlQdDM8JG0vgjmgBjE67T/NOTNlY58nsHLMQ2McAlet53SI80iX48XoTtt8R3q8FGsA2Lp
qUV6OKZYBw7Zg13O3TShXyPhBovMjLByO0zDm7Kte1WjXgbWMXL1M+TrzRW2ADHPTH1O7ZzhkYv8
zXIlMtPwpW6dXYD7JERTLsXrTIDZo62BJa0i4SDbDzXCWEugGAxDAeSD9ozS0hjiE90nNnK4LR8U
jj/OXKl1epzp3qVDecqBUtFzKUzWepnI8gg036jZA7DhVNGQVHomPOg75itvL30lU6xnQoyq1PnD
3lDOn3bdb93ToKo/nmuBwMRTJlF1qSajIG8lhWv4siDw1Wbxrr3JjeZVGp//QCPF+H02OUnlf7fK
lsKHEJoCEwOLw3zCBdMARNcq52mlnAbL2Dtipa7r9rJKsIiUxzEjWU5XYKAitIIrG324szbxQgkl
iq/uHagynda6F7h2jWx80RhDMpM6I/crH5ArSDxedxwRZg5wjRUYFTRVav1Ka7E235EOcPL528gm
LjyWFAAErJbGNfN0wMGsz97TGf6JiXu6xNnjrPDDUgktbvfKMzBr5ccvA0nGYbWzqPXbmWpK7xBT
bRZDU10tR8M/R2+1598h4K9UDHH8baydazBwsgH+gYqyiQZNnqfyys9vOSR+IyyQQnKkuMZQEVdM
mDd/qYjVOBZiRF0Hf4vKMMn3LL5Dqp32H60VgK6tLw9PAUFm6ICqGx8fhO5RZdZOlhOX33jH/wGg
5N4II1/0GJ6GzZXBuQ+MmC3KYopEWwGlRd24jta368jDxBxwU8tt+6QIFbHsPuSRmQ0ecxFS5C7f
Guz82pUwJqYOq/Rh3UmXZ/fKv9icItVb1LQyc5KKClcpeKU0mPBm0gaE2DCwN9+Shsuxy+ECcFAV
hXpPhg37xnkx1hTPYmyl1V/IAChoQViCp85DxjGCjK0SIZ+QbUkL/uvP6Lpmp/SRTVzsdEgUOGvP
HgyEKdqCYsIJHzrd2FQeTvf1GbU4Yt7/t6Os0tGDeHlaWzTSHXw3wnK4xnPoXyGIIN+TcDg0UAYq
JafgMm9XHT3dlAfAB+CR4YZQQrMhTO0NBEKsDrmPEvU0tf1NomSE5OQz3EpTDuBEuCVDZuI77ml5
/9QMrmPGbrlBMERtLHmKIp0jQeuYqlbIBYo/VEjEs6/l9T20uslSCXuA9+iZ7u7+q2wy8Yghq6XY
PCOqxWytXtFz0gF6UkADKJLLxP59nQmdy8Ib4ax0/v3DV8zubTl1fdQcRcWvodcNx/PgaLPUFgTS
mpyE0qdJSL/0+byWHAODQVit6Mt1JoGajXGRzE35AKCcVqqgo7gK0Ai6qtltoDdmIgqBET09hnxs
OofXbNmEg8iDjdc94nfUdUvQcLI+IO3nOM8p/Lhqx6ZGO+xo51J6pjGEIRKlLqsdIM31DY9YsTOA
IlKwCVNQnSl8fkLoxbseuw+nGBkiVzVxPl+dcNznMPbR4m9KakfX+75wlgwblOoViK4sBke5QUma
6db0QT4HgdsZ7fHiyDv4FW9OPXBnlthbc/7Hk2GheisEx9foMpVpwrkkS3VKwCjrnzlh291d9bS4
6JCGpMheu0xf1B5rS/1J87MmjLDeXil3AmGFoWgljSSLhf/+ZrbmsjFPVPDZ7MxmsZQyrN0P12sz
OmjAtEZUAL57tNOlEvbY9eYQDkQ10SQxIUU6J9eFBVZ9xJDxtgdY7nx5vjapKKiRK0+wMMu9IOyk
3Xw8n5Vb7zcgkTahEU1VHcqDvOLll66VuDd38uHm0B2g536M0JwlVj1zBduQgbOTy3IecUIFaVH9
Sb8hCyj0r+bapK4ca3HNmuwdKbJGCJ2ePl3ZnEOuJs62pfVRw3GKPiSP5JZqPhNe1YZ8uLRr1SUW
8bWr19g/z8pSHNeX+x571daRup95+zAkq5+zqMxcRYZW8tPGVjXu1+caRUUMcye8Z1Rv2+En7nJh
OCQ2gRhgxn7Wvgvz+KD+ZvXWKng8COJ19Mj9p36tca9o+CkRvyoXHL+pY4kEdvQpxv7uQV1W0tgm
uL+MiFEiU3TCF7qvK1FYBvdHbanS+ksdO+GVlvdrmehM5GLPgPB4jxnu317vv1xF6I7nsmDXo8oO
9iNACz1sHSuVLbYXE83ejU9wbgRy3aJOJI9ZxU4wLy/Bps7pWoo4l6+WZBnTIkxnQohOCzb71/w6
DY+V9eWLEUlucV9P4Ay3ZBx5P82HB0hg5ib78qzGrWJyVZHLAulsyjYEQMbv4Ra3TUvwlmiAS/wT
+Ut0OUUt6uiD3gxmtmvSmQ3++gHc5tw1h5VEauKE3ofM+bKbiRyBs0NyQdj8QWx/+8DtLlu62JLF
qunjfaZ1kWXx78gKWAxOP7GQ4/6Zowldz3NkhPiIKcKjxGDy8Pgq88CEbsnIkERKUgUf8PaVa/gO
CnTt7R2sEtHYVSsSlxeT8m1yMMSS9aI0oQgJlZQQIEOXfEZ2RRViiq1/yi43Yrz8XyRH9SX3X5EX
yGQgv2+9i6PrErcepmcPEA2nR1nH676ENjYLrLr+NgTGnatmJZN96OUfc4Xg6yqbZRowkfOgGitO
hKqFhGzv0Jr2ulpZXaJQGtJQdvufait0Ju519G7nbG6/qeovs9Bo096X0V6+xIvW7pHJLa71Y05J
8wQmi6Vs4r1PqZlh618ofo5ERBbbuwDixQX5wErA2+Hg4BPd7fzj7YKWlFFdaTuN7u04VACsMvCc
rtRBGyE0bsYFtcx56jUHjH0DFWzDAnENreqXFt+DJpuXyO6BjTyS/TOZZ/B8N/5KoAwRKigPdWNc
IN6x5ftFUWy589s0/9OVfnQexgIqFLJ9JWo52SpjTzHZcXsGYm9PrFjahEqK8TZZFjEVM37yEUsY
R0QPml8Vlb/nVgM0DIjbFtc/WWtAPQevptnHLsfkyPy5GnTN8Lr948/5AsnzU2cx4MzK3/yx0f4I
VJKeivTYi0u0nV3YqN+rdUthA8XidzcYBC0rgwstbaUPKjtNjPwL6VWG6ULRRm3YWaynWMYh5NJz
litlgWzzGNebeR5U0/Wklxr84CipQO1rpbrVG74z9WGVsHxPOzTCVO9bil6u7teo/9qvk0+YI4LO
2naJ3JYaVyIRNQXTP+6tafc2J3jF58ZxxE7ivHRBLfwz9byX10wGP4zYXeL6epH4nYGu2S3VK0cN
rQ2PPj3sfu5Otr9BMgM1698tTVo5Iwi8VuSWYC4fW81pBKqJ85izF+jdyVgXJSjCluwHmNe5QnvJ
tqNr/WlR+2rdzTPf5lx7z5zlJ5Iah9r0mYBo8yhqJF4rdw7JfUEmCpQrtfIyAbofOpkH4CUHWMFw
clDOWDBR685MiufgejrbQB98U2WcWvJwZY6jNPlZ6Jb4nCVjCCbbtla6uToHkZxi2KLdwhdQeB/F
SI15I3u2H21Z8Hcx0l0kHpKq26MqX+dl1Nn9KQqGzZxMrdjeO1fCbJevrKPQ7LlSnmV/rIvTPjHM
XeT/f8gXLiZS0B6QQU9z+wtX7KE4cC+ZzYC22AGFJrd7oZZQpQfPvGVhDKvS1DnwiHYozx3PlMCj
7X/j3Hqa5jYA0zz1rO5NOP++BxCkbIgge9feYTClK7zzKPgBSObFrOtoaUZAXhRQK9bJ0tPItF3x
GR/Y5BcSY1vgA7/5Caj/MilsBmQj1pBcPawPz5vjidxxmyriCZAMZ8WzRzfP4lbyeyeXybsYwg2J
OVmvua/PfHXwmlkzcGHTCjqqHOfEXOMopXASQVkBXnZfdLCRfeMje/0MK/TaVFr4buLx9imc7pp2
YjTtyyK7noEsP4ycsvclNdO0uT/szQ+MtnPElaSESMo0/PsSmt4X3DWTFMZnnj4oUq4TB/Mw/TpC
s8gMn+tXfJvCPmX/mwQs5sRAB4jmFRcWEuthpbRSimMYzuPD/Pi3iNkqdwDvCQIMH+YvYFu25av8
9D9H+8KbE6i2lLmyGZN/DrJksOuJ8Ke7rclycmmHoaBYxCnU+QWLBf5lWeqT2pbaMRDt+c8IQ/ze
sv6vGHTPZqMSS26BXd9EKsP/ZCffaHiiFQqQQ3dA52Xk6RocsFzAXf0aFXgQKqGQIELzq6CLVfNo
SA9p0LuGT1lIWqIanmJyHtGEk59xx9y2PMEMWDqnuk0no2fyA5KGMxwCG12I2ywJX7nTzZ70H8En
GFJP1dodYTW5mlrMLbWreJyuBeDAY7XCBUHF6VrqAwZFsbLs1AQraBVaTf2jOcvEgwSsyxvhPHeO
W2/fACzZlg6rY1sGT1YY10XueW4TJpgTa9SZXxn2zF97N6u5If8OAe7+4SVpDn0m/Jce2fHTojJ6
jDGfJXZYGSsOFm7RW7zBcMwPfR4MVApbd05poumOGWAKzmWxN9UvR9FUe0YA5aYBCmLw9CgJNvSv
cOuAUWk79kIpAQNHK8qLq5FHHQerchTgyMNjWTEYXwf2xAPYb/XQv1SK4L1nKj50Fmt5bqyzmnLK
lt4dBMzNHmAvZQWb2pclfTP9TGLHiXMt1cuZ9jH2wR7G8B8bXD1AtsXhRRSS3g6UW9NC8MfOsKAa
2p54cNnMQuFObUv80N/nYXMIbhPM5HF/PX7BEI8PE21SO02HXVl3KslMfw6FuBXp1U0PhL7x7Vzs
Oej7iPNOIQWfBXoA8g97pLtB/kkMiLIb8gsGhNNTndMnkJcaopl2vpHeS+O9o0DTh4eDF+EuIGbv
ZINPyQtUPcPTyp8idYegN41bsgo1aGCQArSVJBWi0wtRQU0hC9tZ/gb9BP+RH0JK6HcX9Ns5CtZL
4fNOtLp/OvHI2pN/gtoBLqvyuswv1XoBp1FdlmDhVY/HgKUTn1LOGgFDR+Zaau1M1cZ3xQX2ojqS
i8IrNvEeYgcvNanN99uEK84aPQcw7aArS+HtOrEiuTDlZBXUn0X5n0OdF0mUM8++UZbZYlcFJRsq
/m0woifVxHHuR6IawwE0Vrcgfy/gRXfoD3bRqaiAUbct5m6Y3GQHS3FvXUnQ61Iu0qt1LYFFvBL/
HsRioQliDcnUulmVQsCQl6FjU7f47WcFCGiyf5lfraB++es9qjbZtcdvFs9mRQQhijT83sQp8PCr
PitMSTi75t4LF4Yvq1AVKPUI9l4rBZneZ7Epv+/PNi2frswzA7jt0nveg1jkfgqJdGkmHNnjvFZw
PspAwa7MvjFuqxRL7g4mX4CnjLQiLpWKEAsnOhNPxGgrXa1Ff/31u5fmEBUtbnJSIDVu3alx2EiQ
d8s3yfsA3fJUJU+CEqfAEl/icC7MIaBcLcvrZmVNhj6shqDu2XN7ijjjy9B7Ezz0sH7FBkADLNSU
ZLRlr77jgEytZVaCAuO7748MNsGrYyPG7vWC0FU+d/TWeT2Hhg5bHLEPoi1jgu5b+HuKJdzC+EAv
v1O182274wpcmg60uEjkDHQSx28Gs4iySV2V8/2B4aY6pscvsxUlDPQ6cL5iUDndWO/c+Z0QTYLd
nkYtNPUM9SH/LTPrrVbjKTBeH83C50T8ZeSmL1mzH8xiVWHYOsyhyHt6ZXIAS9ryd8Xp/MokB8N9
FQKhalkM9SiB0PnOTv/oDrUCZE3PiSTDr6Lq6/WCmjxKEt3JR8qtzOElR8Ldchnp+dwoMVhLyZsU
Zqqx6OUW1BH1QHDmQCJfM9PhkCCsldk+hU94zUbGtJmkZHtsycdvXaiHkLbMj/gbQrVt5c8yStsQ
9hndjHdOx41XhUCBh3Zjn6yQU+tUxVEMSU9+SofmV1F9l24+In/71k/IleX5HhlkOHUFYP4erJ14
ZS/JvUDnET367ObQ6iVWmhSkSl2lNmWT2Ud5UmAP8eudywnidW6k9Y3F3ZmaOPl+6Y1c7IEPINaB
5uKUd7At9E0ODfaqldb0v8s9OKpZ7RdbsIkknfvLOoFddHnD5vil6/qu0Wkzol/CH1xFcszGO6ig
eo1E4uj437v66WOqix2jAsvTq/RZj1XWcZFWDpTzAWH1yu+ol1Wguc+bvfwzJE8af6qaRoJ+rJ9V
aDGGP5rBfwWczdicwoqCP/EYQAyX6YaU5yluceY7hLNfpflU0hUrS9loBRmbktPnC9qaGN3Ttl/b
O9zCmLUuwcB47uW6J5yKsxz65ONAIHxl1tJEOzF+aMICFBpJmRoXd5ADkOW+Une2I310krLtJgyb
smrqfyN6thacFan9bgW1m5x/EYttpYHdSDT4cNBR/hEZXVqFmsob0+3CaeCO4osiyK3K+VD2lxJL
IwVpuTXpPSPT7T/3IksX4HTwY9RXbMsT/E5CYU+CXrhesTWrLS2ZHdrhozgYbJPNiYtQEIjlQvag
xZ5LfefJSSCQIc6xK0uJ7J2rq3xl7Z3n/TFuR+VSfdEyhrYKZ78ZucWCAYvufCvK3xy+URxXeSz2
5tu7aX2RBaosMzfVCoK9Gzlxp9lfjPoi1Fe2knvn7toBAlEphP9VJoZLYlp13ST+FJKssADFmEf7
LjLAdWR6NTa2XQx3oNlNsXpdPd2Xj81ItJTDpWRWOnETo9KULRTt6KfrsnENVhWO8r5SIt0GbGER
UCJfzr3sC+hTLwiK03DqDQE+rmGYhkriRNhnQhx3F6LVfi9mlg6EYefxDqSKRHuHEAuHYWVK2cdm
HvvsIKIW+R/s4Z9ntHBdutSJJ5BEk1dWx6P2QmSAwLCTV5v0l9LkDF/IBQHnaX4ZVIaqbXsMUJFR
TtbAGXbzy824asKZq67ZFGCvGD3zM5hJj17tBnYq284tO1IdhHT1MKEqHnKnZtvh/E9+5rlsQZ51
KMDpSGuS8D4Kl372EFeCCg3qC8Q4UZTxte9vTo27nrEOUIc95VFycz1cTO7PNnBgOg9DcYHFqc7i
+UzGtczpG0DC+QdjBBQjDFoYv+iLFRMctUXlTdTgcQZyFiW3JABqilRoRpkWwaiBYKz6/TKT+quA
zHkj1bnj+WdL1nfQevg3B1hMJWlMokJXRH9fHHXaHtYBkAzs8vEPV3wDkqj+7aNhqYJRPFQz0vFs
vf/iIUzYhWEu/RUE0bQwJ2t9EkggttlWN1I6uMztTk5JyIf4yi+CrfvEu5TKiiTcwZ6H++AM3pnZ
ZtfFtn/qDkcka23VE1+szmor1gvJ5H94wHTMJuU6fRS2tllEb1N3UZTS+1LlW5eQ5+QMx6hVlMJP
YMCUk1p0s7QGsOm1B7eBrF4lL4RjWEEWOsW2D1QSa5+zDDLpziyF1ChB3T1rgOY4JO4XzI/K7S6C
Cy1c85Gxy5Br3+vOGhcXuQe7pzuPXCOH5NB7fX88wb06YusRz/Dgzt26aZRA2FriUH4q+3iFnWNY
7Y1uptrpRzqCIYHb0j/Xj1fPZx79jCo0SSlO0wK2s+FnyBhMOLOTJ3dkSsy5sDbwvAr84g6+urH6
nABS0CaPR+ARq3XXAxWsg+Kk92rQpokcuAibhWjFA0Lyt0cWlFIzj3PfL2P4mxzgyTQBIgZrQk+t
1Hft7apYqvAzNmtszWTHL4wA89bQxBW9uM2uOCHzsvtbiQwN7MKGtRg455WtpIvvwZrU0RelM2fL
M+H1gHNZe9nrxAMHnEG1kkzqwkuqnhs8Q0R6HLeEglCP0cB67GzuqfaLEVzMQVfexXFhiA/l20gd
e8PBI92Feqf/Qh0RHzTSF5q2Ck3giZQrl3VeP5441mWTsl7kWCFcIaSAtdGSLJ2s9mkleBzFx47a
ukOSwULWC2/XidY1JhaKiaYNSXGleyJZ1aqVsA066jmE8Kx365m/Mz3qi7wnyVNJzfxH7JqxuPH2
mpwlpDJbXVX6+C1PyQJ2I93JnuTvsgq0kPqHIGRKuJZXsGWPBEelLmwfQznufb9Z/wfC5wl19xMt
oPet5lDeGHNCpNyIkCyy7TtnGDAEeuMIkbo/aZLA/4o70Z2ajym0jMp6p8KH8luO2/67e6U62kjH
GjXQGbsWcSxQSJ5sR/eFCFETM4JqzcPu8Gzu/oP2yf318iuob+xJV7yqa6OtixNBTrV5e+Q9IKUr
lb1edR4vNXBejm1/NMGMerzm+AhV6pT4jqbsxx7Z+huqNkbXMfHLtE0uS6e0+5ClnNCW3ncknhzZ
jBbBJHzSHtnyIUDbzzAS/cc0vvhECBHSZ1P9S1mumJedCepW8TW23GfchkiR6BhUmt1WG+97L4NZ
lTinw+wVNVbPfBfgQqtNsiNMlEvhshE6v3UAh5fJXukQrq+RsRppGAHrzZ6vJBBqpgak2CdkeGdS
6XGry65/2WuIbrwI2rHOCQyU67NILM/VloRdnzv88bzhKo3CTRmXcblTLrHR21FCKYgR/zqeceAE
lhIohWkAzbSp5bDSvzU1SgrHIX+QMdczwsuy2Xrh24cA+FFYnft7jcN541G6mXksYkIsyAykIm51
EC2bIdhwGAAqhIq7Xqv+EpDUjy9sSADuICmPPAvSjpGkozjN51a5Pk666ghU6M71utgLVOjNdJrO
u+O5UGzZ7FtKGlAm+KpTxaFObaMtoexUcEkLPj5NGXMuVLyVCAbTrBZgKEvw8ExbjmcjW5vcTgx6
1eRODhRruoe5KhwR3/CLXR5AFLDjC2vSgGvDw9lRRx0Vdv4GEJQLEEOqs/kDfITkAhG6POb2yoV8
C0xMjc8nfOdIEAOlcgPKtOywtuH4EzUMmT+HdGuO+kc0hiNEVoxwaiTElDlfN1qNKOBq2ilqHV+9
8dWBDyDRfnN5vBuYI9wBoztt2+pLu5XHRHgLdW1s3I/O079+wTwzHN8v8NEONJvYd+/QaJFf8DF6
ddpKGLzd/2MQcpgBVebAzHR+oa3MI2xI+q0CoCygrhzay0S34OcBgrH1BOc865hQUqFlyD1IjMLn
zpjRaU5MYNUqS2NyoFWz4k1bgqZkKHNI6YPOYXuFuGtJqIoS9rBmOqLFlBYh7vmJ67U2hicI8zTk
QFIngjfuOBCLTwo2klfsrX2HZs6gaJnM43ew2Bw0pNpHVx9pvcca1cXlGvb40r4T+xnCcxlGHSPA
JZe7FRV+79cHxLmHF7T3xWpcEJFoUVHu2oiMsE/CskbW8nHkJTZr+jjHYha4QRreJLQrvyYY+61i
ogHx4yYF6F8Bfd0HXlCSQ2fkfdxdZGuHRL3cF70FbDJMO+/Es+XE728B1N5aslGfM+Od8+sKKMLN
nnKLuUbuwxnZ/+Ii99uaAI8Iy2Amx4F7SN5y3wSIjVZIMSMFhYWLBhFDEhA6T1ErtHCFocV2oC2+
DMXFcNmfO7z9EMXiCg4uoatqNj2LZ/VnuH4cXmrvK72NBtCgCTa6KBLf0ki1u1ruWggjP0hkujvc
ZMq+eNZ7ir7HC3dUf8mYiYpS9TBZE3m5Ayw2b1BiR3Rrmlbo4FnO5g+olT8kZ/dO6CQKR9kfs+qk
5AGdZ1de4GXKlPIreIqUim85h5y/DbS9jQK2Q6x35TTZaqBlJusrUxG0ZDr8vNbxHS5h8gDx7MZm
LDgRxgwJFKaFchAaKUJLyfkRtbQXEagwC/vgSHAWOTRrdfAY+dhASTSLzGBEyacFqBDPxhC/fSPF
wmMTSNbYyefefkGxBqtREyfhBAiygYGPMXLiTf56NeXXEWXRz7si/Fnlkj195LT3tASqV8gOpHDC
v2Eq8jTNbkJR8D+J2MAfDLnP/9j2F/mUlSdINwpzAAWf9qvuCXtsE47uiMLNNnhO8xNgDy1oyYsN
QfY01nK71h8DFWUkV+T59aDb2WXIfxP8TuBkwMLkHqQKgnG+LwB2cHzQJ+nAr4NaEhyv9eJ1FLjy
P1J6IHxRFb//smNPtdkSPtL2TbIIAKAi6LQ6Z+/Qi8tGzDbavnZ97LeSVzkTkyT5OzDr01j+GMUF
zplGGsGi1UbuM2mxsXxB8GHO5tjVyzt01rtLaQh3jFFjw1QZGig7lgusyXgc4E2fPxZIDAhZQIcO
a3m+zXYyFSbk2zW0WJskiepO2iew7pN1HltEb90zYKN3Hg62axnRuAmwKZ3V79XkEufwCAWESZXj
dSYKCR/FpLmsznmSRkejEkNGj59/xmHeGNKLdLp+Xv6RXYC7bWmEHL6wBygtnGvhM1fz7xnI6Xmd
m+2CWYwmF8MqgPFuMYW1Q6kEXBNBYRAZSjKfDeXK+YBzfVe4RsQ6+S74dh6AV5athrf0lR0owCLf
rhmbmmIG4TPJAVySWUpcKjIJ4SS+meO63oG3wJoyYdB3FSUjXOvcmCvyoBTiUPWb8vDAl8ucWzkH
9rumtyukNmSleBZyMTnl/h7Sj4vqnS4Yv+7wZibJCYyDxNUfBglm3QoP9N71uXdgllcT0rCQ61Ts
zFYFrQfCgJDn5KAhgWeEttjKr2Yb5ahCP7KCRXESQloG2wIUV+9lZWS/a1xeIYYyocHieHP/5cM1
Azrtys24lVTfalnw6HVEzCnTqtPapcCTUbvLur3b1McpCtwv4YBixhIn89lNPNSdsYSG0ApaIf5u
C+rD3TxiV2xNL1uqAjoNan/W9I9fLMTdTc09zmafexuE1KMxdamxqwWS2xVn+snO7arkV9MPYTi6
HYKDIBXjjpharzlWbYngCQxTxYDbz6gPFPRtd8ZXf966+UnczoVnuuhbiHh4Uio1TB7qa8MPITBY
9hOq4YJvRupH//3vJn5FWQB+hpZYyYk30ugs+Ad0Te0ZC+cYiXdy1cQL1iRC5b0dZELWOkrWd6cP
poNOlEC0tGrdAeuY23wHf7yv1YajxymFOQclDICRYOUG8wnLXUO+ZDA4L2dfIzrExtlUvFemtK5x
4/3v7WIDu/dsaAyJkZ7SrF01aM0Ya/xLoy2wOF+x+Y6jJJeThq7M67LJK05/0vgdgY9gfCqzKucf
2bx0qYNBOSR79yrG5gA4RO87s6wsJaK8l0GG0veamdiLHr+BBTm3NhXi4c8Ll4Sel9rLOPRq1pnI
eYZLbMVQ0mzm7aRbt4tOmaQlh7MEN5junajNxNDH7jeBPXGB28VTKf0n8wqEhOWmlq+Co/EaDRi6
Dycrk7Ro5V85mAIParEHRUoqJghbF4ZXDHD6uF/QvcHdthJcPNsNL9DxtugEcbH/57SduLs7NlHL
ZMEnC5drDT7M+vBO5GGwXR5An3UuHcogFtGFtEgRQQD/GhdcN24AD1p7CewSaUGkZNlob280nh2v
hN9qUVxrJMKyn2FwAsHJa1+pJJ1bpmTckRdsfDE5kQxgd7gT66L0+uriAsh6nxPEEbQPNi14MHkJ
aJKy0iZ05DmbNpdO2oHCfyntkRMKv3cEJ68Hy3sAsE/2k9Ge85QnZW+1vv3kRJcPfzmQrZpYHr8/
84p5yQ+Gt+qQBgzjelOK9kTLv610Brn4Y48pLJHp9HlsDvgHNfPlhNS+sFcC2iWPzFzzbrVjAXEC
BsEclElc4MZyMbBUz8hlM5dPCe/qbEirtyT22lpRCjtp1dFl9NG5CsZZ3v9VlemZmevbY63rQhYD
cgfhMmNFUMo4/3+DeicfxggJnlWWEjeMWbH2/vT4zXmVRdzBT+KJosiroSbLJl/OcTvIqm9UZXmw
JUL3bX55pLKCacIS8H/WA0ZV1vKFdQlzmjHcKcdzoeSX5VVXn5Fuol1YPqpNvXj4/n/K/A7oIlu1
g5Q1HRLwz9DoYqWOBr6vaHsCGHPZfoG8LSHwgAaPpXSkepMKNuY+RGa+osMnfDXOkz0HxNMe2aER
QSjM3C4YazPJ9kU6guvUIk0OENWxcI2kCxFo3aQGZY6OpE5LWio9iQ23tbKVLv3rSw3POds1ZMtv
gGiDIK/gW6qP9XmGuaQSouFsK8OivJ3ijnLX//bvse/zSlIwJt+QxwXYLlhrgIygqKW7WdGUpbTx
hvBuDiUaaC32G+GcBDRL977joDTUs28DjMnqNBHpvTbJUEYCUUfeqL8Uxd8XyV66U1nAKSZOnnRi
r0RbSSWI41im1ot7uoa+Gj0pg5rSALLj+7Bfqi2mG+7bLjfHn0scHpGJORD6UJPWgrKmTxIuYWJh
2phPLL7N1tPSL5CvU1Vp1RXP+SkxndSqJR61FRMyWThlBfCA/T0igWWSbB44b4Zf/3ZSplXguwjo
dixj20I4n3QmfCuUj48FMS1ROGike/a8NpHzUjJqcaOgp7/MBW+eveN9xMWWSOGZXYlXHsh2P6qm
YHbaJ7uZanojpBRLl4ORMe01S69Jss6yTtA9QzLFuzdshf++DffibQhziCNu5nQoqHxubhRw5Gtl
ZHBJvQjMbk/BrZe8qPv1OGjPPFKSv+l9zGOs6ahMKJbgykWzNbFbf/6T9hoZ+YVdZNrEZflVnsCx
oI8C++sPRqqSDvLEsRMhTbeKsaQPmCH8mVROMMOBJhGvnOwz5/i32Ws/WIv6kO2MrSNA5G8pmcTL
QZRLzkxlFHEJAywu6kPeVJUncKbruCht3tLjgTYKf1kb5UBpf3xtGWqzR3OyamlutlFA4guQCouP
gHnQIThsAEhyxZaTAdV1TaRny15nI1QQUkpV4DdFb9s/8cX88Tl6rRLB5vW/mu4ROQ1h9Dzi21Iv
7aBCMnH5xs/LlGA22FjxEvVDYIyflHR95j+FfiaJ1rqLkeKUfYBqsgBvo08TH/OxE7s6uZDKIF92
4IjVrD3md+FKu3bdkfPRreNaL2iD9ynizypMCNYEuEOgjI8QoJolhyJnZsg8WW2LqE/r04PX2o6w
ITBkx6RvMP+jcHqdp3GAftJFwkR7OmYBbVA4svwEsioqj89oM3wliCz2a92DQuWCeogHd5CcDMdX
DjhBcl99SqQbEXjPY0ia1iQHWIZA3VefWJbvDL+EE+ZuaS1i1FUEivJf1TVuCYXjBog3Lf8bn8eT
EpLj1Tg5bULn7st9vvWi2rIFxZHEwEJ4xU2QsJpxyo+hishXF81HxHOWDt5FJh3pdXUvobqyut56
d4LhgRNgARClkyfj39mDad2ncaIxtW9Pzy5GmKw9OOfxkNXCdkW1fqteSl0OKZob5ckMYsp0HgwS
d7htA9yaKjT34XKOvl+sMEKkuAvIHIbCcCwbV6Q2dCSKCTaBg41pJLks5oIp06HK/7McJQLqDLph
OFkCd7AV15efzplew2eyziaYbIX7NLr+1P/iqEw8FTtKL/cFPQpv6JRFLcSx4MZAl5AnOUx+5gNY
MOpDB1Ios+l+p5LKtzQFS1MmEGsmC2A97ersgWKexSZ8J3YzKU0shzGKxyiOvybnNbDGkPAc/B/8
4Mk+He1bsG3zXczDj4Y+VNdWVsS6zWe97U+TnfSTwcuE+PdqT9fthfzIKaGfu8nFipE0iXVko9g/
9bcT/Cdd21gCjSpoXmA+EWPiQdKleSzkPfwh4v7GTX3mTPtwcf0Oyt5koCMVRFn5NhcqzaLRBcq0
Lc2iyzWBOZaS223zwejQgnGYpGbsqj0am5leqUBZN0I6Y7Ha8RA8S1PDasW7bAqWzhXnlY8LbxA+
L1n2y+H6p63PGKo3ZFTCbUE+hzB5neQFe/BnMKedzdjllwd9pV4sn61vGNThLTtRJ+Cd564Tn3Hm
3HadpswCwHq75Vvv0jev15PxtCWvfJYh4eWF3JLqWCj5PhvwjD8NLaT1Y621VNcle2QhLELS1zNz
Z0sye7z606GzbM93u/wCSlSznOVuf3ecZVvdEt9APpvF+XR4xL9SGdJ8k9JMyun9Qvy+le52hT9n
0TsQCXn0XbXj0m1E0vQ7tnbd1pF6iXZM4fHIqA3R2Sux2t6RoSN2NHlD9FG721g7uvDXtMHZK877
QLwqW25WC2dAZ8B4G/17zCQGrbObdwLG1DZc/OErE89WA+EYSYM9BIG5emMddm1/k0oImpz71fzo
NuCCdGh2lX1yImcjiWqllwyVllM1TJwGm8HmKUk9KqJMrnHJuVD34Vw3n2IAgxmXPCAqBkQkMbEa
WqYLEl/y6MgG3dEniVZyYUOEt+jsxeQs4x4wvsyr8GxFkzKXyZlito/OFqQevH62Zhto4NFXrWH8
/JBnXHHGOFLd/VSsLU0t3Mi+btn0MDpEZGNs/9XRw2kX9iIWbiR7B8skB24BTNNNqK6m+GHiqCQz
1y4Kbhz5MFAcfroW2Z7PjOk/z+a7eWgyT+kIWJNznxMurFp8U6eLEATgEy2nJM69ximlZYmX5kZn
6DTFL5Vz++kXUe3l7i9MfmLfYtDI1vRXF2VyMToKFE7lv/EvKZcGyjmX2Sgp+JnPsIUXSyd+QdHE
bnBplh21kAOpRm/AZVXbStt7rCnAo8jZ/kd7jfOEiNZKt/b5ZKBW/NGaZqiIVp5PFDRCPkbcGVsz
+fqPydvv7c8BxRuQ5GbXlsvxpKG+yi2S2BuAU7MN+e34Q01ardxTl6tSXVn76DPL3gfPiCzaYBN0
QKKI7wpLu8exhlnWUOJH/KKNwjvKSDYuqyra+O5Fst1sqVGGkpwmjHxdjPYZVCsknm1Ve7urB6x1
nqNcjiAalwsuBU2z3ChRsCEAzAqIkpYOJv5pfV3oxkOtw4SOKzmQWZC+CWiMZp3JXGmSZRfBJnXL
OGI4VHyxtqE+U5M8ei/8VnOjj1P7WFLSiW7frrxH20J6cf2yV7P4WWmPwn9Damv9YGADPTy+Elw1
wj4jgurQH/tn/TlB8lAXP6YHjzxrzr3LY5V/wBoY9bQQQ+w2Vkh7IXT4djZ8JS3JcLahmeqyrCM+
erDdgMFZzJGKm99vn4vazxqdQ0Ji1jSJX4kfoNY6/r9vCG5S4NbUiehh/1EsQOcX+FGeDC54jhwE
+6edJfoJ0uAKq7DcPDsChuG08Dvp2YuihpQ3Ln6QzzRnpojhPmIy+eZCczMbGTo5tj0roSdnVsC+
A1kcNPWdMlMV41X3ZlmzyI7LaJNrG9dApfd4Qx6Jth4aArPn/HPbajkjrw1KKTn8GmNXXjw1iT5s
6YCHLuscsbDQsqInQkyybvmaCeGuW/Y/vu4uVCJfFEaFYNbGUAYXwQ70/989dkoDdMULhoVS/g/X
tJ4R+TH0QxvNbe+sKCUoKFHJ9rLHOM84GnxTXutYzerGjvKBIcDxiMlY3hcKrCCaCP56pbwbv9VV
v63OAbtoTtCoJ5x6ZJGLfn7ZPkIPjNbvOEqmD/CZe+E01+Gh3kWoMnbL89Kywnxltl+SrgQZXPGq
1BTZIN3hTj6Gw1uSRcMLqFAUtD9fZB/8ce6/IHXUb+iU7vSVUoNJLIRoFJL4FIqLz+VKSp8hHPPs
8RyIhuBm19nLqoC/F1ciOh0ljGQhRDZnd5LlDbykxt+rbHepkImDoxdHSli0vSEqj503Gv30zBhK
/gDdms6oeWEkJp/z7aOtI0R7gLDmJ9CtROWZoROTgDazOiBJkHGum1hgOQ7hFNFA58afqdwMGHyw
LRc2RZ5etw4sTqpgLAuzoExxRhjOyCTmSC8mYWnik0oX6AI+elMw1ZAhag9jaMnN2SS/VzjxAvKe
YuqsCAmHzsZtKYYlo6Fa4vrDgPDY+Sw3DAMXS9Q4AS6wRAzBDX92XycBg8LWbrFVnU4OjkbxhiRX
rrGdFrcrPxCwqN8PyI/0ePHppzWRQFkQ//8SYRdDIwHf2j89TihhkJhm4qCVs/XL+zEEnOakWnXd
pRHKiOgm88OXg0M0Pt2KVd4u6uKySNe2Lq1wG3Tzi3lgx5t8wl4DGzPxEhC4paD/fIF54acb7rEF
xxxWt0xX+Z02shZHpES/BMaG1adGiV68y9XOJQe6DJd8plwY2y4Ywgq0nDuFQ/m7xDDlu6GKeaEp
PQdn5fDdOTK61EOjhX2fCiuo68ylbLb03Nw9Fq/gUqfY6bWqEYLqkGFjx/G3hxZ6RVr27axyLbju
dr+Zf+r3qMixkOIZYmQEGrXV1OTpzl1IrSMABayXXtZF1RxOv5DxGHODE22alymU5p7JFGKmzwWN
T6V1uShqUQ+mqbmA7L9gSGdz/xBLo+XyRZFmRTjy0+3+RdLgJ4OCo39HVqspfkAcH0Lc1nQZvYfg
j+t0yD8ST8zKTUKv7yNYbfotZ3vIFS4B0F9cb0WIWJdkPDv/DcqYjvLykaKhqTSY1KOhQzCsIVKC
wBVPUnKLlSoHkXZBaFF2WFujThPxTU4s1ZaOQqbUccZBXv9qHOYcnf9htZuJHg+FI8xoutVgtCzN
X8fBMGfpQ2kUox/EQyJaCGIbcef3Mi47Jm8xyaosj8H0Oa2yQjzgLL28Yk0oBRAmF1oNbO58QbMf
pWAwUV/CR6PabdgKqKBytESi7xkGtuOBk9nhgAk/OQaWQ7MSGd/knP6D3vaCyFU/B2/KWj2fcc9s
YhI2jZ/A3ce10ynpCpnRv2EnV7l83gS1ZsT81/B8YE118r//ZLOK7S7PRadQDaQCAPLtpIU6HNfd
q/ZTdERGhs9Kb9x5/5Rh7OX4fTb3nb96ro0s7iNKpjop96aczsH78rsnjyPoxyMBicQkjM6djd/a
/wiGNdhwW1zVULaLY4X1j3MU4mqj42ieS9/nsve3gFMShosOLCCCsJna8r/pOU0TH3XREPgGmOcb
Ji4pNm/lN8bMNYddfIXsmFwDQJFPiVKP3UOfnwsyDYV1Q3XIhOSj8j6kOIKTRUjb5fQtvT6AdhD3
eGACq6DvfwdFz+2CTQExJHvR3aztpws1tHZzaBR7y0bYGiZbmofM1lvWM4w/Lbu98KbLd9PwumLl
ZxkDnvAV7nHqu7n0Q10cCRT1P42LXnsvypF9V2RSts/GhZb/wYpO/oZMX058DPi8WW7LYeN+momE
QBSZd+GL9rgDzCKmoO2urQlUSAkD5g+d7p2amgB7mfTW82n3q5viGsjdcDNTQijxVaIAwswgjm8a
7Z0oIDFd4DYm/vHSezyoOsCmyDNOZg4jDddzjrOx04IKwekAu1OAE0pUvtjRI4ioiRDb1CC15Z8y
HRHeUpGRGwwCJ8exG+fqY836KI6Mqtxji5OpwSlmbw4yAmCsoueb6Qt9IjV+0fUrovU8KB2U3RU3
1R3oRZbPiDdlnT+xxMs2A/1p+hsPpYf9BB8Gq+QE18MutM1y4w0GDoDiLnAZnh6FPvGBM0CycOZH
lKm7xse4IRwVBGuQmBenqtOejuVjo2CslcgExSxEVpTBHwtmk43Nfi7kStIQvJqtn8oZFNsYJr80
xyj0qRdAtBzzdCRwO/ocOaXzJ0Nfod7parGEMDvbloJ0F6Q/YaQ6gaXwLGaQi66OtFUhHE9gE+jA
Ob0EzeoJl/ECOzMoI5addZLBttFAy8azwvv5N/5ErKaduD2+Fc7E8Z6UbRzSbf6qObKHccPyonKJ
CZktN/a1wNm/hi/PtuFSpIFeQl769FFzi4crGNEXmM+Xccti2b19pgzMF3CX1mub9unhyW1uZ81C
VaMCvYGrHYEvLLvuz9n4NsupK7sA2lwWMFqO7q9nfoh4gNckdmqsV6CI0yghBlqbRU35t8ra7rWN
zUWvQhOjg6i98X1yYn70p0XNYDINU9loOcEyvGt1XyxYkm6B3XcZAvbu36Sykz0Joj1waoUY+t3K
yb6apW+rAwvX2zO6CmY7+POeBdKMsDbNZObu4mkK9C7TE01STJ3vbVdK1NO17QvfZl4riV9/S7ho
YHRWX6Ec+UsPyUE/k3Pjty/s1BgZHZnj2p821gGO4tlYBDHwMcNKGWOUQere2p2zxi0irvSXQvbS
SKEY4zFfebMgwat6cyAX0kT9EX4JkXSlwXSje0HoxoEPSbrxncG4XVhLwo7NLnYejVZfFwlkJkMK
ZwQ01+DD0twPE+qehk6P/sZMmj/cJdyMz1vMefrrRPbLqw0sAiNyBBQVPDwGb9Ityyd4Oa1qhrtn
OAWbxuigylsrZxg6GMQNvsiF7sgC0M/EINqfJh0le+ul9zb8+w69WSMh9teNx1TIJVpKgUdHcw3q
lEzkeRDjqACLUl9rEfBesn96FdX6BMK5g8VwqWxZcfne41hmYx7tdJTEdtRQ2xq79+o9dkFbPNc+
oflbau1dspYC2bd8HhAEeVDDB23spJHSoihUoAQYi5cT5iMc10l3R5Y2gId0XB679YTUkUTuI2Xl
iKNrqsdUWiy4NJTjxHxRlnh7wHDR4KGgu8ZLJqWJEXFYmbKzu1WBp5C5BgNQB4wPaSpyzVXl20sv
lkILJqvUT1VPMPA39tAtMbnTy4fxZieb1SE8RKSU1M8AyFE4z9uYXKKvzMtfjwCOSrIBp/WDH6Si
UGXA+NXWXTuXB36GEjr8lXEtybi5CkjzqGK6aAFSOeM07T74lJHa6PlOr1sjpMOksLnh9jEMgJ4D
vX0xQcfcbIKwQR09yIPpwmA3vCuGo+TJS9KgQjLSfnbBPuBWBDo59AsAieMD6tTqgZouH1NwWq4N
EndERORNs3BK7O5C/5hDJ42nYvEiefJhh2Za3ndZ9yHUiAeCzaW8g0FaFP7hkLUobGyI/2JVJV+k
POUueCM6M+jV4LhwByUzSEhxhAnGMvjHY2llx+1gup2/Rc9WfKZj0mkpXyzCfX+wrYHYebUfCOEV
6VGjXV9oJgNlvMLxqE14jw0Sp4P8Z3r0bx5CjR2b+ZFPhVkAGkOuMowBhiyIiIAcNvtxCT6TNZlt
9CyA8e33OZFgjQgHUPVdZfYqUVNqJj2x1oWDv0vgeVldvFCW66Ai/E6rlfiDE7O1AiCgS+Bdek8O
Wjb8HtdwXHQL26SROTu3bTOds3rA+xfLkq1hUQx/kiDC++zMxEg7kVQYncdAPJw3DHU02EIjEzXC
w1bG4evassdI3kpqMj3rrZhx9tpFddWLa+sdn0Cderi/8TAq06kOs7KLqOws22RU/4QhfKi1gpA6
QiA5o51D1cCEd7FMMjFerWEpKT+keM62dlEReWRfYByJTQJFT99Pz+2csz6mNoSwAc/NH2T3Eor9
eNIWnPNIEdQdeZX04P8GHaQ3H67yscS8Jy6c9WNuvKCu8QBkLyt9Q43cdvo4/7fMzFqs7M8IoPBL
X47aDvP4iIQwsELSNeMAVzcV+PyJyf46Ys+VT28tmp6gx5WWYReozZOshsGkDiEXgEBjQDaAqpi9
SXDJEoq6AY/MPIn1JjX3pu3JboSwOzJ2ISNgPto0TCzTMqsEZztltqHOc6L87m2hbATEn4nu4GI2
jChntPYmKs/Dde0EhArcU+IFD1AciLaHi50vGv9lGjJ9UuLDTTffxXPU9NJGKDZsIqHkHZAwenUK
Bp/SK/BjVkRUFfXW7KHIDyTIx8UhBu9AIiVbojFIzzZ16QBjkr/g76M9HmEK0GFeRJwfevA+Nc0U
5d+sc0W7wShvRBA5RjhQXWRAUaxLeuo2ZqErtrOfrbSOqRB7lF+iWUqjehNJYTjiya67QEGtgUf/
pwDmVdmzpklJKuquTn+bbhVnWqzVEKgVomS9PhD+AnOy8VlvU/2z/IfPMieQQOEDbxt9qyfyPLlD
Qhv883QgMpnk6hQ0HP5tTQv5OZcQOVebKMqM8UMxA8Ka5z8qw70xiw/cUcrV8D2iujmJuIgUgjBJ
ZgnEV7esHqrbpX9QrMXezA/tCxbp2uLr4f305gw+Uw/au/v9wE4c++RhHYJDfM+luhMJRnqi1e7Y
VDw2KIH5LtBzdbJhQ7L6Df3X4bIn0ouOLY8fu2BcOycFMQ4/gtTiCI5qnFcwAny5V+65xR72uAZ9
BH8t/9D1w8EC0VX7ovdsvOoCgKXhS6ZtdKXIxLUPao12fcevsz6YFUMal/uDtTZq21JuP50Xo+aW
44A/G6Ye04od4VVhhpP6oUJe4W7keAH2fvNYIOghOJCWDCleAvvcBDxcoUXWHjK0U+fUAEP3EJbx
HhLq5TMHDKrrEp5kf2RLnwfkBtXod5VaIDMfXkAo2ddx5TRKTkmZPZXVqzJZ6UnniHAs+wOHjcNj
uQFbyBFdHQfx0DYZ9MgL8vyaxocjXvo2S2IhaYv3pX21guFlt0wW8RileaaWIiVgebvVbAy2L5cK
KUvOugQzaF10/mNfEPbms1Z6qpsPxHSe8agIpu4+KBak4gbYIOaTqCNy8Xv7+W10kOtqRtcfZOo7
MlvT8NW8zXNwg+i/biFjn2UkmsCpXC4POhWJrjjacdKXyqMwHluMxgiVlSDvroq+oiCCLVMMHtjS
Z4HpOzjLqXjaWauGtGXdCyta8jNH4MPFs518mBP0K+aVVnwn6E/MudqvqDpRM3bF54/hU1d3b7UE
nEPHoGnmuq437ImD+qVMZ2JVhyw8hchJmltCEV9oPL5kTwzDctFcb49pW1iyefkh84HZUqjM3KQi
4yrhs0+XerMeXXJocgyKzGMAParvkSjwAvrsu6s7IH/zJU8mAcPqIwYwVPRWsTDpOwJP+tE5Xqcm
BESss/IqxrqmQ2+Ag7yJBCzMBy0r8iqI1KXiFI3eZziZ4qXu7Qe3UMUyTRzqHSQO7zarT4E9PI2U
4s3E/qC/130tYRMKjK3bHYa+hlZ7W36VzIQshedxkPW7283p8TmbwSJRq/NfQhDGT1gNUXuS+qYe
xdbT+wEMjsMSJivTpFILMsdUo+WSB6n8LgurDGTYz57TSC1CCaETykgsG60r4Cw5z0dF850AxNge
QXbKTqMhburD9eorb4qECmphHl+e6j4LGZQbqFX9LczDtjt03nhXb3zv3k9RfZ4B20+rZqTVHWm7
hEqMTb9EDydJQnqfZjfqR9hGwWg4N10hu/1Qh1r4+p1FvjkQn4HuiaMJYPOa2vUsOByqXyQ255Hf
beg3HovWnTmfwvCBsy6Mkmokydz60/kgpBxZ4lqGaDLaAX7Yp60cLPf0dgBLO4Vhas8p/IXMyKp2
A4FVplnLUrF2flZllaMtDOYMlEplfoejDFnMaycnHhU7xDtECxe0p+/q8g80IybKMYCQ/g5mRuW7
7bdTLmE2BsjwGT6B52KKic9dN9xn65K+G6BLC0UOdbSCe1uo0DCxI2Wq7JdGLi/7qVHTc97dECo3
y2mQ4QDSwZjK3V+oZc54T+Kf21ZabiqxNnavGkI3KYJpkldFrqh8DTyXXJGdtKtxhhi+E0bOGxYj
h9QKq6eo8QCoAdn8F0rdwZh/oYWbff49BIhkqz9/r/YFQ8orNEak4+AvpS2iCuK1u3t/SHNWvw3U
GJm8QTPKRqWixKJfJA7fwLaUHzEai6488hnF0hl9s+Xba4iUL0FLswY21ACghIJtKf4lTACCOa0k
8D/8W7ff55uL0Z52HLaqtb0lWukiOCJ0UVa+2qX0htfeHHszUI0RZmrBrSdcQVyIR8gEfhCU1SWj
pqVkP+ul9K+8mpV7lcjOsOSxkOJI0HM4v/eIuOzhhbgfgs0vSIngmHhl3J2zgfdDlA69aopjh20w
sR/+7TVx97s5DffFdu0R1/x6wCC+nFiGZ0MCz1/MC16+ziel7Q9vRAJ1ZBaY0Hv7Ld/3WlYQf8b+
ShJFfMPA3aUE4YCeS4aXXJmwReOsJDUTbjmQA3XxTSemj7YjMzNstpj4db5FT18eAK1f2KKyOEPx
1h9AKI+7i2GAyuKynN+ITWuJUmy1ow1OkKQeYlI9MqAc65NFp5LhhgI367AhlR+9drz83jEDW/9S
pqedYi8zCmj/pC71EHct8K0fz/2rSzvphJHcFp8Dpga5lJqQ04ibPMSQ3yER8Zy+k5XPpLv6csjE
NeaIZY0c7EdC750PO7rBYmc5QuwW5+jrzL84VSZs0W0h30Wcg+0C6tpbjbYMtkM9oRIFDy8gMRuU
uFqfWIQ6P6+YOI6eRYMtAyrDfHVavWFX3Gq5S/mHkXSRwlfcaFTehWAPssNnwudQhl9O/LGiWWk3
lMbRJS2yihSGh+9SfEk9160QjhgDGo1eiuMnxadr73bqd9R8o9HULjU/341sDm4n6x31vCuXXpkQ
sUmLcttCh2LXs34m7Ea9347IGzYYsCIiDJmdWerQGVRX5oW3D4HxPOKsdAqUQdALdWNN4LN0twtC
cigwpf+VWAZGXKQeZFRPMtSQJo3RyJNGNDd9XgT2WDNShLkXlrtfMCM9+gs08zMymcaLNOsmaIre
281TalqxQ5EtZJNLO4Q1BjSc8PbbPDzP44ZY2gG+mn7o0e2i5XPaz8zf9hAoH7MNgumPfA/xnUT/
6Uq0DHL7tMxdm2+UriPpuui9GNKjIFAohpOUwPrFuw1ksAr6W0Yy+x/AwKZ+2dNGziweS+ebbUtr
06i3uR9ki7fe38MwYA+FZMAfQETvtEXy2CkLxkK1TeXvsY7f169D+jUmjDPJ5Fr1XsI6zRVGQNbH
iHOUnZT29XQ3axFZYqnfoG0fUP3R0R9qvSSN0wEYzvbcgSGJ3Dw1g/cbemgBzWL2FW6YU1CQ5d4k
THFyVFPmiWcCPd2FXXqJ6X2mx/5fQnaHuRkaMJlrGR/Hpw8oWlA7hSbfcoXq9xfJEWfcE9UGE6fG
nJsc1jLHwCov205930BehFxEZv9A+P6gx5l/hsUKKLV6v8H8/8f6Y6x6Xj8hYMX47n396igeRJvA
6dKJQ3dsYXDsx3uMOP5R3oCEAvtHiRXHvktk8Sc+JhlsZ6O29a1IbfW0tV1jrsuM/1ONLOb/ddt4
3JfnZ50efKbZpTS48Z0DkY6exgeHjRzpUWu/E5RiRfwPrtIip1OIqqoapAgGR1OiR5TRlguPpj1M
TMT9UID+q4EEb0bpScK1Nh7tUPZtS0B1O3kezjzEIhD7wdsY1rMlUjvTTEybyD4vtwEFbv49B0Ua
w6Bf6Q5OiwyGl+bBhRnXgGayT3ogX0FrbtiSAIfx9ns1+nZlK8atQ8TQnC3MlKfkH43S06GcandM
sJJVwMdSqlf42pSetCTWd6G9NUUp4ZJhrURSAVwnHBvvbHrfM9YWHQW6KoyyzFSCxljyVzPOCU71
iQ/d34JBMEghwKFIhzZWh8Pdh/5C7PdQ/LiDebb65I4OWP+8dVsoDnnovzpGrK4qXKOAMYn/R8AY
BUY4S5suYy3J4qKt137yaZW+/+m/fiL4mCUO5Nxggei+kGRx18a7awKBbZyZYgfO8KCGp4noqFhB
HXsj2n8EhhgBWSGl4QrT5swJoQRFq4KjI7UMfOXX9zN9JZFIQ8dB32tV9c7I2pr3k/WINq8lmsDn
OdX5+gOTYqrWnslK/iM9YngzFf7TGikBL5YaWsuB+dCJ3ZahEy9NiMRm/JTD4kY4fcZqaV3G/oIo
HeT1wAr3G2RzLdNRZ7QDZ51QCDUb+0ctgGxxiJgU6Eh1BY1BtMy2qCNKSZlttKRFw48BF53Fa/hx
qL4NpU/DfDdwAaBkJptxnURrc1UXn/hRbM30HH71PONEhXEkSdjJNX1fuJMRhk+yrTd2KaP3fQsN
MzbVztwEYGAFhlq4y5WcDp1E83Nl+fh8r64pg9DKhoZBIyYrqWngh4SSQkzcSezRbsAfbY9XbI5i
2/m974EIExFxTEaBlY3IVck1sM4VCBpx8QB96AIpVbBjhOqwdloIZhLI1fuPWdBZA+/eZVMkalwX
RR119xWoWvd34Mob98mIKpRRfmycm8dkQ/hyHCovubbXs1dGro+QzD8Fz2tMrAmVsNef5w26CwVd
tP4gzH2Yq3knsa2tbNBn0ioSQ+tN1K2rvW0jIRcKVBssJHW4rgmNPYyj4XWqYmj4OQxi8B+cOYQr
0I2Q8jLe8DH5GA5Z1aY4ntmIfQ1LNrht5pRwCBmp17WDhW++8BOfyprHbNW2m/oXqn4q/cKYjhku
Q/zP5akmpLVL2xppRxXfcdX9IkOwizHdUJKMz04FPkQkUNjO50/gMJ0ZzmuT+i/vSg1IniZSv6uY
Sq8bT1DyTJrB61HC3rerRgfSuWAJYFjuIk/pCkhWp26ERBbo63QVTS/NUb5VwHa7RFqCaUwIo8Sc
nN+jb1305rTY5IcWR+mvlTGnw1RHXS709fMAvioRfcVdcX6lFQ9CrJdkkTZRmhdax1GlsT4Fwznl
JmWNRTjGZo/zXXGO8BYyRLSqFq3Uy42PfOzvgdlgd01r1Xak4VjZ/CN0b/+/bm0XYlxszoKudqNE
GfqhESzucPwKbXDRLPRZ4PLqamFuWWtkb6hw6/e2bibtO+a43m0RN7GcTDPnvHn8pQ/lCFHfmsKO
CpbFxcvmW3bqDXJfIGAfJsiWDKPCsPD/Wl5ou8jwMhOzrFtShh5+P2iykY291OQ7wrY79u2rY+2z
/zlbtEPS3j2XFME3KsgEMCh/lIf/6T3K18pqM1Rpaq3AiqAWVL2KrjYOlgWLJr9LNsQIlzHVsnDP
67+SGg0Ca7o0zYz2W6Tae1PGEFeLCYfvXhy+nNBpmkv/YPuEvOLdPHXoNiUEBAP04amx2BUlPLaM
fLkPsfkL4znoNJp+KlmisvosHtluymnGUvDNyXnwmYyWrqyiu18P6H/CdenJHBOoLlo9WC1YY21m
y67ofBMSQYYogZXclP36v03RKmhNY3X5tcATbVdR02Y4Sbp9vUMXnkS8lqqUkTNRs9xI/BTftqNT
OR6I4W5qqmjAX839lpF8ycenPu5oK+FP5lVqOp8zVlulybNQrJ3CXjO17fyPBJxkNoTLwhBXzQwc
2oXhEzbZ15UYiWzwpFLI3nPqLErPgie+txgkBAz7kn9w7m6XYYvLkd2tTimWT+byUn738XMfY3zM
vZ6kIisKrEqXdWfyo5CFZnFYYdCwXaoFJP7I3GcUj9J1MiPXX1DaKbAe1s0DE1nCxOOW+ai0F2Hv
gtGQ8MLQa0BRnflhzSNEar59SKRjDkwcyROzMpx/G8si4JXOym2AFNI2HBlKsNFTUA9mcTYyquDb
rsBAR3oFphhFmw+Br0jhpZDDTYokN1cOhaHTBn+s4dmULlLcH7vSGkDlEiK5+oRLKOvvRobUuj7k
wBholBp70u6YgIEdKgj7f/+YhMrktWRE1TrUFJnwrksIvOUKeNQsXmgADynZY/uoY74/vxs1qWk0
TGTiF/BjWvGv+5U5CqT8GodznifwC27MnXBfNjbdxziRFwQQ+vmnZljUvfeUePlTkzIoysRAsi6g
ZGss8aQuwBl17kYdmtyke77IfYTsQaJZ4DmilO5IuNMMJt0z+QXcVhqSC2JULRDpx8rNrJTz9q+5
Xj/KG5ck00i9YaE2VLxydxXrEQzl+jKpSxsPXIeNZmma2QuPF2L++eN6p3Ksq4bEpOCp0mm76AJZ
lyWMtzYZUOwuMZfNgwERH5AYSA5QJ2s8a4+FDamvz5CA4RX+peufrKDBdVz+8Ee36blNhcOtz7C0
TuGZxt8QNFtfDuRKDMbq35KLVJ++YddHvlaw4MxUshxGs/k5TfHfqOiIw06MaM4qTVwB5sGEKLaA
BlM4daArUKUxxI3ySwa7yojM45oE+0H3eOEpFFu5BcRRr/9ibjm43MmziJfbpb0hATIBToenMuQ7
m1y+tlB7mUTb0ky1aRC6tjDa8FsN1jlOZmrR339dcXXJDm9tFdaEu+eew5zgUyr4YLU2hjoVftzz
pJTiLRQNKfGmztImHBRuPMpSDcKc0zjbxuAc8MjIGnAzPfrttdT8eKb02hL1lXnO3itZZ6aarB6S
wYfLR+SiCA6JnOdPhqI5oIQMMBkjS0hcqLyXeS7VvooK0dQw2vOJBKG24Uo3cltsHd9+AhHw1AUb
OBIbwytUyS+5ECieTjTtzMOLHDYZyFKoN4TKO/5Hf+swUxcWi1vOS2kfqPoAjOgPqEm0yUn1TEPJ
ftdIROCZFOUlYOJ/Ger4Geb+gZEqCFFkidgg89kySA26pgWtc+tTnUtrrVwUuaTNRn4OFu+gDuln
oo3VRYMUZzWpHZals1TnNV5gAfuw0EUp6eG2H3r4ktgMeeuJE8BgeDwQh+MKyYpfz2ODi97zGiBf
AL4//pVa3RRlU1t8rJdgtnFVkOB3o54pbXHheB9V1de9svbscb85rf9t0KZjbdlcUqObsLAZ4I1z
BH2zSGjVKhY32Tv56/5u8ktLGFyMxtr8cmPHIsjR2tht7bskFtzWo3M4X8xvhzIbSeFf7CGS2alS
ZuZC76y2F5Qw3pWwQcOF3P0h9pSydoMW4zcwBHtWa7eqrDX9zW5MnkuaWITBHCBWPoYQUnfVJ9Oq
8uH6s7/dMpqf0rg1VGTZEtCEE8+Q0sOpJYS7tHOK49pgFB5eRRumbEYdT96hpkYt6C/CTOcTJjzU
nJIpfi3nMFOZgn8adEz2ZEPoh/f9Qhgj/QawaxV+XVi8cfE6VG0g31QPBnROlwsUFC1cbQ0H//+c
i266VR7GPG4JO5TQZcbgUH+ZLi8u4S8yo7ezjbo1OlO+SqXvv58BipyVGPGwhxtGu7K3aKHci5Yg
8wn5Au4RQr1u6fG207CCCN/+mD7l5SyXkb6ceSUzf7h7ZvFSDh50Gtv6Obv+tX6ktgWL8ns+323K
Z9abOP42f49ZPeNxqbMaiWFp+wFSZKvv8IQZiATwpS9P/U4HtAPBbBqmh/+L+u4kkZ3naknvVPkG
DWbkR4HWelb5CcrBymUvBiJXyZIQMS3FeDzB1rkQtPIO4Dq589ERBBSgBfA1tet0Jt1sASAueWOm
/s4IZ2dZudHIV7XgOrRAc/z29xsCQIEpGbq+sl2rFtSR3z1CwpUtAfzUf0v/1+nCSwn9jmo+2uT1
iBn2EmLk5Ejw69efJE5zoPp2dw0o+8o4UUpXBQiynfFkiHt+CR5YLWT/306hTNAFl11qSenP7mpk
1xmHN7I7CCXnN5CW34+jhurI6+DHp9Xx/q8Gx7/GDjCVUXzi3tRilzAeUWq7K5JnrtqG6rtQ2Iy/
axfJnkTkWeylJaqu2cRA6cu7EL8tBzq8v6dm7Vw8pse2FJXEtpOA+LX/rD+RRo7KBx+JoNfeN3Im
9x3uU9+66ftDOGUr7yjXMJ2qXnM3fMRIfzatfxnpOuBSSOEuI2oJJ5TEr9C7jEWKig67BzMUoPXq
04FEwykgtNJ68fhu1ttZfsdULSr1amvsYW3oURPmEQPIygOrVg1rltgu3lII1jZJ+lVwULK46BYw
OTjtq+0fGKLmqus/onQ4TIlX3/heeNAQMKUZwmGAQsJYiGuHRL8mQ9poWy3tLttXrjXflJuJURQv
E8ATtC51FcrJFyVks70IeFv1nmMkHdP3TTmm1aYv77fyxmZq3uF23x4dI6ooJTgPbjEZZUPK+oH7
0LKu0sQiWiDtNwdUr2SmMHGxZBeTnr9Wq/btXukBqG0xM58u6qrMCbKCTrjVM5SWQWJNzLSHY/Zs
8HGkPnpXhVU2VEEQ7lGaAJ6u9E9yxUfEpWGDAKk7fNy+tJS1fYRxRYbM9FLU/KITGx5nThRnSGLg
JcsTTaXKVOaU98NULiARaw6hng4hUzdb5xTEQMhzVCAlUVjsDfhh17YsvzyD/ETbmnr/ap0DcG2o
NhUcYypjLA3xZgIEJHN59slRDhIB7cB4OSrSc2DQQhzCE0REI2BD97daCLe7FlpY1Nga0zVNhQkj
h+tKuevP3mwj8wbFKZsPIJgXz6g1+l7ToyCTQdNVhAnQ6WUmxCrGDvm+fIpLBTDxIkOs/kJL7n83
aAcxZwAYq6TaGu8hDlYSLeLSMkin9yVzknr4UBsVr0NyJIEioKlHFbvOwi9sR9BcrQXA0R3UaieY
qK4ktJRxR7lRLtv/WBJguKWwDLvxQazpx4n8MkXMQAryrdEu2W3ZlcyDrkkm9KVLm58myyXd7v0t
SnfZLXI3+ZxrWUkNf3eyPxgvPizpcPYG6nj65S33f8U/x7RI7a4GX0TCUO5jr5kIHJaMG5s3d9dj
NOTAbXAWEZJWrccI0XsQqPu2YJH4TtlpdtpbJTNwDrMCLcinV5yxkE0Oo5mcarfbwZL2HmfdE37q
HSwxPpW2LWh6oLHerbv4s3jyhvAJa2YgNa2wVfRY9TeRF8IhL3m6MDUZ7oFhgrALnRwseku2jSWa
BLkt1zQEZ1Q3aYFbkAaR+e9u9Pd/l2/BvHGZ7udxlbpVe+pFx+FhUIxH2hYFZ4fngqm0GCqU2yyT
G1wcTkJSUSrttBKAYLDFcYtQSfAT6JLFyb6gn5EvUP//J84QwGyZ+f3YO5yxjQJ30O/U+ONLe+MD
WOQZ0AhOSJIhe1NkhpIkgtomnCkUigAZic+zx0M9JEuj//vACJvyEHli636uJUwPKGNpWUBa07tI
W/Oq80QlHq3Kv6ahfTzsXidLlkR6NiHCSueRRyGRaJda3D9Z/j9To6Os2SPWQy85GWyOhOllUSfS
NTTh7stdZU3cMOFDjJqVjk9mcd3KsS5mCuSjROB/WEd7Jh1vI3Q9w3FxuonqbTv5Zf1jGGXswiwz
CCgAcwl3wM4muxyk3MjK7slfGHHlhmbEogoqtQ3UH1mZTBXVjsHNHLU++uodWynOd2IcsYRheF3y
koIzfZWFc6kmGJp7xeJrnFdgjH7AqHG7XrSXu9DRwueUYb+wO4OZMr6idqHbkIq8/wKSQ1svnLMv
JDzV2/o5npY2gJlwTolk9VBoxLbwgDZrU+sft/ixeFCyYtg94FSHlIueG+jKTyUya2opCuVvhEPw
N8EB1WYH1NwHFECD1iAjKEKRDXXCOgRHcwhpOmNk+GUdiVMXNJhgv+73fsFT9c4TwAfiLZgaZxAc
oGvhKJCiIpE6Dr/pJ5VIA1RGRjdSdJdeLPegkC1g/Xr0Jw1vTkszDpowlbdT2dqRNC5b1FaGpif8
2QtSJvsaTrKjtOrSCfRK3G8YnHzB63d8/GxTeCOfoR0b7PiVIwNcuZnMv7iWi4vFx4ozbFWBFjxs
rM3jsFiNeEHEnK51wxDnHilWRGOkOic6Y3n8s7sVqnyCwR3vIPdjMSGMNm0FE+LgwWGidqmb1853
WSNHjPOk+knPqRrfqS3J1wLJNzI4mNzjTEdOHhMJKUS/a1SsDkP7tv0+hMTe8uNgMfUPDjj8QEb1
jf8FjQuNTC1XCO24qNnrcVzo5gCCzVPmbkfeVlrwfWxn76eggv9H+TBXGukVNTsmWCpxFrssSjX/
YmM7X2Mu7e/ikBqY8WHji0VvvQ0738My0ctjDqXjuJ4gEqUiwoUmp9v/1r92Skop/W5qZwGHSmj6
YVrDun8UTdFVO45EbMcTm3WeZ9Ymzj1NYViSxkjISCdpDLVoKjyRpKM4l2N5Oe4R3D916u4pW8WV
UXanYxxs9tFCv/vx6n14qiwx6Ey8XaZn2xyU4RlMClz9DlS+5cW7/prfCz7O9z4FuIWMxCh+D+tP
+wP6x3npWZAY8GNFN8jePrrAaEwSjZjVtZr+A1B1OHAxuN2KQtRH0DHRUrDjlMnE4btjWreG0jsl
S/oRNf3deJgaebUotJB3/j47kjSmTXbSQ3ITxIudqaPhFu/BzgbBmQN3U1WkzssKxO/GxmCX7Xa8
MMKULTyThZNsQ7emt2WWUpM2co+go0kWL2JsYGAm+jxbYGxRWdCTFW90M+ORjMFlfB1nSkoKyaCe
ZVCivtqAAgfs9tXgoJvyNLGSoM4JTC1fDA0K8l/9JcJUFrj1oN7vEOptV03tAX0LP/R+LvjbZOjf
yivze4HNZOR0whf4wMDef8TlRITw3bhdpdEJjzwfEmLdrw8AWQufu2xUowBs2/xiwUbP2x79s7PQ
3aJNeSujon6KtSiCsaWSy6AtAtesdggoMQkqmgiPTxYdDW6C+i2IJSlKXoIPODN9MZVNQn2jdD2v
bhQscM+Ciq4pwEToQVMTByMct6BwMInYMcBZm5H5Ij/Bn2UDzesZ15deAQdbvGtiZ8QpJkI+r2oa
db30UyqH++d5d2lPLF5VsWsjJQhb7vC/PAaFm5QT9yBly/qirTk/xj1W0d1FzQcVyAyVC62Nug5d
4/uThXuH4CcblUiAL/I74ZeBcFzaFaH57/3pS348Jpl4T1TomY9lgeKoPDHxShZ+CbGZF2npfGyo
3UfpRlbxuU3SF59nQ/BfmolL5dQX65EBt7uXA60qisA2TIkpIf1NwnufeNGn5t8YOVPEURcCn8gX
7ZdrccQInl1N393njmxr9W63YJkibPwUEvlyAdPwBEVQ1nzMckUSMW4EHNXjCF489ol6Pr7f0U0A
6cgTy/PGwCuOGzWIjmTweYYyKhdAR4MjxpZrcH7/f5L/kQAiLKRTLmuoiE94mHRDmDaax4U6wTw9
k/LgLuOauvXZuAtpfy7G+SzgzoWaOlkFN/okUhH3TizTh/wwQvEIBJWFQJ18Xy2MMUl9tfVv5zST
xjjDux+SJNId/Q73ZxOfXrXGsQSul2/ALQkVFR4jz7f6blRHlemHfWpkbWFLQQ0DnNZvAnXkjStG
EMHxHiHW2egWE8vmqO2jx7Hrxh9ohdf3EtSf+FOHFkGwfOF0Dn0BgTsogdbQs7EEeofP1KgeEghS
K1Ru9nwJBlLgsc9Hac3YyFgLKNYfjGY6OnSu+JdzQafhpD+2CeZ/CcT+KG/5eo3ZK92F5Z9dilzP
7BpPuK2beyV+rjJcwHM9o8Q8W34dtlwywN/TGXCY6HStOdcoeDT4VyTrEDfvlVHXQwA9eGErL8ju
wOXFtk4Sabyvt+zNUSmavrShu10J7lhYkmhbL5pAWwEbq7y6thwNAA7su+rUS0LHBreRCClhFHu3
TPvJVLW9Lam2n1dyidxRrnLhwSa6RKbGPECi5yvTQM2dbWpwxZFL54CfkhbM5rH+irfLdQ4n2nlC
6xtcKyh/SCsoqKHVRGFaWe8y4DCMmHczpmAPqWVr84mC7KP4Ecf3Lwlg+fEVk6tRttfMA4Mikc1K
XoxD1xpyA21j61bahjhVUXuYFuURwHfDATpquMre3Fs8yvdPW1zs/mQ+p6MoRvBdToKCrd9OIjwm
UXWYW54UGtlKmBNUNaYkeUwXzLJ99H0QNDuI9fc58YfJdV3PVJf/VZycuu13JuN+YdDSUx4WZmYz
LYLxu0a0jpQFW+/IrJ/UHvyTQyYymWf25y7KNNie0TSouLtzPE1etOtR1aaDtOR2I4KoFJpkn309
hFhh9yguaFCyRak2cQTKBvbb4heEpMxockuoue8yfbQJF41e11Eu6swCFSDRNZCotCnUlKjyaO6e
9Do6ZGa51wbAmo+L4Q7rfy9/lD3aDwAX1N77aFhM8Zuj1OE0rHTO4oK6QKIMle4U3VIB1bNKnLqp
OnQA+APvCQMkbRvPFjxF+bcDZJLDdlQnJsAxNZC0gn3+ne/Q1c2aYpqUIJDvfgx6qcX9GimzwffD
NV+CUygJ3PtASOGv14aGz6yuiPfR1gSkMNfzkKsRImYgknt8fUD0uHaJyWVK9rJJj9VWNBdIRJg6
NR2XDmmYPF6mVh0oImuutHbCWFVwBGRGJdbT9viOCpQ6BahvY318PGORp4vwcAy3+zPW8qTGI/WA
6EQ80fLSdTy0iy/S5Vf0AwW+yWXUhdCW3pgjN46LmkdQ0uaSQDSz7715iBhWnmzQcCtsH7GpR+sb
Ukw2GP+xQoQpgrYbgotu5hATtir3qDFq31eWHD0OcCRJTVJ0TD68WtYKK/LatWhxt1f3+KVQafwr
IGqu0CSr3K2huXylQJ5B/Sut9zwUIGvGou6tsXIKuvoM1/dDR2M93GxujjQzSnAwL9iS2dAVFtEn
jXQGS8UhWbDLZ5mUTdpIyQ4sOyyIJeTG2fJM3r3MUc9z+R14Imp8m8PB/rBPedtFQ3jdQOtvOQA4
lq3TENdMYoC+Ey778fOJEiIrves+utMr2/9RZ/nFla0u2zKrIQTyD6fxsLXswYUMi83h6A+dLpTH
5b04fPTJLN4bqPz8xVtxc+WZqYWDR6bp6Zng86qJ0rz0GbG7Cnan4zDgwvdQZpswpydSdKqinJIW
h0YBEENdgNBj3mR8ylWVr2070tc0Sk6Du3SQ2d8/Xa6+B1LhgOIn+X27dN3dmfwKv+PGOuN+lAa8
SyW1UZhjW0h19w3EoNyv63poW4IXSyrEfL5IlHWKhSj02+abNfxACYr97qEgI8B75HljvxvimW/z
4nNtuXvyGQccraVB7lI/SMa989yYQbAicFgq5Ch09ArSTvAskdPx95u5JWrWAp8V+jXlwebPTVnf
yd3dlLJSPIzdpsaYo2+UQRL/VcfM91vUISNWOHEIlKGRNsgt9AzFwVTz8MlFK5rpj+DDPJ/mMJu+
HYpx3h5ElIAA/QA0NzIXVpGH2AEzlBeVlK6pL0G/cTTwViwqmpUg1Q1KTzBdVWXuyYAZqFvMz+U0
4taEtnbGND+p9R0wSxdgTq7RO0MjAYPJ3gdLS0fjSPb6z6eQULg/R1xeMoGygx4YizeAEnCjtf5S
BlG7EMlxdRxPwk/a06lb3U8q5h1f3Kk1Xe0bBv/OwvKp1J1yFvl7p7RAJrZr5eNnhegPmbC/uqVB
pwqV0OeN5nKsZMlMQ2l2A+qjR2rMUhF2idKPvDNCMcfYeVVq4bjXH0Dowjy36GP2BTpHF+Eht0//
/PGBuAaUmWQpHGEHCvAxTGndXJDO9RYBUa86QvG3vyt6TEzR4JRIHRXHBM3Ay7N/4lV4m8drhB9K
Dmz38cRlanzJ8RgfckFOt8rCgKDIbb0Nc/B78HMf345MxFgJXRKSz9nfQLW8Cz6KqiPNQ5ha6y5W
dJO7ev3/5VimGmWuYi/7zpKVjmGrS4HDBcZ/84LA8RBWa3kaE8sRdpZXZ0IMhtR/GJbDCgux918r
J28C7jYMAUDbsSFhrNSZ7dYTJ8lmQyFX8SHl/gEFTgQVsv1H2zS9mErLcrJeA7g0dvr4Sf+3FYZC
BZHoFUJI4ItpKxPAAjz4yW1bfbLHNZQap2LDXWyjfin3oL55lKYAgGTrjMXwvpHV1segLKpGXM9D
OUcwpSHFpDPca2ZyZp17IqyvBFHTEGevbqsbKoQPMQQvoZ7cX86IDwTUy/UmSimldJLBR3PnBnCM
wljdvsTYbOA/tZxU2U0/HUig+uH1Gpe5E5npvCDLOFVZaOpUq+YXDZqSFjmwDR3WSaBVJwHRXWkZ
q14tgmdc8v0dBcUrpKLN7SDvMX65L8WE0570RysUNgjy3zpR6icY7thwleaFbREr3lXazM5Qfgqq
vneKfVl25+UCTrpGJDo5ba6kaADvydvNa321n4YhYZFxi2NkItB7rnTf2uQN+R/HVtQIJZyaSATV
nvh/JMIE5lycYwnC9kbF95XTH6OzSHlj645EQ+ygUd5nlbBaF8Zu6Q4k280dHP6OpYlFWrV+ciFh
Cur2o83i31uI2LmDW6xqKMf4cyRU8nPQAS3kVtXe/4PTOrMkeIiShbIkZkJRcrv6nAQ+jA2b/dDW
l5EnNJi7JilE6PDvw/J9wUh56RwnUJ0TcWuDltPZItUrz/WFuf1K78J/4PWMSfmJqbRDarCzYf4p
cHjFqhQC4Czt0URCZxfA14bL9XC4w2hcQJvK0EKFwcxMchAMiKzaum9h53XgXeimg/h6QfyfQh0r
NusmYQHeQmeMmyXu9NBOqoCMTvXLrhLEjWtIcpPRnn42o1AGdwg/wMkSg5O1QZdzB8huOMu3dZaA
lkiAgpma4KFg4df6KFvFD/S1klffDS4GP7VLQyzWUpHTz2A5/rDT9hZ+BDdLQPhsxDFfw4AuwdUB
Bs83Tr+AI6IQjdloROmRpatHNvCHsSfAHwPRSjB9mj7/tWcoi9+wCUSBbmPeZIBN6LSVPYTNvNWz
RIW1UHmJf+qLfyMi4Yd9/eo83LFoNtDSq7X7S3YmwlMXPSprkPPR1SQgJCeQIeqMfrTTszUHrV/u
O9bgRXMVJC6lIJWn7RQd8GVrZXfOGnS4CFXK25lPtJr6XyHzAlw44ADDZIr54c8RHEIeNVH/Y1bJ
Bl4h7xfoO8v9UDfPiVoac9m1PdaPsVPbeTY603cR7aNK++hpcaRf4Maymftb7xtw1k9GDjgwtYOV
4+nBtyETmu5FtNfljCMKy27rHLNrKWOISzYiZuo8CLBHtqACfDjM2Kt+O8didv8SCnmTFEt/Rldo
a+ixNFXYXBz6gj3+bTQ1bG1OqsNziFkruafH1GB5DGuqRVL6KXlruyJFp3H9fennEn6VmvgwCx9e
Qk+hamhPM+CKIBBnTpTGgIw9jZ8UUxuwWO7AO7TXBTtjW8oOl7+r+f96qb8XN0/rNKNYaiADN13X
x6T4p9SH94UEyYdEFqz3DK9IR64J8aY9QlUDYAbARsF0/Fa89vvMRr1SoJNPWhNnZaGO9x1LXCKR
1KWEs3GzBItwT1O2jMHG//fRyelPmKRnrO51E4zWkE7ierUMSgjQI+URe1CRWBiOYfXIiEuy46NB
GYmKgcgncu434lv8Z6dvfM+u61obcpjkJH3jKEUVQyNTHKh7tgyjdirLXLisVshcGgkVqtc1Vw+c
WDYfMempIBLwm6lBXZ3sU0njwXfPLHNZRU+T3bpXuJ6UaYPir2OmAu+yXZqqiMyv0P8gj+y7GRIU
aQQGUZ/hvjUNnY3JOPJ0UCvMEJk+lsnoFKByixpTLT3gslvHdV8QMF3zo14eK54VlAdlga16DI/F
aDMQj+/bztkUpxd2OOjlv98U9vy2zt/N5STfNCM0RQYz63NCm0b40CX9fSBfKM53qnWpdit/Pg9O
DhoBNxrHCGN53ZrZrPMreY9Kp9rkgwQmhrkJG1Q/f8Wwm0FRU6Q3qn1/QsHOZqWbzFNYUY0Dw5pg
BNx54R4vzDlmRMiX1RFZsSKVNpsKyjBdIpry1Eo+ouNH3Y2X6lF+Bgx5qR2KOT07JX+ckPVxDeGN
Kb6iEU+EG2nMGYcKyAjidPjgw9diBLMSKLTtYsRAlWKe7KKQT4Dq525kOI4OoyunnvXC4jEf9WgE
N5GPWVPRlqHhTWOFz2Y6vAm2yCG17kfdoh/e1cEUZGWKf74NEXXqcrRLHawABWpGt2dUpms2o/hm
8idSxNbE9g2PUwxqG0u4rBPjizOcuh5MNYL2sU8iIpIecIWe5YSd7poURg+yF4J8V9yWA5n1iGAU
YtNdG5FaszZMcnVzl3xLO2vr9FVuQtQwatSiM73s/6dRiWUE9rbtUN15ruoE5R7jGunjGQapayWs
z3bXuVGBsLNHsbAgcC1UvXscrdb92dVsvAe11ZBT0llo01IArwAR66Sc4OOfw+KC53HbAON32Cm4
7nDT2W7yZcJ8KbD8KminAT9ITr+TqFhOvY4WAsUNtzcVf/g9nBkH/4BtYCwB3w5QI5O9aye5D7Db
VqKkx5LtB97vqev1nSpe/id5Q9IZoKacoezfiKZ2IGc+pWS7pBpvcsBG6D4eaAfjRCvZYe3YXzNf
pnnzf+Ey7L+rPppReyn6XxqbWECuNFpFFCHCMHwoSJwEJPOD30DvZnSyxOA11BRF0GgBQdgswPYh
jKkQ2uYrcyTg5Bmi1AhulUeonHU/QEjC6Cmt6tD4EnCghVfhjZIz2DxxvbJfGtFwSISGMTeQdAvn
SZ8MLXR//oWBHIwbTfS451JGfiVr+tUnw8hSyqTHDbrgoy0FIaL+N4ja1Gl1ebGcF0NGvoFwmg9a
9Zv5ZVxAZNdbJTrg6dlgRE67VbWamgncrELp0iV0h2FEuda/W/92TQ6IXI8+YjNtjmLw/m4f7INj
XMDGiHqCFAmyDuA3hAwiH6QeOKVKT4zjhr+HyO8qBYNfR8OGxMHnjfbj4gkDn+Exqkm/fcJie/8E
+rIiHUWmRtynu09ixbO/J1gvt+A4dGwlsYdYS5vDztLi1odTjSoYpt0KuFzyJHVUKOzVfkF0xZpG
ybskrfDrP57hKSa8Xkk2yrKf2CgdyBxlfq/4hr5rOXvAJFrfohosdOd8Lcln8+F7Xu76sJzK/koB
eLCJhOS6+K267sgP7kb+jzbdPNSyIJpVg4i3YNhPJn5+yd3B30Sb//MLsa7QLC29/kBMOkZAwfIE
GnTn3Ns/OB/sHpZysVS3vc2uEAh4fBEI3HkNxqxOiQvcYVPvhLYioYplMcI6i2XRYRea7azQFMSj
TlQ4CU3F9x64WjIoGMyoJhylzBAHjFEKRBMo+dCd1qiXFRiHfHU6HYkZR7vsVmGnI9HIZlQFFhBE
c/HuxkVRVpC9UhxP8PTHqa5prmtKmnsnYIzCAKmikevD1FkRdwFrx6/r3lDkMfx6e/uOmQsN9wsY
wDfgSkrsCUgKrkrdif3wzaskNM7wcy3n6nViNMG0WevjNNy3uNFE4jP326EC+7bcTipu4CJcVq0I
R72LjyverU69TCN/VltEcD3zGGAQVw04BasCSt56NQNjzJ8yEtkVogjABCINWJZUhYiDfQzyP0us
WJbe2jydQJLWj1ki6CO1fWXTaH57w4tQsTDcvRHYZzpbH3+nez5vB4v5ES/z83QWnqUxnv4Z5aZI
vVqAayW3qWgBVbeB3k6/BJYw9JD3HFo37373K309k9Y51BglLkhoDSG9zuby2klRFuy6/L8CQGED
3boTKLlSwg7TPB7sXuLrdp2CIgTv5J31tA4ESptlyH3a5Me0voXUsQ1zJeKp83FsCZSrkb7H/ZJd
BFEqB+JybaojcvGtKVhWSiIcR4sht4r7wje1trgTgxrLtGPi8S83i4NWV2Xp2YbZ2IP4BYNZVz96
SyEcXOaTGXq80lda+7klLlhL0/A/wlkGmXBKeXc65K1IQXatD3YxpeZcRK9zOYa1mtDofkNmBK+1
fIv3w47IIT1SgAIA4Cv+GL+Mt0SMOd3e2AEAIKqDl0r5di6cduRl2snpWEBtu8Re1fJNLiVnu8wu
/KQMbBZJj0CxjZLfu9hWJfrhXr5v83pxPjjhmovf489rojiRMP4wKSklr745E0Vy/cTdwBnki54m
BobB3B1//NQFjNA40dj7XhhC1bBGV9A+SQh+84iu0hYt6kRz//e6Y5anNUeNU1LaXJiJegGBLAYa
9iVjs+Z8Js4sApVxHRuxnEtXfaCb9hq+IvjoZNqzHipBx1bneiRBdHeT+/BEGaeJndT0qcUeENom
5kPokBB0wx1FyZp7naa2PUQEPlFNVzX3nfqvAE2vr5KQ5c4K518Qri9Vpp2BpQKezSIOSSysxatd
85jl958elFknFTfaI84qYD6XRrhg76sJgZx683Ml219P4THVYbdwzFgNVtrq9gug7YmSN4Zcl+Vs
bYCenT6mNGPA9jlx9dYzJwMhWy7VqiQcHbn/qHFvo8fiW3+Kyy+5kw0Q62qgo00rc6zpIV7msVVf
YBJ9fAGcUVtPi70hp9iGr+qfui8by7h7R5sMwC+zPRSsUtvlUyHDeQBNDWL2qmOxcwIJC5jUJUF6
7BYYyp0cUC4qIJoK6W8PG37CvZ1ippR9nBY+NDlK5V98u6okVa7eRRs8JdrIwhIMobuHV84/9W+c
rhNhjlBOj9o4R0xEhb70eNXotYHYyzPGh7/Gu/dMmXSUt3BIrS6W75vS4RE2UPYdnAHs3dbA88fH
GXN0cVLjIKpnGH531o2ZPf/BaudS3FnPIAVuqVidJhlq7cLRNrtA8UT5j//VN984NLPLrPmlJJiE
8Vdo22YzP6cy0XnNNUuIqLkMNWLy4IWinVjDPDh6CghkeH0YwnSHCKhX7AWLu9vvgdt1AQt0GVP8
Rh3mBlGTm6rMROf6yfYMIBxfgOLo9uRTHPujQk5ip6/jQUs1lsCt4KZVH2mnoSOF4fPpmSTFrvfJ
C9Es7v0jNVNiwIzWGHH3A3cwBRdpZ+cmViBz/VTRigLDSAcxdvje4ork+7jxLDk7zb50pbVf6OA6
POrksJ84yQm99sUUwpVwvC6NvSy9cmwY4O9G3QHSRWEpsksrV8ZQ+A0VllU2ZEUpOHOu1XDfDnHd
/jxbhM5ME4Qn0DHxvh4iNFFVbWwHgIhMzBtoHEtEDEwxOSEWZP08CX91zsCDZ2z2QcAcJlL8qrfD
l2mlbsWovfZ3eWIlf7Isc8uXk9byFuEhLIA8ZbzMwDyVNvlrzV/rkce+eWQAEFLsZL9pw9Wiia5P
aRVxYhyBqoG0skOtFExb7DDARwu2ue3+CR+zVkBVikgiJKDRJkF82Hq+LK9cPbFhRT0rTMWmuARG
cfParV566bqoA0AMQ9QrQSH7D4IaEc02UGjo7N2Jpjg1UgtdF96QnnTFD9o2DyVyDNwal3H9Z88c
9e39lh/2uB0NGByWy7W706GJPaqHlzXyx6Rxa8DHJKHTD5EAexlX+P1D1u80WyQXQuZhkCYS2nLR
cbOLzOQPhdgx7MqzI8B/ttTgm5C+madkM/fB9OEkNpenInzn/yHQCA1B1SeUQhFRZteryyuK2pR9
btldTVGHecTHQ7nPOOv6Bm3uKoj35+5rnS4PHg+lfQNHJYgtbhcQRimwjfbh7eTxr7jQfvmlmdsf
BNdjHlW/8c/mdCm3SPtKn9lw+X9Q+U7TzVir1keEYg/pf+uHFJxsrHs4AvvxiYmNoKfbqRKVWJiT
tibAf4LnHb+IUYAg79lUK5uhMJXYP+huZuCeqlDEvLV9k5HBceukXp1uao9pZeuXJZWtE2BUKmNT
FtKkFwvfciJo9TISOty+vtXlWgAca63w65SLBD5xQYCsnVfql8nzETW1pTKMtGGANJdt7l/F3KB0
QR4CIRGrNXcTJTAX3hs4lGDQwo5PO0DUH0iwc8YgBOh2eFlOKljJTaxVGrARRmPAvvX+iFkXVYkH
KhDBNzYf7itE0Cc74CJPyYAHJcMj+dk6GEsrMZY17rKWxQHSge2ofDEGSUgB96lyAjAwjENnD62z
yp3+0Alw32djizIqmelWN6jPQtzSLyxmOzUY9kC0PvcQ2ch/DdCnDbjq+38Jghc/CwvaLvw2tP4s
uVGSxUKy4fcAfY9/Bzmo2SeuKoQCNwrdfsrMPRPmFTo9o0Gp9VcMAVAfap78+H0NXBnWGpTzzbYm
WSaTzO6YlN82ntOdFcpDq8HdGnqxEBQzGSyiNtdlLljfSief+uPi7D/2NGH9QfiEN5+DxIripsPD
TfF2ISpXSJiak4fwhWhVcS44dyY+cevGA33kBDpka1eQYzCVqqntdepf6VGbgIBaaca0sCPqOuZR
gAugiS9GT43IYi6lIUBUrhZjfD6m25EUczsQF+SZ+F+eq+V9nH+ijyrXSxaywuCUN7UazSxKo3Me
zflGV0wlNHAh9mpy0zAEa63PIO6/MeBbDRiYpH2ryfTy0BX5Vwi3m4cgskFlyxbwCr/dl6qV4dbz
ENPBxw5EbRj4zAWWlLyPbFpH0lkdmG7RtKpPe/pe6ziFH0lOB92EhoSib4MrBQnlc1ArTsSe5YfR
MkiePCck5CuIqKZ1JJlXDa4CGZrXPEHvGk4I1lvhvy1gVV8tqTunOWASayE1NTkLFv39Qk9m8/pl
ZNRrWg5YA8GTkZBTocSE4Su9Dj9uWsgg9lPzPSMP3VuXZlhn97Zx5Z/JZw2RnW5ahuI89Fm5K9/u
jAcrsyvcJbFO7tludYfmrwBcFLvwwkXGvzaPIL4HIze2WtojKH3nd/neXzkTQ1z8jIytfZ/SN53x
xVEGZZu0mAQ3+CaeVWSwtEURCZFuCjZnQBeAj/bck56NRb16Y7wyHpmfOvU6oSTqR7lv4ZabLT3/
Q0PRzV7w8rRedOmeGTBJm4uylKvOg6BvoWXU2tWAC4+OngOBcAkFbPYOXJATtbb0EecmMbzGFgN7
dBgHxF59b2VrVEmGmAzYgWUwiEYfKOdVIoCr4CtR9RUWOjGxhzqDngylP9R4Eq5J1E+xv4eq8xvI
DDjVRIYybL2lrpK94TWETMNBPqXUVTk/Zj6ARbURwLSQ2fUl6Hp+2W+1yzWp9hjhbDzq2shSVxo/
O6405mmgi7hf0CigBlfMaN0NN33DsC5HEobW/eghCUKA670cgt1mTn07xyd0vRbCHEcPQCLFA86i
uxRXT4lb2rOO6xWkJm1YO3mgbA3UGdDIp6u3IqEMIC0aqfenUg/n3/NZWcfcs49XYBRgnvZ5Y+9F
bcnJ8LclkKtiPD0bjHnsJhn2+a7Lyvciu/yLkXB29CDxOfrqPQARF1q6eHZJ5V1a+uAStSNx9KP6
9G3k28Q0AYueyyzqZYj7Nd1irOh9VZiVx4s/34oAWGNkU1jJU0ISOb6m42MUrJCNEABS1zhsXQhB
lYMRuLkuNqH+HgCSVJQl6eEHzA/5HENnDOSn95s4ZAKWQg29Q0tih4mx75T1GFkP9Ym/IiD+bB4i
uAL0zm6YcQmVoTKzrMjfgtTWfm3v3t0ICz+MgrJNXX5Ioel2f6F9LS41ANB1TVuEq4Udav9oyg5z
PZKGf9pIV4rbLca6UKrq1nKXPcV9p3E3QHuaKJglz3zbm2WoyuUO0U5W1K3LNkKnmM0yRJNCQcYl
fu15dpTtdtfweVeztq8kS4VXPHRmzjwcvf7fTO+5Jf4MQV+y9pVqY1e+SxNXuIcdOvg1VFgYzggi
w/DWyvowsRMa7o9R/9fUGrlqzHj5TvHhU+FRWPe0pAiK/wmefaHVGb7K18SwmY1nNO0N3SadPoxw
g0/TGO5gVt5wPl105ElJHxDAsqh9onWmJogmLFYS7hLVHPvAVXCbvzghOaE5uOg9zfjff9A1JqgM
wsDOiAkrS+6BtikQ/7yxcavpUs3bg1HOOh8MZS0JPutMxwrX8t8VA3UVrzUweu7fHq6yU3D4VNoy
IX6T4cUTNq/SDoVVfdYj0gDDdhy6J1P1Xekgr21ZCqXRf6hqXanOfg/WS0DEu8S0/wxhYg9TvWjZ
nw4IVuxzA2GU0BgRUmKu0JuS3prcqo4mTJ4WfPe3Qj8E2d1pTOlylje38lBvTqqX3KPM8+IntOsS
w28HaP00s2RlH/IPz6l2j23huSIG6m7sACqufO3Rreete7Q4S6buTckVpjgcwSblQ8d2r3Hschpy
Zh4kcvtXlpR9X8VCYHUUbfT/oObVIHP7fs9oP3VULD5Y4KP0THpvollZvP8BJ7WdebkXmdFCR5fg
vaufFq4g1SdoDCUjIZRWLr3UioysHQK3k8HgmPu9NPPdiF1V4CTKLkYVEYPiBWXN0YdJEYMfDxwz
rIdhBXbsJ1ByXge+sWQuMb3dltYlLQGkWPSu4KTmxBcWTaasFVMK+im3RUmU1gxRpY1Yf4xeHSng
h25a3kZgkOdDODi1MZJxuAHOeg0fQxfON4dCLuZOLhAb/SVCKlMO6lgupqdUry2HLtVBIpBsJ3DL
2QN7kQkaqZVHZYRBMmH8VvFjw4fqTtRfFQ/9KVdNDDN82qWcBZFYvxQDEHFJwbXZ/03jZu6hnHIn
EfTOeeUPgQ0wv2lTUM/lH5znAE566VJ3kZOR7pU12NF9rMHA7tvxbrtocjvSxeuIw35G4kXKIRUK
bgBsZ97OZkjshJsu/4tK479Fuv7QA0q2c7snbDR1TuBQgg+Pai3XV6n/tXfdk4/usmxFXn+8H8f3
w3NI2NlSqlVprGfVy9dnyaD+cvbOSUITN/YKCm/L/PnL1kAfySR/HXm1LVqR68ihGtIgdJiS3e7c
BFN4CTGz0YfUSyfKJetbiYcQUQvkqmelJIgQiOK69He2gISN5Sr6VVt1rSNRvuaPUUoQ6C3saB9K
H9ufdC6xSNoXRPuxRyfgnHfBGis47afI8zqddjkDA12//GamU0N9DRxxgcWw0rGFSsUnE1bsvZ5H
Zio+XifJjfys0nktN/LNjgxXydyoD7kclRx+/NMnQnztoUDCa1VUyh+08FJmh1m/QpMhbAjGLLge
6OgW7N+D8At2imvZYfjmWsOBvD0PAfuWh3KT8BmCru1NpQwBDfvFRhDivYqz3h7By3c2nhI3+umg
Gz/bwFL56IpgosrHIWf/2LF6iGHduEJeKEXMZ3/ms8KpOks1nXjhwIkTY7or6+nnF0earW5OY/lo
igV0VFt87/qzifEFj7Ql5T2H7rY/RiRNGVq7CxVtqBOVRxe1UpPY1Rf+PYRNDBATJ7gd3M09TFml
kEnx/jP62DGA47s0fDpS1bFO8l7nQxnlHC3nJT1S+zMHXzFSyS0ZIXE5TfKK2q1RpjkA6+IuPr/u
047KeFmPdx9SNY9YLBWK79sLGSOAjdkmlWqQYqrLf6K2dA3TcS8kEsZgA/GBRfx9rzefFjryShtU
eUV6tcz+iU+WtMBvB+0spdK5e2qsu8/QGgHvwAiZVyDuiODcB7uvXJr6s2DNEABEpTKcubvG4qrQ
eATsvud5Dh19bgj2HSlNlqKMQvZvZYH3SZkz+bar45uEWnEfArPs49zxG3gzWGsq5u3vDFi2W/CM
Lx+wDFiXWKok3JqLhleJlRv0gkNiyAcuywRoqFCsbEYAvneMEcXsF4gzyokSGPNOzXLVvJo6VQ2A
DM56s9O+QtYQFsgcM7hSMTC/8lXsiRFrHN/9ja7EYXTfAGS9eZV37Byb4oCXH+EBSxhwsBAUPFeA
uJoEm/MIZRxSNhiq5JgLLMX1rU7HGX46PvMc3GjSqoKzLwFqKc6nbJy5rzWCPOFzUWfOKBWVaGFh
1zpwoEHABua23BwqTnxFAAWCRcTR1KUzSmJymhPgUdAJBcCIkNtpk7Idk4oOmUcQdRqeOtTGgoru
eaZdX4oLI+yF99hPsNXbvv6whficH5uz6KbIlCURtGitZv8e68Hd5BnfMs7TZjlQn/fumRjuaOO/
sXCuYyj0MI2+AX2S9dsongNQNWWr8274xSo1bipEfNu23MAehmtXJ6Ei+zlxosCz5CNJxvM8bett
IlyPH4XmCTZdPnx1366Ls4l7q604eeyh8zrRWl1oV4ZMLbliAP/7vpWut/IQkZTGaLEkPuP0woKC
X3W9bfJdGnMqbtj7iJQs0tmaOIYKLnKQfMh5atXkwATjRcb90hDXXsmBuzGzD/NJ2ZUOpyBmuY8u
rB+0z0iWFdcoA9mwPFJmbj6W/IPvjRPLVcdVpLKAM182k04JhaY0U/p/HyTEMaqnSMsBSXKxzQQd
smoGeTLiTxVRdfPdtq0Uq47XHPDp2LVdw402Z+eD8xt9b2+xHKKMfVKkrZZisNIt/m7+5Id0bepw
0NRWF/AM7XzcpsH/JM1xxgQVpOpKVTFOZAPN16N6Utbe/EXhh6juBXKeOLlJpuHSewZy2f4YA0El
hSIgTpB56Ks0kVvqntd8jFWoy8nZRe3J3yRMYmRI16Rj0iNAszctgXsxLosYmr0ADsDJEecZTyHJ
mu3z18tCu2OemOTpYwC+gELxVuiMxb3VhyjzEi9qDkGHU3YNPY2P4oyyvspbGc/5WdAJYTL0GNLd
nClVFcLYfZz5snP4Tekd4YtmwIIcaXV98aT5LEl0bWS6WLidTDlFtoKMDpXtySUexI0aCSlpdJpd
eaqjaLBCSsbVDRVOG3h6zgv4R4kbDmbjLaRPGJxOAMx4WFvfQPxRpvamp+1Pd4u9rPV28yju2zyD
3CTNRT3uQ7REd/NaOKkzTYrSMQqQfXNL8OKWtkaj2bL1a7IeI1Y9lylbgOEoFxCoXNlajOULhOJq
oZeyYcNg6ryPFFT7rPu2MLljfd2FPQx8mJRVwsfYHAno1SjtfNRpTd+nu9ov20fZlWkSuKMg+Apm
H1Q5e42M5jbciXH2LNZpUyU1ykk3KkJYbXuQbZrOyLw59+lcOTAZECLpIvK253QL3Ks6lWXxnbA0
e1/Ajgk3ip7tcEeZGGNBQLRiyXDKl2e3fyIiIEbtUYnmLVX+14nSolUTx5DFM93NeRYtYj9vL+YE
93q+c/c7m0Z8pxtQrJIGubdChazSMslkt6PEFC7Bj97ONFxlrXmzpEGVx1yctNl2aEsq7ZApG5nu
vAWIuRBQuzdgSTfZ06/zjaW2gX0PQnaeYiZhbYdHp7uM3t2G/pJc3raXsXvDbUc6spY2oS/EnVII
O9KbWHcp5EgcsIe9cou2chYBI9b2S7XsfvunO5maamEYJ7Wn8wSi3P7fCZhsncfgVm8T3zeCJSXp
b3ymcf8MhDHRmDBOEbBPFeUTlgyZc5nIeScL3mbPvy87zen6NKzuW7x+CCYQ2+rYnva5I3WQuMZI
Ct9hBiiqzK5hMapGF1SRZ6mQH41WuMo0/3i+teSbxOajo5v7nCpZgUtvagLRxTmQvBOnf8sk/IPL
oWclbdfS2fX0VwC2Yas5C/+MBWvcS00dC9gLLl/MelT38HKnrdF0jp5EcGfmIObXM6iRlGp7Ow1m
BVWHq4X5D6gFNCaH/Gw6/p24mRHtmzhri69iVMD72VbGzwcQk7nP97mfLSPNkoe+Pow2NyBHXxFb
c/R/wJdUDHNs1R2d5I+Y1YWW1IIV6nY+1SqGefmBIBLeennzjMtWsl2vgPPxC8as/cPND8qC836Q
FuPeM0Nxl62lvU9SZnz7F9B2J4f7d3Yr1EBIVNuxp7vq09h2zlewapqTHkrB4hq7w1k1lbkgPLfk
dv/DAJM2/882QT+bsW9zxiteZPiPPSryTI0c7UBlhu5O9K49TsrVcYkMM0tLgt+FzYCdDVDRSnDM
j5197N5zsel6XJt981ZU1/LCRitQl7HoDVRlheaCeoq/WjrmLYoaNfFtgPmjYaC30Fce6PdFXS3s
lvrO9NB//rlp7y83cra7uOKSAtXDMbtY9iIshcyDw1wdxFnq6dsFU/Rr71Ldhiif/NYGPwYcxWCQ
8dHkGXlq1YrdGGNz11ggEd3qnFOzQ5fJfIj2l4q9OLlRj2nPu6Mh0I2YUGbU6Khf6mZEeTWVu996
HEFkZoMsLNs8OoaPidgzl9NxOpXNTAJjRvrRohPCnciBuJX9rzPInnS3IYOFOpekU5qvQ6Q6ciAM
p3GHDBYYtpBDqH+pO+UgEH4ragdD5WTdjUIVrG4t2KZc17WoMSo9HFbb6jOOlhH1R1FER0R8hXVf
dHDjb9JrJFHcRXJKp+iTGDv1/Z6thlmy8kzb6qDAmugTiULhns73sRCKCKCXtGdu/am7z56zvmSX
H+L3E1nIWD4whbjMV0aUboIiiIzB82oXg9k4qUSTpfT8ZAV1/OJLiKOIg8c48oq3YE29xb/GSHP/
riiwVKLcRY1nqeYfHQT06CBHdgPicTJkM4pBfO99j+icQL22D2FtB2D9zCJjw7lO+1nSfQyE11KQ
1YfaYMsuaeTCnHrtavnn/n+iIiW4MC5eIWCQm21l/qb2S/yh2y22g+/h0OGKHa0IuwQzeXVisS0n
N3sMRiEjQR8ii+bdcfwKDxmuFj4hkmRUkcyqyyAL3nv2LyIhGXddhtI9dVz6WyBXvpjkla9s8oRu
4PnCwqkqpG8OE2C9W9ir7fxVlk9grXotZ4o/QWtEcVs6uWeA8Zsdl8c/eNeyUnv05ls+6R8AS4Jz
2KgZpgCH5MrU1xm2bMDSv7p6YjcuTq6TRtrJYJeC+AZouJzTxPOv/5HLVtHUOb0F3q82L5dI4Mdz
U2m5xUQZyFUlFJj1yAzSUGURjeJ3OdO4NM3yp+clPhNQv6DGCaSW2s6uS3ydvlrm7WKZQZDVBI0j
QjeJo5kLwCI+Ohtt4iLDD+9EPPTBRcAvZE4oOErWPnNWuFE8+R8q1l43sfwubt91AITv9x5/ryBO
OqF/IMOpmjyBQWUF2IXdQ9Nea/zuPqsJlQq7tlWMVUqATWkUBn+LjpeKFPywo9xK13who5VTHYEv
sODgj5muqvJfgHaZuyqqzurn14l5uC8ByW5j2+Hwr+R/u7abERaO6J9HT0uqGrIwjZtG/jsjLOlL
qEULqdboSzxu1eUR6SdsCZgW50exfMZ1cza4fyHtJlKN5RF+OGEY+lzU6MHvRxkvfhZq7zwohVk/
WuWyAEao8jlK+flletge2mhFmv726xPS8pAc90C/pLsnN22KK0JVSkGKvQ6UiKGA0hjfSGVG9Jd2
0oFtAMQjB0eXOu+lky1S+AeGBVLktmU59XBOTBBouJ5N5+crXlwLP9axO6vshDn6WmjB9zoI9ckr
kFoyCtAvB4SfGy9/OpOM+cHPvXJwebQNF87gt+GSdWkFqVgHDQCJBwkUYSgiiTGXD8yrd1IspQ4P
fLkdtrqUxAppDIhTkFS+vfzpltfNOVyeS4LJP9wGNcHW9H30onVx7GjZMlHFFtk4GxoCIg/0OeDD
lXiR0az2B5KsnlV6/xp7Z46V21xAO7d5ZC+y2fV53mpbyTsi1Bfsd+drf0azglGLtRPY6VL1f7aB
+Nror0+WMbjBngxLOMCpKZh8v7pOQRzsxC1vLGwP1GXSO4qBBcNHvl+JSg1oy4FGGycLe1le8Qd/
oz+L0zZwJTs1zb6IBS7FY8zT4rdbURjiRDlz1ghQiCU2AEQDEy3JXRmWuLtv5YumOjaI/A4/NNpw
or95P+6hfQIoVqKlMEOQGth0T+btZ5Lpz2HBYcAXTh0U4wTweCBUfS6aC8rMCCrLD9G6cG/BlkO9
71aKCzOQCB1L11YrKLiGnkyaORRBs2IA9DVTL00ND8mZUP6fUgKBNLSJPzNw1Hw6QqKxmybRC+xj
Q4NGHVNx+7S4dbxf6gKgDQy+7wqLHY+ZcLBdj99t0ZC5uijiPpwsW7ASv6XFgb3fHjBqnXwPI5IA
QcAKVzbWJIrqXvuOdcsp4AQpkzlTyFzM/ZTnW0p5jaZ9M6gD5lPzyTgQ2+tV7z2gV+U2SNa6Fves
Du2Vmw+hYpwsmpUVGVMf0RP3PsDaEeOBzbCzKwT8VcIUlnhyVaC+nvdJWiVNd2pLz1v9abOxNsaP
7pK1ubQQdaZhRiryrAhG+YIVvlhMa+aU6RFx16Y30BxMlXr3w2Pac1jSJf0GO4TqydH3KCd9RqAO
9AF58p2J1X5R6oxL8vj7QESTFJkrBjDGe08mZx10Ju4D/OT/OhQY/D8t69bneg4nlTXC8Kt2PKY/
uRIQ6uEiQFD9w9IxHm0scZXZRMJw8GOO9BTxL/mQk5wmGE/07M+6HBh78ZuvUqvD3iyXy2e2azeG
YXTxY14IBsMxIL3+S4XajKJGB8ZbDEM676Dgk9rucXq1HpipxeOCMXJYYx1T4HRKzHzh3Ofqkwr6
2CdjcmhUFn/IN50InY1MuENbflrnnAO+c0PAqbbJIolXlGoBwfpzKGcLtObks5O8Zt/eONihc6x5
ricnJ1cjqJ1yRADikeTLtfj4QwwsJiQRExZ8bBqBVgdsphWUjq28dP7hKsvAnT1AWTOS5cP8AIo5
35LJpYqvuCrGuXPIrfmkdkdpCYyUIDxNYpCoQ6RaDLlD5BFlfiz0DoUYjXCzjTLgkQpFBf7RXQiQ
NJErrqlM2A88DlXHP9PCkoJsHBu62k9C553L/v4ZzmmUh/HViIL3Xu+z9VSYA5mtDMf5cgs6VYOn
+cF+eHwAKRKrFlQ/N4cmY3bFSPTRVUSqGMuGFf9XMk6Bw2IGer/UnAnvHdvaWZ2MtaKJBkK/7vGs
LtCJsjP4Yqr/+pUUfJ66qGx1Ttn3Y2KqLo6jZlP5Tn7SJ5WrkjhDA6k7wEbBah4k19IX0fRudM5w
mjbsXjClrbskdBB/59/EARYplHycqkSB38dwfUda9qdA9QUFTX8dcZjkW4e/pi+Tqol45ZWMXddN
P3jRIkqNC+rm8fczzYk5Z87xt5Oofc99stpo/soHWMom8IKoAxWBl1Xth0pGr+wPKK55MrQiuF6P
7L37f3vTNFB1QiGs1usvy5fWkr0u7Aiqsc6fOeA2T3FfjT19jYk0meYTYsNnCs2bdtmGuHcNyuTI
a/qg9MHjYl95ytxUfk9O/WXYy/lJoOQl5vvTU1t2ga6ndOndWIoanKSY44DT5lblSyBNb8fKcr60
hSabSQK65vqC2MOmN4E2NCqySG2x3mK0DKqM+/JTfdL8hWYbYKGVGFryKAy3GZB7ftG1RTNM2ZGK
PSRhtI021wWJu5ZTBI2x3PewhkoxRjQeKfZArHHZBF6M03Ly6stgzUCAHGlQVEf58yxoxjvc+loq
1GXVPzgna9ruYoutD/m8cz7N0UbuNEUHgivoGVEePb0v3h2XBEnoGl6Btgeku2otXknSTY7K+4iw
My78qEomHH7K1rFteUyOJIbGckFbtebiwCepuB6yXUECYUuw9aUXSPW9GR/5tcdH6c0r6cnXjZEO
tD0Man//jP2H/Xlq7LPGhYkA4mboK2puLKPOOkEbP9O+ODNwEcvFtpW6Fl+WdmHB0o8pfIGSPjHn
wYfqHyaxHnpVyhiEb5PPGUZfdVORUR9CWozyKvZ5hrPLhS49wQ/28aICab6E3wL2ZVZKxe6ZaRNd
nOXU9rmj/heDjrCryj0md+RZ9qrOVa0YZ5NJcHu/UZxAoFi4h6Q/Ip5Mx8LqWZ5wLW5gxiFV7sXw
fD5DsxXl1LBcocpZjp4QXbjivnKvXEP1QXb16lmMeorrwHIDe1p/sQwypXHPWxDPlqYeQnOwtu6d
1k/e7066pPtMKrif7Nq2J/5vXQEIl9n+20RGtrsZ6q80sMuv1N781gM/5de08gOcnxauVX45MYIr
CkDrRN/I3OBU2jtcSy3QTPB+cwZEThTQJkZNRGN0rbv35UZ+6NP+p5iUgJa1ubHI09IHobPWRj3+
pcLKZZEJrRVE1EfZkCPgl6u/BYYPH9CE1650+BRLFp4ifdV85OPREoRJUFWv8Q/Ycqv6aiy+iqRL
sqeNVVgEr3vWvLVWzoNvrgr8N9WhbTkqdPXCEj3rQI+UD0Vu0qyXtI19ZxM/qx4/FqxAIZwfZI6t
Dn0dNp4SABw36h9SttFGZCMG4ovLBz9a/dgmI3VfiwpCdS/nmFNo567jpBZCs/fWON8WWg13Zm/b
cMrin833nwAPGtwc8NbLA1z8t3s0dhgSZlBV4wbI3KE1gCwcVjNabhvNw+XXDSQ/O92GtrmJ1NVv
I1leK9RIBZHqd9D/SgDEWQCWhtr/3MWXFNlJUX+SjMTJgs9X2q8lAXX6DR5BokZfkTVBBqFwPkft
MvTXYijPQxJbyDEaaAx0C4RnD7HLh+6i86J2woUJSBsLN8LOjBBFoVK2VnG0E1iFM8sdol4Nu9qj
mSSW/cJRFAGCMNC7MCOfkwju5wtMYfGIr/KUxsyC/tXNb9fNEAUI9X+v+3l9/n+XF+LMEiAUs3EH
91OOLaAZ8GkFZHgAVfD6aPbJ2AACK5N3C2e1Mld56Zk46gYtAK++dHyeVAmXzBz5hKmH/1fPVmPb
Evs6yKP3buNRO18TA7WXxjTArDzDXG4DKTeIwLuDg6tq9Ig/R6SE4wAbiPDnxe4vcySD4ZaJdJGk
SL8BbdXXcM2iW74JAviwHWZYi2UuKDphrNFbVxatXqfaO9aNFQvRrzOkB6jIXiOdg1B7B3Q2XEek
I2WjK0rAdg1H2g+W5tcC4HNTOHlVUog/X42HA1SB9v3lFa/YR4tcmCFWuXiWOhZ1wKn6qwgsxjC0
lqcvo02J82P5ipgpUcUsjCpSOrhHX4RHLnIYPQNIj3zW9kevrIG0lYltiQBzILqe/sBoAlXsjEOA
UXCrmj+eWjzsIzl4mLVncxbZ+HTgZM0SgPVR/XTLDwsq5LQQ1XDO+/RECenLH2lZMNsyYYwwAsYG
MWg6uU6FZKRgH0BYzHskdy4X0j4w+RdIFg5TuHIxIUFOuiky+iF9kzgOspKR9ODX7XQw715PfIEd
6QP6dPQny75PGIFb+JasRWlGaqzd0M7XTf4Gg9wvylLXCHMjQvgndTwQrawBa3U1lf8aXJVGGcH8
S1Snl5DdO996UIqyEBT9alQj7qA9GznRomNjA2eildabFa0BbNQB9Gzwcon9LgMfbq0ev7mm/DV2
3JTAjmqGZa4UfwVy5GEXs8SEXkjExWoWWq+VPUlmBG+YbI/hgGg0B9qxwPUL/VL2YCfuclh811rz
UcOWJdGuZaCgxEv/50NF3/xRge7ldO09lGU6tKocrtAzB1JkRKP4pymgmPWQln02uXEeUdiwwctD
v0TlflzPrbi/jtvTFZNUjxYvQwbKHL6+uHuzOX6qd/HFFzMjqFdtDq1antvmGDF0buhOxSfcuEGw
t7dmB6hCN7tw4uSBWeRE9fIW0pqlKsw2a2rgn3yY5zio2o1Z8IVkRV/5Txix0dzbOvWtbRx8tzSr
aPBvPkjFvcLFFcnnnMuJ6Q+knyVoYwu/Gu6H+3L7WXZKHLOlUfXiTYd0WrOut8jSNKZwSsX30o3x
upZwvj/Sk65fxER69bMgPGZSV7OGI4mH0rHu9vvab/2By8PHOzti5jSqQaq3o42mb412Q3XJSE6t
GBb3/R7302tG8+JsjtXspGVThgR+OQVzWpi7kAEtvoMEdf9LajnCQTaH+nLADOyH7rqwWs1bU0kW
eEqcsJyePFo6IgcrCoVZrU8g+Fw2nST5LHEZxrl4N2qOiWEPk7xhLChRFVDARv6bth00qNY0f+tF
mUzNVTi4VIqFcxbGSvFx0OC9ZUlUSrMck9WPaiB58uGUbTjOGNcH+ySgvIXWHSjrfGBZn5xnJz4z
VqAtdtJVRk72J4TTr4vp9g7fUINCeHMmOWwfKE4os0TVg+BR54L2X9RXctEM/qx2wigZ1w1bheA7
poWLKAtQVuLgjmPmI5w/3zG5MWkkxcEBahuYaPIXpAC/sN/zQrJnLZ+938pUNki9Ozx9tghfXlwG
IBA/tDVaiZcDBX7Xu4r9ospdpD/s80g5rWdg2C4r7g4HnldtwsFzK5k83exCNDdKv40yjmWckKw3
ZFdIAjQT33Qeqwt7f2Htu5y0NQKe3QV9TfZVyx9oDmzoEsSWvcemsoLLUEjQrMKQzzWhwQQElRU4
w2ekhxjngd22VGggfm9KK9QkG9id53jJmHlRHEXUt5quSJ02TavDyi/+qK9yly5rNUEmY/9ccHFg
AhIpE92TZgEcrUZ6LXxCwGH2Sw4FiTtklCE+okzoUrvID1Rpsrpv00uTihI53qzWaP2MYj0EDKn9
CuPpPhEsxUbMRxyXz2scuAnBeH392yftTAXPUZIEwkTWy56V7WTMamXUP70JC5/rDG4PLf6zhe4D
gjCFaSmjVsTI0FnywrK+uGIX1Px0Qwk/5pjuA35/bZ5V3EcIdIo6gaBcn2gSOx7QMz7JLAJFvIMl
u3Vw31BIHXyJgBqmx/xeDDk5Km/YrcQFlTwvgr3FAmNoihSR7fENxuOOOHB9X1wsh8bEspyqfUBJ
RZYl3TwVUcX+PrwUKtU5Qc851hDdNpMifIO9lbNXjsaO+NwUliaLyjpn9sXviZyNVZC8pnLjm45q
p728wjzuOkkB/1qQx7Im9Qp9obNEAqC32z7EaoPrZowkcFg2KKlANFWiazFcIbfu0o5vNMZR/M8O
b9XpaxeoM1UXJji8OfWOImaJZuMqZn3A3b/a8DxTJ5jGfcjamraL/D/HApAu1NHZWxPAKtz770qb
J0P8uzrm+H2XiGadTFAN+1DZqRcdrZL6f+n5wPboOxHcHMhzu6vqYx5BiIP1pofy196wrzKVyrqc
zBITLznwNWxPlhcDSDFtoSEnsdyz8EjfriTl4L/6ADZjDuJeBhwn6jtWh7THAfFxW1m1CN2rtjLw
F1vk+navsCJqt2BhkI7BwkHByFijT5nYivAd1URVhKmNgKBkk3xkccKGjaxbGeLcdTjL0RwThrim
PnStZVBv5Uj/l1CMeE/ezD4lzcwG/sNFg1h7rBQNiTsyqZ0LTSrKIrYIep5TcEQqvLvIFLWO4RM3
3fclHhkdFb+gEtIY8mQ7u5KNgehQcls1vCwBO68Czj8Bj9U8fJQ6LoL+u8hZY2Ry+FveuL8HGcu8
DnmSUJi4/IeqLX+avXBMw6CTTU9wbNLuLkrtKZPWxfApQ/a0kgjxSpbAB0gudcm8rX7L0pXXGdgj
LVARIfAeGbExOPGKowCYPc4wN+OFKA9wRe5f6Z4/edMdN8rlqmH4oPSCuUB0uCRTQnxngMS1iL2M
hY/OZa9fY8ClJ6hzH0iCYxzc9okXZv2tEQbhz1E0vMPthlADIAR5OJPch7A4JXryX9Y2oEN1CWNb
vrASuPOwnlUYjSP3OOmxCzOgfv4YTVeHHpPudzkoq97vvtHyu3RRlFVn0w84k0KVOJ+ct1tgP3dF
rzZAsHnp4q7Hx/nOFTCOEWkyVB20MLvvKPwECDXDfNirGlLxCFHWkh6HcbXpZup3Cow6gbN2gfrx
xSndju5L9qbmuKo4DJ8WK3laj3Qoz/9QvxCqXvVjRCvxROdAEJ12STxWdEYvYzIquOfIE8ZJDrYs
Arz7NKlQSvNSE9Q0dOexCDA7oePM3sCulvUUVbSQXL59ekBnJAZPS0dumo0g+kGgut/T0vFDZ0Fj
ofSipolrIXO3+OjT0LU17QW8cgEZYxR4i+PxqcpS1FmGVMP1GBYP/3p1yetz+arijAgf7HSJSj6G
ReQRjdAGJNKB8ofY3bRueGQn6zg4DSrVsf8AmFngtc/2Vb9Lj5omRyMxkk6wwmfhpYSNb2P9sYjs
odoXOSHujr1nuO9G8r+hM8KVnVFEj/pAIl3G9X87EBqS1ttDg0D48XlSkwVJq6ZywMBT1buqX+EV
mBB+3Vgdy4ajcfx0kbZd+xZGr89sWrPm99kdjGKgXkdzcet3Mu+YH/fnrInjq3VmmJ/yjxfeZ+3D
QyRU2g+0ZDaEmVEurW2biZRT+DawjXgbId4+1PvAzADocPL2C2wkDdiOpyV9txoVpjJiGdMk60Eb
UyDzXOxQYQCRiVYy4HSqE/8Y+KSsGMAR32/eGFd0uuUm2DPJPMB2/lve7XLXMN5TCQsq061h4fW5
oVpDhQ+b6F6reCXuN/hASoyjUGbkf6KxC6yAiGmCUq5qbQ5XkQfb1CedzKuGjqa73T0YBNAMKm/t
mWmwu5SvMizse0CxkbqKNoDgDdooKyxp1vvHRtAlWBS++syCGvH0RwV9beEZcYP7fho59kFAJdFn
4EO30WlvJCrGF2eELinexVIpRERSxi6wPQo2tP3SArJTOelYrosVPBlxOjvg4SxL1Txzyf7ajUwR
So4vGO+davBvgI15zo7nxenIWYoudVyfYTN/CG8Wh78A4xESM4/coXeQDZnZslP9HDALDV4Fy9WE
BFIFJ9Tx94wh8mNWKac8kTj8L3/UPxYjBs5vZ3/6kq9PMqYV4OJ7Mex/g0QaF+WmQOsRjjMC7zGj
mRgBwaTjs6hY8KDHGcTwdecYIY1s0F7hq2Au2fW+7YPGzU9pAB4h089bD6f5FLggDUnhRuujPYjS
I9Zqxqc4f3goh2yDPfyRsxrVmbnAogVnKZP5OXVrtAa8utvNKd0tylTnbz8O/blgM69fKavusyal
c2FJu1eLPtz6Jev9pGeRP8W16sEX8AUOTdl+5daF2V/RbSbikEKbhDF1Kg3oGkQnwyHTf/xtWuoL
+j1McJs8Zv0jg4//ya3I8BkWcRc3sTEjomTVwWsYx6auDuU1jCG0bHoInFAaIkdv7Vs0Jyqeo1zN
URt9t1AH24Trsu1etODLaPC1BIxRxAVDOVlNtUUjeaJ/DKIHcmXksiQBgAHdlEfKwnEjdKGcn8sa
6321s6ZmGrDG825G+9dwJLcJeGuJxgtZ6siAkH6vTEW/O4941T2Tgniw0YgPR0yYNcv84WJUMu3J
DQ6vJ0LEFwXl3iz6aZFjvbWIiSbSGIAPWCPJQKxlVwbTwbd1mW2LrdqK3SGk8tmFHLo4KRFp0zoe
n3NaqyrZmtcF3tScOwnWrDYUTO4uez7dCYdeLEKyTvb7jS4oQzbjLZgTQ0RKKRgD89hnlaxu5VJH
bo2ARa+TG8d+oBd+YzY4Gc3QyU/EIxMu1la71juh7Fpr+46QNSz8HBQy/Ae8BPKpKD0brjQ4Pv2K
gXT5Pjg4wcdFkdVfk2Gf5EE4SGMViLMEbGsvdrG9PVZ0mFV57V4zqLXfTOHgQiFC5sVP0p+rnMj4
K7lK/LEOnjwCHt7Ri8KwJi79uR4NRoFbZqK1HDonO3dYisrp+jLkd+46Z5KRv7+DHwXu6Nslzi9+
eenrNjcuw9rsvIBNcH9jJ8qs1fNoO8yZhoqti1rC9PlPJrCTHWmS0xdXccS38cfP8ptjmKKpDtpl
QBPT5n+bvgGHOIVmhehluSTPdyiJRLl4kpPOgCX+pn/U7nMtLcJubd9Kex89/r+qJY4Y6Q8jTZVG
GxJUgU5hnaw/lv3mexCCX2txaRueHXBxnlAFgtKIljxx59lSOOFB04CRVz2u5x+LiBOZRwNIucN9
kqBdkjGApYrFB0jZZDlGPCpHr6rWG+EkxrFIj4PojxBGtFTvMHutEDQcwjb/KY9KZXQol0fnfPUm
TyW/CSwQlADsvw/KoyuWNUXegNMYG1qpl/+AG9UdvBrBn6u3uY9U4iOdavPN2xr25tsl6VPlns7v
eg/lPa+JqxxhPLDS1/0CY2Z+DsPKPzp0PMgsWM+nNpWimZCK8feOT6vwH+DGCGl4uMeE2QqE29cL
/iRN5sklHw6PXKp9RMQ5MnOdLSS89o5Qq3vFsdWIhjKjlaV+uDsxLIVSOCAvwcQMkBkBWA47cHyM
ibLYQ677vOr1/CaROEkXS9u5CO4LyZpUtSFUFMITFMx9ehsbFGsZoTnQXQx5BEoK0IC/k5B6I9jt
S0Gj2G3rz5rVSyZo7lwHQIixnpHAipQ2QklzztxKk/A8gVP8G6n48IU3v3EeJ+HLHN+r9dDHOKA8
0JAJnOX7PZ3TXiSloBATUQIUGKbN9u+hCvUBMfgN7Chs4NCoCyQOWHkPG4+zVHgdw/yGjyGUgYJW
LqBaMTVWQVKled8BRkZPpsyNfo8GRuCJGF0DiJNC58Si1Hx7gGut1x+XH5PqeueHTIzNlcq1vbPp
JL5rC/YER/682cbkwEIdccAOQILNaccBx/7WiMAkuO2NR0O8G0nguQ4Lgz3nke60eDtZZCUgS7iv
lgWvHLx7+eMFAmmaQT2xAXX+uZ6oqi0l/XNgyd92fDQ642c73jG4OahL5lEmsoueAMuByg6MObK3
P19IreJ8lt6iydjbEUy6tYY9N2J4eoG9iWq1WLVmb0smMMrfVgPARbkngLBjAYLGZeq8/8CuFqq7
uG3Qfq29+wqRESrncnWP7RF3rBSESpIMrFnPbNEu4I/deRmMo4XTxeosiTQUbAstnkoldSIDO/A+
mDKFGST/XVvXIqChj4eyEmT3PADXV7bXtBp5pop4yKg+6MNXfdG8mBMl+qdSPVQAXxnzG9ZrEwM4
jHq2oVVdER3rhxd8dKbsv2LTEc/ChboHHskin+JKjdG9sFjqajSboQXSipJO5rv3n0e+F0F8ggV6
pfU1QeQovpz9UGcx0Kg9IBG7npMOEgD61InsAZdAFfea5i4UngsrVsQVyjv4y6cEu74oHfGBhqTZ
x74a6PwVdIge5YEphN5B2EwiFYZexcETRSwcsdSB2W51Ld87WBHSe094kW4rIYsB45tH5PxsjWnV
QCvw5tC4MoVWMRaIeIK6rXRYeuh0qQza8RWLTss+VFEQC9BXNT0u66IBoUP9piUMZLk2/B3i9TaF
TVmBJmDxBFQDBZ+G9qU+62FY0iC7ubQpc4qWqqbcd+3QlIwwYPfUDYTDCmO2fD5VaWz+wYsOQqn4
RT890rm/GnYrwfYEKqiletxJsUGlSnxBSusOSEZhsEuYa730/yeFgPp7+cHIvWbLloHKrlSk+zQS
GByZbn8fLKb78RRdc0HKBfzodlCFIIqfLZ0gUuQAHLJyoy8CotXD2HTp6/kAKYkDEyd639LVSWHA
noXN/aegSW+851T/HeXd/PRlY5KT2/hrAnLCAQYWVHq4SP+1ZoOe+MPYyXB9DsReNDTGawlopSJF
+84Re7Sjf86W1SOYWVZ6sQLRY9i9Ryxnkq/VAZkQWH8L8YJ5J3AAx1VMmOUQoerUPwhiOlkgyraO
ByDIpqDb8ZlnRm5DizyfKPfpP5hV6Eq5DM3y2DcZz5B3Y26Z3NfgGnqRQl0Gu+K3jaywCMRNYYKO
vk5osextRpSdOmBJSM6tk4iYH4MA1WdPbo6Va1xdXnHAA/xigokAov4ExPzy3kHHukJe1+I4DE9H
ymnVYxW+YGL8Hvz81uBkjI4mq1mco0tE8IGrORxxJGUSeP665eh/tCoC74t6PoknLhFowiE49DZA
BuTp3W2oMoZVa28vZtLAm+lFhHWtKpJpWM6wjcI+VYU3ilImyRzxROPNEmpELwu9KwLW/J6wbepk
5lxjAQ4YF+QICvV+Nb6Tp2Fdv672DDBZaL2CLx+ez4nKlY9LHv4wHl+4eYo8jQCK2aJuQYK5V1kr
df+vF+pt011iEsTKG0DVOmOPhIWgDG2O31VPPmtQBjB0BjzLLXREaZqHjXk4Q+uHoqDnKtoF3ZCD
XoKw99a9wcZYhOBoPRgaaLG70hlc7ZOnMfNVx1hk0ZwtOovXNIH2xsM5GiWpWvdND904kqph7kqT
JGKrXQJ1bN0fI3th9akuxhr8hk6nl51RLq7upD0M6q/YFp4cSoe2WOvlZQ6Kt0rHRClPgIvKcUYR
X3TMUzAHgFvvLoNCY7rLrWS5VbmR8YjJxbncr+IR2F3U15Xte5H4yaRV9UQizGUStRAU9ayHN3Kh
6IwG3LeSCT+Z6zW22ah9EcaPGgZxIj4FLwhj9XG4k+ScY/D+YI6MNhReIAC8pSG+AuBaIcuz9nmr
SUEjFzuiVXhgHXvlCDco5V2Dv0s3xiaAZYXbxjW9vqhINYy3RFkS+EARE7JP2igCN4OEq1k0v1BS
YN4Mzk/b7IBFlIly7pC3s01wtau8cCm9WVeWTI5htoFdVstiT32EP6DCQmg78lvfL/18NN/3XXJH
UUx9AqTuTAFleJprFXPt3VZCmsl/hTvKZRhCoJfJLSpGMepjv7IH0WXobQb0as/fvWhnUBR0ZRU5
QJkyFUl/lnRw8fL8xsQOGGuF3C5vLkebF1WyKev9kxBy1McNoxjvMe1LJLxczSQLlvlL5DP7r8xn
jbt9KMqyhnfnmtiCOce5BxvtKDDAIxcf5W1EfNx431AUOAgsQOXmowd9hfbJIt51nMejO9hBOrfj
BXU/0yP92XzGBPhaY9w8ukfEgb4OB3EWq2tugH3enZkOgT/D8rKIzZCOBKHgSFhIyM2XLJABoNyU
y8d9HnOzW3VYmRNh+Fwe4vHnZ68dyUnGwA+qGQ8bi5CYVGwFcXu8JUAKFYLN5dNTskSLsE9i0HyN
hnPKxf36gH5b5gNU1lZ8whPYiRzXSw1acX3VZv75OEWcYzDMwBIJmPnmccN5OZhqo8XXdtaWlNd+
wpnz3OfGutVzyajWZtr6JuhggaX5SD9K11RG9cnqsr+wdIYXEG8XG91Uw7coMdjOesnYMGQ0kkvu
9sWqLIp+3nO5TgOU9P6JEMOv1xdtMB8G0VYUyaq69Z/nYcsAFMuFLjY45xoygC2oK4eQ/yc7oIBt
zFB68UOOJB/9f4cVQ4UMjwMdHGRdq9VuEf0lumawk8dZ2qlgHecVw7ic9oAwNRYbY/9gxGIfyB1h
uxfXlQMjrH6OEy0fit6Mr6Nu2dpUt35l7cEEAerBTeoOPiajflb0Qw3Fj4rokyD/Rawzt6jpkaB2
t9EHJIt1TM8Jg+DKhBdu3guaEn2DoemthjvBEk9x3DS6DflUkn0cNYupnDH6uM3XRKYoDxrMEQL/
goCV+eyTYuYP4uIEmn8JIGC+cQfy65kE9Sxb3HGr9sh6nf8LKtDfYbtUL6AzBAaNPg3FtgL+AHTN
PZW/ujfTs0sYKMS1F2tMV95f4siFKSneKQqrwgVeCbTJpAHyDPhhXJtoOrbBJGufxEaPutDXuzEX
1Ap1+ySojjvTZ7qK+5LWElpLTVzPfeubE9dS4R5bDsfOuYJ7/Ke1IvqtcRYUBReuH733m1RO4c6w
gemhEJgi7NAPozcOC20HRVBWrOiPjwvXU2Qj+AHJR4lCpAkyXNWDNMIdEIrlnPT4Br2nSIDM1Kqk
cOsAAvi/652oTbC02+h9GjA0poSH5J0fr2ofC1MCn26nrNU6Y1ON/Y+sXMzBcPIscmmk5iLffDY3
PHs6q3fAW8+GIHmfhgHfjrg4W074apHVXOwFr5mCNBwpNRhXKl5xZMjSHp2PjpRG96wvVy1QRYsm
K7HDeCXvy4a8moRUabD/LrzytBiMslI+1iezanDKl9nmFk+FPNPJCtlqwvWsPNXROY2i7TsmmAaE
yBZFaaSf7BOQEj2kM6WMar0WUOE0HRBPbx9a3y3wT+zZjHeh7nRd/0P21Btn9zi7s8k/kj0RmIf0
aPN0bsRbhw4lI6PFUWOdjIXWOBpbx5lyQ84X9oOYyiyXu38M7x98RY3M/WXJdrqEJ5CfPGp3J+7h
791s14fWqypTF5xhn4Cko27vqKown6HXhV7Kj3JsuyJkKMK0tRAroCeaOiPSN65t0o7uRQD5e7kY
yKHBH3tqLKmv164LHgb4zaMw0Ub+9YWhXm05rqwBOjB1et5SmVX4bHb2hMQsqzlDji+6ibMjwve/
9b/X9FjzfFkBwPd18tI0mpkhnFStkc8D2/oGdYk8/oRIUD6prdCnkm7LW+5TkgnlZn/na65lFqgG
wTkIrgFNhGa1sRwahu7fiOkVKhSlVezpRVFuZvgpMOnGulwY/9rgI0qfdvz6Y9E07FGJdAyCFV90
g+2b49h/OQFdlJRhEbiKlT6Hy2H3elyx0/HA3VgpEIIC3GkSGJLXxR5ZDO5wnESaejiSDGqGOIIo
gS06eDKCVlOprUvz9rpsXX/ZKQ7Ee5ENhopdqqOs9ih+MN6+3wsgZYsw/a2CRZFZVAsU1f/tUJm5
ONHaMcKAiDjBRGUkmBIsC2Soe0L1ZU7j2txrYLz4DRzdgBvXw2aTPDxjfD4mBFS/ZsanrOAjvALr
xWE2z0aP9BSEyv8CKigdmgJ4XbObKmSNddE2dauStdkwnEZhS7ORcr7Fa/bKBUzL9Qp4n2QIe7L2
I+vaC3sA2+MHKjoJWqVuSU2GOKTZNxC9EW++7WcWA11E67/3cG/As9KiMuGX/JBzOPxdoMoOkszB
RWwkWx5zC+HFCa3GeuQwzW7/w710BZ89fOfW75tNtrFGXGGrJSBOR2NiaQVFZ3xqIgnytLmzeXgT
sWInTtbOIQG9rR/OomOP+8Wyw54LlTUV5B4cxUD7s296WxVUazLlf8Hv56K6NfnImS97h9srIWTW
3aITqO5mCzl4tW5PGAKIv2B9dtsaP785y14u8SB8qGMTdJ33livtQNtt5kodBYW6k8EsGVZdkN3q
T0fxOuudTbzCqTKXK7ta9BxrOWDETyrGB0CUG/ITpbKMM7fU5DTFO2n447H/wd1/7UsdMYaYvb9X
URPehoWw8Lv0Aoi/m9Y1zOtI/eqzfCgqvcDMeu79bAV4pEuOXB1rdSIpffYr1Ld1ybruU+VZtJC2
zk1vmhK/kK84VRrK4vEu6JKgHadgx9iUpiIk77X88UHnn3DjfDBcwE3gZRhlE0bt/HPjrjq5vN9o
GV5TYWx2Hom8GlDDVyz3ylXVFKk2JLAx9VQVpHYt1RoIcwE2zP4qyc8Yd8580QrARv2WkeeNqlL0
ouPofTBC219BznwWYIdgU7luUtPu6wxiRfa3km5aEKLS596uHT1CGgvobTe5DekmPN7p+2+DICVt
pbFilkIMuUAVWL8BnEzyMHVXU/Nk8TZxTBbqWUVHNZIDt8uH68mfO21j6kt3x6pzL4mn91fZ3S/x
K1OYBdjuSC10904PDG7WiUv2srMrwxPFcB32ISmiAbo0qalSsSVBggfpcPTeyE0ap9D/vOSNLtgx
H79Wk4XKUSXl3dn/MocHFAYlABQUN7C0nTGN20V7y/wp/dNdLwGykJ6J7jg5j6P3OuyNt4JvSqcH
/63SPs2gOS/CNNYCncY5Q6fUiPf4JuvHDZaIEfF4Aw9PutB2Os/KMApIskaMCjK+jVJQfozKui27
lzNfBOogx0Dqec/wGayBxQ8nHbELUO/AhlcTYjxWWgNXdP5Sk/dnOMrVYmh+IVPBwMoPN/VUgLJ0
PmQ68EA47/R/SlarH0x0ERF1y/7bgj2tNjNdZd5OrjiOiHTlTYJ0dgsJh0StWK72XKGwH4zhkRRz
uaMUrYgi5+1fHA/UNwUWgvgLeZyBX87K5x6ysBnMfhiiNsrjdhE/cEPV4eRZQJPL+PUgHOmQ8H3S
LwJa/4o87dOmcHCPB4quevWEl/yle8qeELOsPWnQfrQ02BXHFD6UMau7yAnCVLpSzUnAwxKMWuxR
rdqHa9KYm3z8v/FaRVS1GaehThJr3gQn+eQ4yvGm8bcuVzJ2A2Z7agcITv1rx/cuz5qD/SFNfwJS
IeM+H0CC4F2roFVidzWo1Qvx9vWYW232y+d0FRmKpOQ5Gm3+Vzy6Eg1uRmfBHCT2pC7S4U9RtPPy
jIXekdGkBEgz9JSOVufyqC5Kuujoq3sugZQ9ZCbtNiIF/pW1yHELgQGxAacDw0LIStTZPLuRFlx1
0kyy/zH9YHzsFrskSM1CNWzfV2mS0y8Aa0/OY/dYPj5lEMJNY62TyY86oz+08M3UUKwh11od/NNx
CGyKyhOcxyLaY+BZiKttdj/4vCfrtl+r2dtibr7QzV0k5uIYQXH6S749vF3iqgsV1Zx9ma6KMKMx
mu6kysHUrm86M4+qC75lOPRA54FEIurqA0SwRTF7hDWx5N9CrrKFvgJcRoudPT/onl0WgrdtP3PZ
ULHHvmf1I+0ZCMjqXD80LzvOjD8g+JhPLrpknMjfnc5PYgOu5zLGvDHnqRLpfiEczkQV5iJNUjQQ
yBTnxaWpYoOvaTKITZk5SvDeVbZIFykrQKTneZulgsqKE4RlLBjdvELbbDoXPiGdzA+0acOPeVL8
HYcuGNRO5gFK81hfTiST3QYDXTRF/VgZ8zUcfiJT2u1UFKdLOaK0KxyRPIiNJ5R24u02eyX+7Z/X
frx9hU8cSPNpeByV5l630SMU8T4lLRaCtN9Q1X+xMYuo5/TnTq5+caTWB1rIHy5QZwnN4t4Ghzu1
AHCijBh47wT9XzXzpvWtoB7KXV31NuQ4fb26eprqrUO6qG8aejbhSq/j1qz1SUYI8HOnXGE3N0Vj
YT1tbNqi8SEtufCvyDxDob6JFFx0zLMHI8esd3pV8/yWeh5kgAFlc4326NdHogKNm2ghN5+nbuHe
7gyvPhDyD86luDAYDrUmkjdqm25cDVXCE3EvEFBXYcCQRSDs5dWO8KQ+tj9gkusp8XPMeJpt5+qG
WR3d8yaXI3URVIzqnuz9v/NHpoibOpd/i6jWO4XQu+EfbPaJV7aF7YitpTqtJMTEmF0P86t1UvSJ
9JJU9SsN2XqXN2lVEA93+gi+ZmZuLpbsa3AxZ/SgXigWVea1ddSNYW93eT1b0yyZb7J8QYnT6Gw6
3odaeO/abdoeRDQ7phmKX4temMGg+F+fmcb8waK4NmlOvATLXwaSRQqe5gug5m/NOp0DzF7mGjBv
Hz03ySW2k1fI6g+FyOrwTkwDcNadPk5ODzkX7GUOKToTP/eVw/Vcp7yZnx2HGGc+6GRgpqOaUGCu
lsvRr7J4YuIqZs4pCWhQsAthB038rRBx/Ya/NQBL7rjFst6kJ9pJ8sNWOByqDLUOXqleMWJoVrXA
DJEzauHlrOAromNt9ZkAuPy9nsuAQvn7w07E+Tqe2lIPirvcXX3BxXdtKx2ocEGifXuVCGB+67Wb
AUZvEvDoxk/sTQh7+sN9fqM2xoK6ZKNpjZDXy3GBxQbfXNhzxmfpm+jO/p7HHPgMTI4VFqeIRQAN
sVTiHHq+u3O+pTGiada1ZgupfkSU1vjZ8o5A2rIBCcTGe4qF5JFf4v2zx8THoraEKenu7rJLUvjw
kCv13EsMTJuF5wetuHw/SJSGQrhW7IjI4ZSdFf+LVnJ8pvkQ0349mPwruu1ibBpgtspOfiDS05x4
nYJ+LcddzXqupp5pPSNb+LJqfnHVQg9JUso34Ux5PlRrwmZdxKp8m//+RxpfyQS7F7uyUJYSrzlC
T+7h0Wfqxx4FC7CS2ebGhsIcrytqztdJgBozkb3W6exAYlWkwJKGFeQpRAS7rqWKESW9kv7OLy0l
m/jLDv025EjpmZyV2i51zgx0x5t14idC3LGd0/rdd0bUFDhcrjK5MJRcvNNXiMEkLL3pvY5kywc3
oGFSvNycfV1+RApIEbV64lfhqwlZP0gqfH7f48GW1xex1gqDwgHg3skaXUONbSQCsxOFi6f7S0DO
jLFhcW7YLD4LHSZUaIF22WzAocI9vMwxVQ91ziJ2XSWaNvF3xYdqzgNGsO0FIayeSsWpewsfScoa
mkijl60DivxfYeeWGu7yszn39qqxxjR08xlvePbSJz29TAojp9t8bsjEm26hV/H5hpQLiNsQ6lBM
M74JgqGMYoeqLOcEd/x24Han5ta0oGR+GdM2rfJe2ocQFNlq42ePqs4w02R4oha8IKCuFZQ0Xjrt
YpKxTMhhN5Bf/BoB1H37CQbHBqWG6+LPSCNQ+xWXudCpvh1EwJA4bi1Ugyrk6fwkyqOYWgvhzpzb
pZPQ8lHwJCNd/EpeU00VDVdZ/IC+YWhg9DB9w8MhGtZEBnW105WtKp4Zyg62OlqkNnMvCWqomuhv
J0NUR/4XjAiWoJTUoU3L62htnzj8GbPJN3xHqyL9hw4QCEw6+KHNhv0O2JsQzX0Xa8mu4XkqBV+p
vvkaL2HN+AyUwG2rczyq1t6+4yMsc6Ai1nLEdrZGagUVj3lxkNm2pmwF3VNA+A6erZSsCbbrEolW
1NRtabNbOCBZO8IU8ydN8uXHliFU8Aun0p6xg39v8QLOV38dTqlwlW46DAI/aZTAivVFs7trkvYL
DzuJJe8Cdy8DYgaKdjAY+ttZMNZrPK1eo/Y4Rm3fqzC8ltrqWVVNEWPlukkSEr9PWlVoipnzUI+S
z4vhOpH4ohaWhdGAe6vbHdDjM5iJtv0IBFYuI6PdI3vM3YhgheJkZPkyCp3D59lW3h0Gfa9y3IXy
P9/xIgAE55iKE3Xw22OBEW7+eO0OiaIsqUP3ApxxZz8k2x/iehWFfMcsNixFllzGGeohEDOcKHgp
aQDIykCT5AMfHSfiIRBJxRS7Kb4t+lsWj4vYZ0VMd9ucBtWvo77B/n7mxbmcLe+68JuOkh/F1+CW
6vdZjHNg4nuxBECpdEd9lRbrbzkHj8x54C1x0Fv/wx4PDFOGvjQqKK9zrT7cEg2VzKgIa5dU7b0c
pU+Vr2kFHNY0oZ5vyGuAjXmzDBkucpi17aYthvzOuy8JSQido+OAr+1n4GZycMGwX8ILUDBlySSc
wutTcTmkLXRaHB7NMDvSFWhYuinRIQHQuGR/DIxogzSQp3hL/8Ez49Jui+W+gcje700Kz9kW8+b/
2QZrhO5ctrc7rDpsSO5P4qY6pby4tmQNaLNaOtjgRiq4mCyFphimvP+RUuahD9Gjllw5RQj8pkVH
1iw/A0HCzlvwxoCan3efdPT7X4IORzucKOw3zRq6g7fF1b2Z8yMfpDqLfBXEDMUrtDhvm2C8ecs1
pfnedtY9rCpSew/4GdfcsZ2vm5j8J2YnAuQOTn89nh7U5vWQQaqfHCJjVCk2/0SdEO01PsRoI/05
ntOlDwH2YtbkQ9hEsMAmz5AMCzYQrRkfrNH6Y6ilArGZ4sNqwPTllMYTpMUOhSqIQ9XpSfH55cpv
51oQREGwgfJZGfOumtVmRH4i6AtIyZS9xcPQ5oj4Ss16+l8Lh9jdRsQyDNNtptVUx/YDTRSvhwvz
BwYMk1hCsEmpUBJ4I5nabTEZ5cUCXQyJjsAC9MnAZzxGxiXaA+MFmVFnLwjT6wG8qrQVxcEQsNsb
fSS8YVjl1lAKru2s+Y6MVe6TqeRA5f3qlPGvy/dXqnDBLJMDrCgnqTFnU9kkRyj1zj5VuQsHFWYY
iOlFwWhxrR53k5OSpMaAcfsh+7RXWT4Jigp2XIuen/bE3Z0WksfjAptI6z0+WqsrMwTaqtYs3VMO
Voz+0JS464Ma0OBcJ2XLC+U5n8tfqFLkX0+wSmqpXaPEaZk9d6xqUj9TNBBfUryYHWS/rB7IpCr4
owGGgxt9DVL/3A66yZ06pqYfDxdwlgty4c/BZ3307qUjyBVcMJ2KX2nYtN/vmDwlRpQX91iE5+W2
KcRLuwJrWHhgNG9jsLOgRv+fUYNTswuv6K8boi02K61lw3BJeWRSI2Yahrsm/MFPZjfm8MJ768YX
GQdszkpTlhce3WrjZGi3J2s1wATGXStvdq9sYjm2gLCPpeFn/5TLPjomjLhoRDcnKlDR+S5PRV9K
HlxaqYu2cNwJInFn9B2L/T6rpW4amp0NaktkxiUEHznznucB3JJqksy+XvdOtRxVelA0rtJFr9Eu
/ScQfpIMrakqKzrD7TLkO1+Jh+1M2Br2sQMKttDsItQKiz+kyQKFsGRzNjS8tqCyjFMdR8CRyNgS
rbVbheQ3enXne/NTGa+sBms5nTf8AeFqwgBr+TSBEbwrgQQ+JmqOXxfLdzkKNxt9YVZXu4iehhm4
AjqCl4S7bOK6SpmgaGzuStkaxlvzVslvXcsLqZqmOSaw4uhfRihpiYf1Fdr838C7tR5CFLYpEPaj
qSbvgoDtJMDtKIMLGA/cqZ6UhMRC8j7xkQVYLE1Rt3GwBOlW7l8DzSLlzOa99EmJDEnVVzYokiIc
rHGAphKwTDWiEWmiYIvtchYjH1ffywBuMa+hnOYAwYKpeikxQkfth1ik0ZfxATnrcXuYjiDXxHZy
VI9MP6KbjbSl0gMcJlG3HvmG9OoKPLfD5UMqjMJV/rbxLT1DB8i5MweGhKoqlHyVmPof9xncGX9m
+nMnYhIiSVr2rsaRBzv0X6pYxPwk6kwGWBwDPTZpauPBkCDAppJMDGcsN752JvezbNLhqPKijlO1
ikiYGL9u87g54RZuiCgdTDby50QWQPgn/Fo3adNFMGopyRSlzPFCL/wJkgCSPgposGXh8CNc9uIc
c/ZdcihLNEcd4OfxyqKXLXPoSWIUfUWyBKpuD2lix174OnXizBLEBllfO6g9vnzDeGmdOJY6wjgx
yN5zgmQs+KPWdAcgw7KmvstzioB4ajDkzHEjyPjzAAhJ1hZ33q0an/05CyshTtSsu0mMnZW1KflP
1h1WOWXgd5bsp7xVgDrpyR4X8BCoU8mr8bboPGJbpoJS4CfY1BeQ19gItMJKxh/1vrqsgXuvS/bI
bllSKBKrbp0+TOTSv6yXVzBVvrHOqig4U9Q9IDwauHtHCnbXgzKVF1syfuSS/ZPuUqnZQ+c3X8pp
SCDfnahRsEh1jZl0fsUyJki57UMfz9SaRMJyZiSdaT+cwUtPMFkwpRpRDsQS7pEs9Mj6mZ0dvOrc
RZ9Su9P/k98+Ck8hHTHjWUZQf40KU2pbMKdflGSksnOKMmUR4nApd5rFSKLq2ZI0ugRtOY7JiBIl
ZPVSbUzE8UA4O973qbkGrnqe1OTglfxafNFeOZsCiwiTpfQjT5xIOkDqkWK3fprrhm8M7nDPUDRP
O2iU5O8uFUYy7+dik0dKwZL7zW2FhMdn5N/gfkd9ZaypdVCwFrBK9mzRhYnBNEfvoE2EPNbJq/oz
XdunoxfF5TNGMLHmmeT7BWtRjGSUXOCuinPwY8wAB6nrWn6djFrR5A4kcnCsVJm3/t4a0pC/YvF6
5dkQ4b3d0UvPRhSXQwv2/x+gimeSMcPPmVElwukSYS706KJjPK+QmuCDVoX4a0UE8IFzHeMJ0OAe
3ZQTjLDZfg5MOKG4gxyYbW2PZCAn37qrl50qptXJXCLOuazG69Z1X99VCIFyl6RXhnbEIQ8VSaCz
eJwBNbqP09kNDO2A5un+p093p3kSgDWVt5EsFbGG0qlgvvUZ0R2mDkSxHqglGSUZ8vJD8NPe/P0O
FA9WnC1ElIbpgXLbcfgJaTLj/n1ffQeOtsTEwXmdTiECaEXBfnXeiinuaaYWts+Q434+676MlokV
Nd4q9hSZ5EMG/I9MFw4Sojn6j5LxGxRl9fPYY+nHRT9DTBflVDq3mOdLZG4b/hX6uVuaN04WWrmK
WBrZPyXEM/7FHVyJIDbGCqetebz74AAVi5FBJRavSZfJxhc1EkjzEN8fFA2l40MRE95UVPzHowmh
PleNE8n9fG4MvW2d4SJgquy5XPivCcJjrXBWBrcGVpJP7wKROck4ZTSkyQ4Opi5gc0N/yhFu7dCg
uMSHII6ldAGkCOOi3LHu3T4MtddIfa0hekptYn8bsZ81elfYhb9nnBrWTo6iAFWoyJPz/O9SChbL
SV1Ap3obCz6b98QCBou9fezkDHDs7+SHvkPXw0YNMl8oJb+w3xdVXtkJamsMiqcVJml8a6BIqMeu
tBk87qGxNAQsDraBuhQRbNAJOHli+iU7ZeInAQdgv8Fa8Z6Dd+OqcntZhhrKZ5KOxPr9nPKDB093
6O5vP6J6daDik3HqDjMs2aHTr7uatr0WOOji6lq5zVmDHHU3cO7eI/UP/bbBLMbfi6aQznMO+vE+
GkU8UVfEaSfAb789uTIhL4bpDDbSsFFbkK9VNIfZXWsbnuBtq2d//Q0hakKDGuJqevzPe2WOAzez
QDdV4A8p7RJYWHgG30ZjsMFGJ6jVv/w0LqoCLGqKd+e1ol77Rmq+7lQDIWInW+Phcw5XsmzwvpPQ
GxaBEhVoALImQTPLcrEtDe8vYscorfLIEuO1UInZ6dklfVzC5KnlcdO2If3SY0WTzhLwPdwvmkia
nuOQ+utr+aa2IjnuSzP5OP8zTcjoAoxdqz1c46GSKIoGzrmakedpdJoFP0gp7Bx0XkO4KLRbQWAY
L7qb3w1mcmDeBzxRfhG+0XBcty8TIdrwuaCaNhGICTEqCPkV732dfKz2ZmgEwAMAwKP1M3ZygprQ
HOlLsNaYp/x2LdzDpHvqrspxT6RtS8nByTwLt7Mgr+Lr1Vsl0oZu4ubJmGL+8rSUN3tFeYJ//Zt3
0McuRcZ2zJ00DG8bl9qwzgEc6adie0JUsUlM2PAUGNRfpVeYuEERo0G33TRy13mUH5d3mkWuPaNA
vuVRm8cKie4kqO/lATdOIBBSaxlixMdEDg9zqyOxqK8SHbij9ulloK8ryfGWR0+AJ5GKeIuKLvmj
gK2AQ1Uc3FG1vXYEiUTTd9p+6R49tpogq+f+S95/PJG0lzZcqCDwBXNTvg8rZldnCug2m2nYvp4b
tgDqJy8EZ8i3oLVVmuamF/o+8fhehi76Rtdsj7oA8S0uiSQ5Cf+/R0ONrEksAHyn/aWxOSmGrL+3
dswg3+TxA35Bmil6ylgKXjF5l88LdCmBLA9tl32pQxSQT18KTj36oKp8eO3WFtkBVawOO+OtAKlg
cehQhAByF4fniAcJHAdG9JqVtiHzR1xsmLDlK20SOxz7nA5mjHWlEXWRwDpa3Hpw27HljML2bhVr
furllPHzHdd3d1kn38HaZn/TPZqfBaM04jqXRsxVdJRIk6cv6qMoBUb3exhrX5pg/kF0mCh1QXST
asXLYqYHYYS+K/bYf+SQ1ubnmXA+6dqAvHexgZ9ATDL1R8V+cHR9NwNgva1VWW0N2AiaAVQ4PfyQ
mlhBKXqIoExk1yWSUVjXPL0FAqHaEyWu/86RSswt+XGXaRqTsYTYEkqFc3PE36/aNBN8cR7d5Jm+
Q3zQ0Tkylong7Epf3JUoVMy17NzKIdqeTCQaP8Y79pcAh/TEWNpYIP7CPGZ3OqSUmJAlUdyJnHOz
V/0M6uV0ZdTkMfzWU7DGN23jk8r6i5PnKAKi72XtChauZFoeotbUSdudDPJAwbc3c+9wmghXTyo7
AYtwjA5e7MUkmH3Lwvs+FxOvNDzZoiDXQN28NSSQ4Jlsj2sCsboMtWh1OS312+XISPf6s+PSozqt
jmUAzMUo2gZWCbp6Hrw/gqVHZX29oCvrs2dDRWTlomUAAzrz7OPAW+9ZTm7nIHmH9O+mPXZbqm47
S1+F+/UbprxMJ2VqAeF78xoKOx4Fw/h8JsCDgpwOqiXMMYrRmsK5vBhymnbwlq3Rza/xsSHBfAtp
Vhvimqg88rSbaeH+M7jAj2ETkTVosBBkD65NsMk/UCjWKaOfX30DnaGN6j5HCh/fpssjyvLTWJkA
D38kpgY/6nQhKLpzwQRvAzvDiWKZIjtDSuhagBR3pxPVgeV8reNVt21YqsUgYLGJyvlnnKvf9Nrz
OieFe85lyOUeLhxCe6tpZs6iNUuNb2JpQu4qmejb7DEASxAXbc+yBkdirsoP+a5CylJhoLhfZjin
Ds5caP/UoeS34h5wg55fkvG8mtXN240mWQfSFQoxj/b6KCIVrKChmFb+mBBzo05K1OBa7t/R2KVT
AJJ7Nhy1SaGYvDPM2ion4e8eIT+qyfGqS0AS0Yzq54crdbjNxvQBxb4LOkNXuBs7XudUS4OiuhNn
vR9b8HLMPiU4K363Dt4OCO4zmsdc4w7MEB8EoiCOzJRWrw7b+P/n1T1Bo1+aSRzPop/ue0Q/T9pF
rHGZXM9RYKHp96JAlgYEeN2+szwDkd9wV2sG+FIOTZGGT25bHUoApXkcWf9OBCyBgLTJNjLopUx7
YsiIKjlI8IxB6i9ymClPIAs0S4v1tsbs5jsWRD+BDJmgQDubr+DabvQaiJuHQv/TDs4RHF44DmJC
IzrKXaofGrmmJWp/FJmmxt0Uvrp6ZqAa1GJ2rJN9Utl7IfllaKP/W/P+qzs53he7mR3kHCJ6pGYm
oMIhovqinqHH/6AifGLluwXzSWsaAlwi60AKS3IE4CIhfqt5o71CxuIZcofo5c1CUaDHGB4cqVOU
SiE8vRH0+WvLXf8NXqV4ODRlGoNBF3OIPjAbiF/mJOdGZnCBkA13e2J+sMbQoiNpDv7zhzGng+yQ
H3LniJhsNWFMJE/3y1xitAVsujKs605iF6adJJ3c6jhWRWnYczyrTIJomM9kChIMXVzcFRZWkXa3
VBxFdoAjuJbsJw6P2NZBVHxj5zf3N+5aCyId4em0Gh1KQ+DAxeNyCsplECmet5bWhPQQv2mOoLDq
l1Grcb7z7Reu6cuvopvG5aRXUgF/yuq5YKWBwsFbrcqBeta/7M+gl5P82/zAquhV7vt2OiVvoVtb
cLiPTlTHaJeazbJPW/5NfoSu7TDIMSKcGppI+XoCgiZdiMyRz1b2fxv+N52dFrrpnaYR9LgWQ8F+
9e3/bPIM2dHvDBaljEmube9TrGvLc8qv1Tfgqdm3VVXqx9MZITAsc+P6xQxj4gnfF/MiXxRFkF2Q
VieKmR6zS0zIsohkIg1IYqTGNSc5xTvRy2Il9uVC9GRLcGupFN4smGrxC03hrbMisY3udESd++hq
NDk9v6ErK8B+/JRmksc7L8Avco4eqiC4iODk6NPg6j7gfhX1xNmnXsMouMcaunv8EhDAzNvDURIy
Ayzx1hvqqmjPbU9IbT8v4THeKqeXs9QXtM0kypsjWLt1nWc4jNeBaiBuEoTwJJHIrKXfyFdz8s1O
qOHrY7vi9T7anNanGzPcyWrOnpP9JxyWmuFcpcNfC9Rys0Kjxbde7r0/akk1ODb9nbJsczjj0fIX
w5UopPaQae+U+uq3poGIXewo8g7TZQO7qqiS3ba5dH19hLke+SnMlYSPSe4dhFyocijUeQNxJXsL
ZwmGlRfHSCmftNL6SWubGvapG9OXR2AJdQUhpES9PhLA+KDcXU1IRlObrMttYVXxarPApnpWJPGw
H49i8TSLUmupIF4QBjJGxusTXJbNC28oWNLJ81zREMoqX2zWkC6IPbG22lthWogU2gsKit5b3syi
oz5hAZwyoSneurUFvMY/i16DZYPRWKXjvPFfxonXvgC7aRuSQxQoakco8T97CJ9fKGB9Nx0TXtFN
Z1tmrsfnlhI9j42MKLzyRrn0swIKNhaMgJ6FL31wBZaR/X1koqxKF7almfoOJ3zn229BfYmPCZ/0
/l8XQyVgzlzoV+t0tdQpQE9gGCgFnw3tTeIYD+pnFisRSGdbebZg/7QvUJRLYng9ysX+ttdS4oLx
T5rpyiPLEppjMFbZReHnePiLUbAUDDDkM3vwuoYoHq6P2CI8ow1hEpb+0sXB2EHh20HxedzWZOY/
48WF/SgL+62JUAzJ0Nl0Jyi1ZqWvKei2ofzcLzZqISplwwNjAfQrhUXn2XdCHFbvYjOx8865PQ0W
D8H2d/DIVBMBVnW0OC5+6SBJK4Dfi1CfvduBjMZvxtxTvurEMA+FfArNA+vsxEf5PdBYtjShrK7Z
t8SYjEXKJgERZHQ7kDIVzvhaFmCDl7+y1roa4NFxMFruVBdGhp/auyrrgUxvaaU6pMHenS/t/0v5
b64nBYbwQocAq+GOOD7ZsYx7T6abMgW0JvciU2vdNRpEJYCKGMNTYnT872pD9tWY5ywQy6kY9Cse
t+OhZZLFwWM+6SXloarBcO/2zzlhw8xRzjuazR4hsNaunJ3bC8Pl92XgMsNPv2Cq4kx/q6pFN17C
wGB7Z5Kmc1R6CKriOOsriuyhPGNUs0IhV5Zcf1l6DioK8aWaMKBF6Rq8TOWt8gqN0VPU4FmfjcPZ
aQTH2jk/Xl/A6v0PSjCvhXuJ3nT+jEmMqRcDwmp63VwmW+yjh4EnXThl+ZdcvkTomNcJpq3SQG1z
QQD019KurS1LO7+M867hkXrsnp3ZtucpH66t9PQ95vNI9Qbqx074u8EcIj560TBDUfUQEJZbyNhc
bRm60J+4+XwagUpNA0pYaN1Zy4Ouvo9DkXuhRhWda+awGeKS+QZY7yhVkZVYO3V650WVk35uF1Gi
Yy3+AI+CXxhJL8dU85dttH5iZWSmPItBSfJtuiP2EDZJoGQzOJAC7QJbwR/ARIu3h+UYmQZLPDxa
I8BNMQlE/Co+VWCYXW3NpSheg8nSxhmVjc+xuTK2wbzrEeUVkH3vC95Hp+bKekvOHxzyumJ2RMHc
2jfR+1ZLltkUJRtPoqcgg74PD16AdggsyeHrj8kRFJkDvJ1d04UA4x6A/Ks4MTaW1/JUI9Pd4ujS
n6hx5exvti3yv40NOTlOOSlt9KKdEyhreN20t1A+x251/uXV6Qd8j4Fp63PBXhT1Ye985RC8wnMl
LVFjVXqpKRGU7XA7cbhtpO4vxNdE6ml28at60Y3xce0NmwSH2mH41UdXSHWAu6LleohoCUFAubGp
Co6+aW7ha90aTqLoANTnAFMm6rw16nYTg7d1hNk3kWXLEglp0NHIGAnUezUf1WcDpB+1cAOtPyH7
Nu3afBaXhT+RThQFnYw/F2cnbq3E8Rm5S8lq7YPlIxZZkl1iwvdJ5cc0gU86MqBL30tmeXBKfvp1
+wgZLQTl/go+wF+Lcws2iKMysoiSENva0Wl9aL0+cZ1jPQooIdCYbzGkZ2hdZ6iNxiSYVJYZWpP9
1MQzDx2jz46ID2cvpqCScQogujxw5ixXH8Ro1e+giS4sgTg/5nXrlQ8PmX6J5JAdSLFWDBjNqZka
nSTMeDCwMbokEVkB46pZjmAvGHQrP7iVrjmkjMeVsrSrv781SRSl58xg5/PifDhhn9zgdA7WjURT
mc7TPoS4mizpBMFpIUb5zO4tjQn2YIZAe9V2RA05FX/+T+7hsNsJqObRlTto7tQ28ur6F62d5uyU
w7C5Fa21e2wpnGFYyXVZyur6aeMELCa4GixRtCAm48jjp3PgkgVwzPbVJWI8ift1REvsG0JlRaZ7
uw+p0UTzhYOVFeIG0k6DEztxvEhB17TvOFOPLsg48LhwqOa7w8CGzOmAT5M6MGO//lytVMVFriUj
uyNRm+AU4SDoKABXLoaudW8bYI7yUQIt4y74rtf/kylv+emtmLYsum9rF0rsMA4xf//1W4inoPej
l2p6DllJjG6ibfzvK9fXEVSnVByFErLPPrT6NIzq7FebS8LNOltEF6hHcxKCVJUk4FNIEkE2yH3M
JiVx2oauyvCNEEotyXKGR+bPDO+Rp22R7m/UwFTacfKRGkXJOSGaphe7p0rrXjTb9ATWrkozPIqv
K3N9jh/Abzb4A5doJFo+/WBBNuozodSa1BRhRCL8Kft8EWEwgK4mlO3eq9TMHxW3KBH2YWZaPGJb
sExA/9d7K3gVA70BL9n9k77wWrpfknNIzhejyuMs7/QKYQu5sQ/DlkVmnJtl4p8IIv2rQjtUJgtF
2YmJ1G3vSZDftLuwE4gfXfa67yEwxPmb1V7q7VccAivB0wz36HWdDl8ykVPWHQLU81kIigbiGent
GZxgvdXgeKfGh5tElc9KP88p7ehLeldvwz0+/I76+UiECyg5IrmsvzNxTr0sNxSwzVQBHU2WS2tT
cG2bgmlTfF+P9mFUW14eKamdTYQwMeuWV4lA7JTCAz8E3iXMA7wxsIxD+a38j2vPNswpIRqj07SQ
iefXjVtuozd9GcRHsI6+IoEY4sKjWd2bd8ClMhvQWnEmLbKROpNo8Y41J/27MhOfFd02mWkWzbc8
ChudTRZfocc7KrVER0FaZWfUwLXuhLlZt+6Klowd4wvQskkds0k3w9KT2zbR8j1XwqM/7jY7r4ti
R7BBFbOJO6rO0Or6erp/QzH1SWbwSp7jdV5mwP0tJBZ4aivmzxPEdOPOOVZozW5gA1bJpk9E0N9A
xzuQo1GsJDBZPLZ4KGGTHMxsKO7lJZGbVcAiNKVv39noxhJhyHebFb9qOldMCF8N9VoDAsa+VnwG
dOJbd/MMlU4DdXYRcOx3zWdlRZGebh0V+LXjSrQLeLJIBPmYy1E7XD+YQFqwwiMka/R4OBW63IiP
1Qc/Abiqfx87XNtb6mefouzg5BXwoZNKUJJOAt57WryDULtVNGozRmaPWbpaq5jWVGLBuoTBrRLU
juMITWESmqJmFhuXzYNwkYnJGDRCkvrkBXACmrIOVFLwq3eyKigCsnUahgPReM5UduXwpsIV0gIe
qkYNzWrT9W2lcgzZCjgPYbEmQX3UGNXwxW5QWV9T/c6s8vEyJe9aWr4ARHE9n1stcSPIz2CyvEsp
J5LFgxm38Y5+7b76ZSpT6IamMyn0jPA6CIQZQ8dh0Hnpv4PdAV6ac7bZNQbyItlQrAG5VgfzcP1u
w7VfrejT6f9vImeMe3jUs4+f3nxxAWoOG7COsgbDvIFXcTlOPvnIxDc+S48s7dzLTOd4tQp24YCU
cVUVS0jf+uaS8QAFJf0EFSHiP+iXYt7JdxF1Lfsgqu76byamIO7Jk6c+WbzrD/1DO9C9Mul0WZHB
7+Gei6WwQ6YhGD5sx37cdjMOIhChqbSkxfwtep692/qwJKX7K3b60NtVoRunNrzSetNPk83iR+9m
cCA60s+QlWMsflFb4M7HaCm0r01qDszldwa9sfspnvMndPji+XftM4dwS4b4TtoHikOysQli4FRx
J6oXgd7UoIAMHqwGF+yh42jQdFg2sGEw75ytF+Sv2DGy3iM1QUfDjbT6HL4FA9ui0m+b0+ICT+Rn
k9aNCERS6fieajaGLH8+cXnQZUmqbCxAD/MqGg4dmiaNQJOu+wqUCJtugYqargAjo5Bmmyr1msew
YG85wUFfX5qp6BuQXz3baY3t3WknOGTSu9ErTQX9ezb5+jH+fjgimi3QioTM6pTN6BIgwiZYMWX2
y71JGZIvYwHKkuj5dITAVS6jBux6qT3v7wNszD8IFTsyRKVmSSgWMiwxbN55qvYCQyecIqA1vlO2
giOo42p+CUZfkUrR/QjUi8JPqvpmz9VhlmupOJX6E4u5H2Eqo2nWz41POWgBp8/02zK06P2zAVr1
2QtE1fykI8Y1VyYtf934CEPJSf9NiKtUmcT0blU0/7OY9xt/VgtXZWepIomR3bzzuSmLD/vryELW
i4NEWB6sY6IPLoZYguISLjtzAWMyB2d/J/IehCYTVP8Nhvi+ucQ2LSNnO36wvg6PvP9z8raD3gTw
U5L2Zrn1DJw8KsNszWpijsks2KtMlB4n5JetkCYDi+DOZ92JDXw2Kxxa3F2nqGdtVllxOgvC7a1C
uy+JhbhvMGhTKRcVXsAOHpIVcWtaXpxneNsm4rFG0DOmf3UfrPffW9CtN4bhVWAqz4vu8J5lMtXM
I6TNx9Mi88vJ7eQy4c1czYcmK8+o8AV5KIuYYvr7fNvUgd97sGWG7fkw54zQn8ij+E2qzmSwC1MU
PKw/Rn/XG5zFEgbt1aouHDTkb6bm7Eve4v9aZpdf06RBsWWmmX6FX1gw+MxxI//gCYD+8coMGkhE
tI79RAlzx8a0uDQOjF4iEhtPciW4DG+1S/elfZflI09O6e4lTrcQ38uMATpyiM22js9UiDf7GEOC
9nTnhu+OBhXGvEioMpLCTXUGgmB0xB0p48D8cMOqXZfy3zHS0GnZWDD1XDQYvm0kXYXDJbBD7kbA
p/N7ATatspt6VuG+rUMJS5RU7lNhpmcce1X7X83EBQWNZp1UwidfObxPUd68lCOwYhn6m1JN1Bml
CndXYGUtLYSmLGKPXehXSNOaRMUwFK51JudzPU8F6nQrH/9zA/5bYhYsnzw+yfdkHx7rX5uvislx
eU/B8mFoloNxoLEuqzfEBm75FL+LsAhgS1oJ1mtDdWXtllSooaI0Oj74EyxXhZruLKgqzF3mHGw/
aBCglvCGoDp2fBOt+uiBLRoqo6BivewSz7tYzRh+kWA2178ARnq9TzrZXeUtfYnuBa52dqmMliWG
Gf2SjCMepqcue1pyXuizwssgpT/wyxlfq9Uty7LaA4VCeG0Wzk6/jpOUiQAbz25yZ59/+PNFkC7d
ixnbi1spAIGqDT/jnKoJmmNdqBOy2l6OUMcKPOjk/vLNKpSkUS9bvpH32HDKTBaJhpd8BZfAaOim
LBU/lulUBKvk1kQEP34SUANmQ8LhnIVmfmCHZ/RYjXCJJ0jTLZZbAtBmWc+zvshMKqhfv8XnBIl6
NddztDa5+S4DjIQUbkZT5J1lV670MzdJZoBVuTTzVESIqY5xBD4cpBRXzF20pyoM4ly5Bkav8tIK
3ONGCXJJKFUtT/ln+i5UrO07ofjd+9UI1elsSdnzMsVG6kH6dINNo3q8djaoMg50DgKU9WGCd6GO
pmGkW96e2ToFv+iWpK2Kt/F5buf9AOysdHKMEuMS8rMK7Wz9PSP7JBgUHxW9JVvgYDzp4PQ0A1Vx
hWvvgjgULY9eidblYx4+DicFlUAhZm/3ztVg2bOtdINAQwnUeB65l7HVoI8em8KELOB2HrWTk6qG
LfCegMt485hm967yNIaZW+pmyc16dOGkepb/V+gkH65dO3FbT+9HF6a+LQOSpwYm3Lnn4Ae4tH24
PK0cTQgXQwRalNyFeGSqgz85vHOzNjbpPcIBokqvodPdNajgZOIuQJRFQ0eZrK9kgRvKPm76TKs6
WrBXNm38/nGKqrFMud7uRCHBXvW3RxajK4AJobYjMS9f72Y6v4ZKmjJkthoeKtSzPvkfgIWKpscc
/sn4XNkuKOTBwAF0EZIaW8Om7tlLV//OIshzMYwviqX4rqeWToMM1Psbt9L2KkSwr6gra56zuxlK
CyRVP4OpRtH2xTTT6Re6rtEiTGLwHQReKrYn2mD/C9rBlUW6RvoQ8xtdUkiVOTW4c8+QZCVuX3gA
/J0HwMEd3BXWVWqwy1avCTRF0zpVf71/AOiez007d2qFh2PRYhlaGp/WbMxmIsuSU24dIwDgPmbi
k6HN6H9d+MaZo8GBbSTvB2dOH3Mf3WpsExSfH0mjyCVpjvOE8CDfJAx7ZtDZJC32BmbzlPd57hr6
DpWFa8MuzhhHrXdaSKPO+AHKUId/UxugJtpxWSnrxPsVhQW+NuUX24pu3oLH54Kii3Xdh6Oz3E3Z
GH2JlwyIDlYKNw9Pt/AFrqRBrL4f2mpr5uIMMW3sbiuRp2WAALQwj3IVh/fnpgXbYsuiBK4qEs2/
ag2KqDSZa0lgWPsquE67zU5X4fqjXyxvRzkFcujg8qIME2KameAv+6Hmx7AyRW2pWEkSN7glFREA
qAt6xgYUn3B5N3bJdxNf7wF4yEDcL34KL2r3N6R5uMo5i+0gABUHS1SHUlCttdebNEklTZKyq8sb
KSpkgpp4MTh9TzP0cyGm5Do4m/pNYEY5CIw+wLYVG+LzMvSjc3sGXbd6cIF5j63YX3D4gw9IHF0w
MIdNJE6xRO4n30F1xgr/49KyHKEB4XJPx6jovQe0T9zOYj2xNCbSbscyy3cggw1IUMZXzQL+JG/m
cqrZytMSPdPAzyrjxnlP/Ow2xbZZB+nYz5YbbDgM/04npMzTuTb0Pi85JpRl5z20uMIivSJvY6f5
ZuFy/0tZkC5rZjzn83X+sFRCrds0n0pib3IAyh79dyWYaY9ywGh37LL8Wn//v2d0kUFqa596Ciuh
StzSPXwhAmjBSDNeTHog7k7bma3OKXlPCK6Q3YeCoEWmeN4fAWr0tzHt7PuJS4cYdJ8PjhlwwbU0
eRkDkc4fb3DKOenXodBfRtKCsaWfyc/9XlX0TOhwE7XgzUztxkrBZ5eagwWL+2vh4z2bR6On9Zb0
Itko68kGrb6s3y9Dhdq/8MLegNPmQpGgpGiivHMDjKjJ55yOMPCoh7N+CDkiKjWEcsiCdWQLFCCx
fTxawZfR9KxznA+Y5KvAdKtTpfL2adyzZ0EIOk0Q3hd9B15OPEiO2ps1/4fRjGCMmM1oRGwukBHv
M0W+jRYalAbcE292e95HJGemhmLVt+kvlNt8r7XtJ9sbJGLIZyL34pvsRelC3wx659w1/GrcEU0o
n6bYvvZOAPuhOByXbKSE7+3VC5mcQDxxPWvbGj0zsRWXq8eDEumOKmvAMUCUe3oOK4Ws/IYQQTuF
tycf88iNAJcL1PZre3WtE5zZfwkqTBx6bdp+L2AScEkO2d//HjKbNRWnH4UC1HAhutUWfejlsoA3
Ew8JqGrOifYyOfhy0nKzc0ZJ6oUGWaK2oCIVQZYouk4GjRF3pZyajWs9p8JrNPZz/hka1qSmAQqH
r2QYElDkzEaFU2XPxOpkdIdih9zW81h84rMDDVmMTlhjO5bbSwO6jdUaswetvD9qMcyx+LH30p11
FFJUwqGBv2F5cvmvvvCnmpm8YwPrKs61hhqcSInzaQHQRiUm4mE5sRxdcsg+6gCPWGbfpNHcLR8F
5BxhoaQLNxYA2miuYMxjxL1/+pnd03YqVTVC1bVriXKHNbOBNDq3tVWsOmaItdsEE8ZXXt/Xa0rv
kTTAraWdv6xdrDsvzAm30xPvOaETFgfT+rd2XRLT8G4FBrTPKXjFeCbryR5SGT7M6rnDVHa5kQLo
EFcuMXKIT7TzzVp1XDV2Ey0eRe3f3vHMitS4/v6WrLLZoUAiVaRLWTp9UQaT8Hy0EKTYn3gM0IBx
ianFh/O2ysKRpjlIGDl1EFw3hN6vmJ3N+LRXF5toNTtvET2i7cFDpC8soQXRANBcNmx93ISdZLOR
1wkRVfJfiKSEhEfyNf5aY7t2pSSLqi6ZLwaMQsj+xW26Vs5y5EPEydpL1nnzODvPv7DLDis7kBjU
d3Fi8T+BA8IUNkto7Br1Qx6OJvs/JmGoBK6SIxQKkaMDju3SX64Wt3DlXX9sFo7FSCObTSJE2iUR
K53rtPEzVOdTvE0HLqD3h5hIRSWirTw9AZasNhpjdsh4n9bh0QtIno+Q6Y1aU1xiv/gDaktH39/G
S6WHkkWQ342SKykR2vBvm9zia7z/Dfuxefvt7AeQ6ZIFvv/XSHwpLC2A175tNB6v4i2eKdoikBSA
DdUKy1m+9JBi+66rn/LdGXxGIwojw6FpPDIlFT/D4Ad38CzBU8904MIcUW0yTajoegsjaZC347/e
GMbkHEDqKu48oVw1se/FNQipYfAhLhWICprO4ubr21ICeyO2YZGEsMkok6fW7hFBxxxIt6tecPNp
Pkw8oG2SEkoLdIT72mkWqmRcSNOhqKJRHEOqx3kbozzqJ7K/Sk+tAMTjWcGrQLB5npXJTbWH2CPh
AG736Cr5SLnSUaFMoWIy0QfNmxu+cFRtYj+fv81QkXj6Pvx20kVN0tWEYK0+PLSySoVYQ1q3Egci
EnLLSLHym5eIZDRBfZQn+cV0S7gXBBYAQ+72NL55TWfK+5cujFVvbcYNU2mlaLm1gFsGeTzGGZep
Z/YbHBPL8TGC0vxouxBEXjkMLTM9ytLDRkL39bPfvn32OlS7U6haTWgwUzwC+3V1lMnJ5EpPE2Fe
6BOXirXPYiiCzC//pLwn2n7C7vbTAT5umXRUxrOxKtpHtT1tQ7JUm72HJqW2dAsagfY2h+YxWCMt
JAsev7ss6xYonKZTeppzDV992wLcnxkTLel9VvHvcJPtw6m8b4DNBik5GgrbXBF0O2dwCTh3S6dB
Y8KdNpXamoCtOVjY0rnNihsmC0XeXfJqPEQDx6AqaAKoFojbIr5lsAQyy2kkf/uDa4pJbVKu0VEf
r4EtBG978hf5IBpkUCRNFKj4RfSG554pJnh9fy5ZsvL5bsPRe+oYLSBGIT4TjiVqu6JfSAuxfIjo
186NIVeVCms5V3+u8FG83OeRN3c2vLHMVEuehog9RqfnZ0KBpPUG1pKxgKUfiMxgi+sKiVYV/40J
gW7btkMxLl4efUF98wnYx9h2zgzBfSxtZVOQNarcNzU2J4He5E/mcT3g/gSE7fOk+ehk2GLYdfdp
jGHJn7zUCf1QHApby59L2KWLBRVDeEtS5AKzCyjkazEXqqWouLRja+dHCGEBknG39U8tx1xA1Mgf
AXJdTCJxPo+a36eG9uwiLKBAdY+QUOL4Y5KU7rtS0BRx7VSBcuXFflz2AqYVqxX71w7Lxqcrf5ym
Mz23E1tTcNWe343939MYKLAqTrwjMM/pKbSOVbJww0rMJB8S+b84GbNPxRWGMvozPK3kM7uQ0hc/
rqsErLh8f6Ty9rcyKM5vOe8vcTmFusw/cnZ6lagZVnJYS1yEhulyoDWnKlK7LP7C3EtewKC8Mqb2
qcF+P0ub1gywXNoCec+S1QbZEQnKy8QK/kZjPFiyfNDJkXJko+o3EIqxWcCHxRFcuHwmNUvpS2b0
Iujj5ujXPlaU/WqjIMSKRx20RYpU+7s3aJBJG+fK0xFstMSZOSYecVaSDi4bo+D+xcqvZau7yPWw
6dh5Dtflj79nY8YEmAXbTw8ZVaWyPMqqU86NyUXeB1fwF7ljZWZ3Loc40QV9eRaaAvic7/zh//ab
qx6G4NPq0ip1LfeuMvt6FdrmXnwuiJGtwQs3Y6qrybtHpQHaLbgmoJdKWuKC04RVMf3lanb1rrIi
63gELGIszVtjMlcx+sb2kNnJzdBJgxlA9IHtJzq+6sfM6E6v6uuT0Mu04g6q+1lk8s+2J8ry4Vn6
nX+BfWKjMxEc8hl76zCvYb6vhCZxt0Wp6P8DeEpANZG0pb5XuCdtf8GQOXSurRpNmpjmhO1rkLYn
FwrrEBU+2ho9rWom9xNUfDPfkZMzcN3FWDjiKg4zkb21ZgKidjuWF3ve0wn+6ViEbqLCgPEVS9U0
wlTg4eZWkUqk43/ytRsz6KKzxzMVjBa3tiQvgyBKywHqzqfnBgGBvG2Ree5OGwypIZ4Mz+PEN4h4
Iv3dZjUsfha9R16eG0tXRtlh9Rf1VCqBFXjh/csUBeOJiSxeIRfN6xPa4NHpMpOdGMTZ1Pk43IDd
1eFn5k2FdoU47b0x1UbrYoIJW0FLO2Z6cmxBtRlNEXmDRypypfRxYdFTDbn58vGDZnc+hHs+JLh/
PPRCnwHCDUGQK+NvyaN2o6XRLiFnbU9kU6jIlGj5ahQPrlOyzEakqAc/N+CHCleG2XjWfvgCemSb
kaknqFlKOX67DWoARX2xEvZKuuOJ3hDzGrNloeT/aJSTwvEwN7os6TjR11FI2K5G1Bkb0oMJiTOn
zYlwif4D8CCW2tPGLWDqRtNghTcCb+Jh+Ag06X2TqNHFRjOF+oMrv3tdT19pIjlPVtXTC7oCMaEb
wDRGUfkQszGx0YsfsxP8jXTZamWm4oeTY9fgwbyR2n/nItcCttEhGoF3aCLU7eXIXscRTey79nUV
je9OMkbrbu4m5JfM6d1dMgXlKInZqSkIzdV7FCv6anC7uzekcHWNNTTfe4z8dhZ3tzwBQ71y2MuK
Jx0RDQjeWzgkniON9AVeZezNOPeWxgAbzI8iOCDdrFaRvrI/sfHcubg+0z4LAXzsHvBGICIzM24p
+bLKtLpG22TGtEaFVmtKbm9FQ5+PbNdQd2vOLMoaOfyFU3DA6dTPI5QQPmSEiNZziXTR0xMcj8Qh
+Wv008V86KYfCKEQ66FLXxsNm4Ptt04N/RXv3MojxusnwDXA/sUbXcV+PHV3PbR21oHwyMvupAtC
TjnsBNpAM46RHQ7rlS4T+lNfmrM6xYV93hiu7kw2jpRoFycqvaliI0S1KSoXUk387Uzc9D9CdRos
G69+0poRE3Ke0nxNeMn5WijIJFkt0HWEwhme2FynXVh6I8NSG1dZ4mOaO7k7qlDkhRDn79X1vvFM
ze816tlnXPTxp2YICJfzfwOKcmfobozexW/p3katV1C7QttKJGJRA3yE2+Px/YJLprZnKI3aIjzh
Koslk3cpiG5s8nZlX20Tj309SHsd9B9o4cVdGlr7XMRDiWoFJ/gln2uEBaEvyatFjJtPdlKCWWS7
GiLoM6S+FEu/orrCA1UrbqCVQQYmBgQvNrwYYMbr9aPV+3EsDcHP6Cu1R69nuAmns3xE1Gl9jCeK
dX8CzUJVtptE/8JGLJ+uQzbtKRxBhc7SlyjsL14Cdk5pawU1Pu4X4YKQSdrHS8MujQ6t/Y9VjHUg
vYxw16wdC8J4YDRK237IfsGOrLrfoTPodq+tjhBxQfY2p5E7QyJzOLQmuAbaWuwH+WTwe56DFlMq
iYD6zC75q2xfIUjuP7Zn5JG/95WvnFZrjWGu5xcNthrismEM7k7uZumWE+f8lT4UnGVa85hah7LV
sm6E8md33BOVugRk36d5TJuWzXGVMfeC6Ee9eErk96JWMGmhW0DLyYFy37ato8PDJHiHZapsjxF7
BuKS4yDShv3KptHZ3SP2VEdHo4pOSYjRSzCUaoY4SvuR7DPWNr8yaLXWu//BKAqywIU0ftIN9pJV
o4+PdwIgjIC0SmUCGZZ8OImF8JD/OI9ycyDeX/DlBb9R8rThkdjpQin/H0WNUOnuzWkR1qfmkH6y
5txJGpo15JuLrKNcGhHc8cUUbcVHS8q/Xd0FCwv3GoWbkoQ4Tnz2W3km8q37Tbtdy6Bm8yF563NX
6WaFTv6b4TADe/aJP+ydvqFPrLZk6VC/6mozu0Rn1aR8WSQAkik0CI72t36+oEmk+lOSL+4mIx2O
qoIbF29NpSsotsteR9j8FgdzKncnBKsR6+J5o4CfKDgp3LjtqOWwiMqEKNW1CokxBGemqAP+Kspj
TR/DlT/hIE7gnlYFoP3IwAcTPOTzbtms6pz6uFE/HnauKaxzMfa+fok1zjQNn93bmOTny60GYJoI
OI1NivBMKLVolulYtnnorqdIlbVOFWgY3ZxQCQxs1wL96LPSiDKSqsbuM+okWdZHyR02Fjb4gSrz
h8uDnL7yqrXy8J+SCA3kvj7KT2lFq591srixHL6FBSB5GGBrFI9Hizetg2Pln1o6XDOmyWWa2a1t
iRBrEbhQ+6uxoN70ldxuZv+AX+GRnVLU987VUQp6FFvd5cJpD2eVM+jjYpOF38CJclFNEwrz/eED
R1DY3ATzx63f5pvuYDT4WXpnx0YwurIzYZLA9b8qT0Flx9f1UTAFcaB54R6l4pbjDAUSmh2AmUD1
DtUfbYIBX6ZMwjqVOaB18B8A/fu3FFRxJ4CJmprYdFUjN8e/K0pIA1Dg1qBzXeIoktM/lEpg4KLg
Y+ceehdA+EWX89DFXqGpRdIdx5ni1G5NOET5WTaBK5235Hhd8QfUQPm8z8Gd3t7h1swiTcwLodyJ
a7ia/FkPM4APzYtnqoWjumJi2CWclEQPe0/B9zLHrJE2Wbs1b5Vj84t9t7eNR/nh16eaqBgLVnAu
nc+bAQW4SREGA21ojtI4+zH70cb8+sQ98LQr0d3df9BX1nHA8esGzuP6OnrpOzJ0tKVRJwMLRbxa
p4c6mEXhBp7CKrOAEhwOW38ZpeFNOWCqV/dnK0nNhUHKVdhEUgf4fAdONeCedj6Sozc3qwuq07Zk
pWgKX6oELBxs8dOrOLjJ69HaOct1VOvZsyM9vOFLK9J3Tp/hulUi2d7Jl1i4I9uPdW+zt3Ke5IV8
v0QbBGPtqOlGO9VMc0/KchTEk6ZM3XNONJaywgjdOchcwgJpO3QPpugTWzZe+6LCuLaywli4mrue
QBMdemGPhSbpHUf0AVEhuc16jdPXTZKiEdStKbpohCorD8w3Jg91sFEiCw6MJLttWQrPZR4J5MY7
U9MLnUpa4g/SfoDidvU+Y36mGNgsCHfBs7RarKMoV53hPQCUH6tgZEAWa5TRDdcIiAmD8lYM9oaB
XD1IprpvfDh4n4PcUq3Z0BoBs1RvgROcNEu34s+hz0mdKTH7nAvdvpMMWhW1EJjpLbvaLulUA5KU
oFYsZjnb9KpYPUyRCmZ19sOzOoWv5fHIP+O5YCuacoIbnu4f4gjiOFz1Kc6PV+ZBR3kEI5pQP4fb
3E1AXr1ETjkhftZqNyjwPE8Xv69gd7gcR4Jq8H3RyKMhBItd489PWqlpIHivz/qhFBYzfNWcr3Sm
2Gx18H1mMMO4KW9KSHL1oKxaa67Uarim5+B37/OjPCDxd0g4qswdSCrAA5BdX3TjlFXoOMgDP+ks
UgBcYwuTgZBTPydT7qrfyQaGidVLk+csnfRpNzTNYDrqDVeMPLkrNNsqWtA9+UkLobPP9rcd+4jZ
Qz+uAAKJ3poziu2ZII/gl603MoSKqY6aYzjAAoqjqAA6pKesvWiLsJtr0WVwx1KO50TI9CUG6Grg
weTRZ5DXSyr6nWin+/IQNHBvOP1+CUoeuQamozPu/in9qDUfX/f8F99giLlKnaAAFtSi4ZbvCV9E
wuiNJZR4SAIhOcC70gktZp+KPWO+WfaMXMzaEtI/jDNC7KweASP/ILHvN/U4fdeXmpOmZ06isgn+
eLQ5Vs1DaRPvWQG7Sf4DEKFZv2vqGJ0dgz57AsY13kXCwECXPP7StBE93jzERd4mV8fcZ0Mw419K
dTW3yoFUnjhUgmutQCfU+9XJAXnxo2xeK7x7aPfwAwQ0F7XsYZb//PKvMO2qyqdUIYf8TwACm+Qm
6WZ8c1Xwm2pq9NMhyDUt/uF4YYfo/m3kfRqOiA0zucObr9SpYgtIdPAoR0WHTW6rldp9qm4mZedX
8AdZ9mi8qT5txKoqpMYgo+heG1NSIy/HeOpBIu93XFMZGCHu2mdv2GIg+yYZqNCWB0IMPJQ1zZMa
ZJsbl0SehvlAGCFCh3zpaqYGXn1rkAs2+6SimVkb285Jqd24IXZmyO12K4TfUzxFk+TmDz2TRn7V
cZLS7NR4D2elgCqJ1JQvHYGcw/KyEYqqQc0MFIQiTeeSl4aPMWHRMSLBY5/y3fBoTQH3if7l/RXc
y1brmBBPN30wKrf+qfujJnCk1EhlX/NyiUxMVZQ4HOBDxb7l7DvhrkPQJtPNOYsRM6lW9VcXSsqw
efEzvV0zOwOUG0qRwgDyjYN8OVkcRsAsSTuZXtTsBb8JKvHW66eh0ctJtFFOQhcGoxz6Mjqq8cmQ
IM9RVw0JtHZh9BTqOt1iqDntmgLN9aqY82g2gLKMVvDPzotvmFmhp25NuTkgL2aWBvd+ACu4+izm
EGO1hn5QxI84ieG2fb+h+5kUlZSqiKWeQykGEgGrHWLd2rgWy23BHSsJAT6dXRYTCFeeRahqJgPs
cnW+qSMLm2AOkhfOXzr7sryUvKkp4QA9GHLoNJRU02W3lMQ9jg+FhWCERLTH5f8CZy0zVAuMHUr6
vRytfajFXj9AEIqJ6lOygAKml1r1uw3wzcuwSLMRsQh2+E58Lr3Lyen5bD68PomaSk9BaTI051mJ
CJ+nqh46GaAufiLN2HxZCzP7TfhHcucJWqqiezB08OJgX/1W6gpB0aqCdOzupYnbjUjnsrKgFS/c
C3Xtu4tnJYhnWqcQfBM48ZinDTp9j5DChluulNmLW4f810i/vDSt303Hkf0+XQy9NP0adXBmD297
6vomTVH5+WUSG6cMoagkeuGGdsrp37Nj+gmWV3kCeC+3Mlfj3D4cc/XSejvtHXOqWv1wL8R9Obhe
87C4cZEBQP7OZQmssPxk642BHWPseLAUdae1mOdAltCf6l2p/GR+VsYeGoAUGGRjm6JMn0bx1nx0
DR+EWJWcXcrbNDlyv/xwWEJDq114Y8ZSIiDZHIUxuI/OtgByL2oSYXZ3+uhzD1yN/topHaeJyxHb
mGH2iEqaUWhzmqxJCihpoqsdjZc8ZwTW8XDaCrN4pSggWEjai8tjjWBzltTpWi1Jg4DDYw9o6osF
Znp0qDoHzCD+6ObfPZyqOp4h1Npb2OqBSHb50K1JUVOUarfAOqF7gKvBZBQ8w6/goz/bDVGR4BBQ
jIKGYFbEFsbrzuG3GHdum0RlHH5gTAzYR061TJ9G9A3Nnqpj3T+yTCpAVqU5wRoWeevnrNlWp9mZ
DStswI+Nyf7Js4qv0wCZ+41RaW/btHccsJ2ga+CAqMRC4yRdfaOdtif4vECzTLiJMDBHsRvTi2hJ
igkDN+/lKYgbE22XJkBM/79RTkR+l32Miqm9WA2klD4zKgtSOzsWFfDAMpqMQ+jZZnJM4gpNKks7
iA+7aP3k+dEWNuw6/1i2BjGAkH36SeDiTw7yPulJYeKgBU0ntheH8YpKyTA2NXWLRS/DffteWqqi
BImSxynZOQUaF8nfgjIOB6sVKvLhvQgT1b2r6WCbPjMEzJC90HtBF4lHgdTBey7/ZL32iZvax6ZE
MuoQr6zbv7Jm3Ee1YDSNDIU/qGg9CJJzWQc+z67M6MDR0eLIQYJ/57nk5wXWNxqdAdZqhFs4XvmK
KrVVKFsBo+b83fMUDDvYByi89SdxG6Vb0UpkPTGWPRZJPS+XwfJlncoiFe1ABitAw+r8THTz2MMN
5HKd2L5AboUudmadr9yDh6mbTHhGjY3AqgndBMphLOissbit5zKAVzGRuwPsKCAQ1RaJhtu6JEG8
NN0nHzuD5ZQBP7aAJjzcomOssl3buhbJT4B0P2RSIq3SvTCPcJvoYqW19wjMURawt9KzcAvmbMAa
Fu3ZCHi/FCo5SEAdy9mjSj4Y96BP1GbrRtILuH7rjs9tqaCFVgB/s/FCSLUautmYp+rCVUsbeEeN
OWlfJeUHl6fyhYL3unfxlF3LmkgUw6f5qCYmK6KKXzaq5STOn14yCR3frbhNkc6RRHPaEqHAeaQz
g/6OOfJZEtwH3VXy8sBC3CK4klc+8r2O8YMZt3Xd6nODIjhjUnDxp5joR+N1VvzqoOPbGQzt73rl
BjVG9qQMxRJEWm5cf1TmQxp30Eeic3WpLr801nPwoGaCho8VugkysH47MS+ibUhlx57m/QYEz/0n
AO6Yy97su3qpO84tZsQUX6ARrFsQyPaF7WCGCY1qxjdaSH6bHbBg7Pidzeu02qv7+7xFn8K8uD0K
16GExz2aWOZnTmaI3VRGFB+nzfOe1WI5z0dHuptsd04p+uTo22UZwQEsUiyhkkj6a2rO30Gm/qYl
/0s90506266mZ8owDUe7kOsvCX9aOi3Q7MjHzfERGau/0JNdJZ8Tpp5HQjY5OlVPjBYkxEWeZh0E
6ZCT/pg9lly0zGPXL5K4FMNbXeHYJSLRtdH3qAV26OqTowo5/WMA1FrT4pmzUXoHwGJreD4p+VMB
0A0YZkRabkGkN9jd3QQveWSvdAeCKQalBX3TpQ1Z18oSM3LLkzK0fdQehv9wZknU7fRQAq1k1/tG
KwRDgro6TMtrr7JQXIe9UK8XfgvYcW1Xjkg+it694DmdxcNUTLMchQJbilyvbCzoFKqAgL6Qm7rt
s/qcUxJsxDZDvbQ7r92zKlCGyIgat5NNNe+RFzzOs9WNgWifzrizpxAOg20ag6ROSBtE+9ctz0MN
a4B56bmkeFh5PlrZrsh0aSVaxKEOcg6bnsi2gzx+KH5HpfBoLgPdKfnRGM6dmKLg6ctP/oMvhk7A
Syzy+sTZ72MZ2bmLQPKdwfDEHKchExZyGHsi6bl0ixX7EuYTOmgcHGhAQszKlEVMF85Xcuq9GTpq
z1ak6HR/cT8uzSFQvOJFeZwtxG5OONXx8f98CXWmnCg9/LxEluxFLk9thLZY19f9OuFFW+spDOFe
V+YwtUW4/XWQMkJJrWlkubELio6xg3fY3PHx/pGcACTkjPygoJCh6ylUdTEN8QUl6Vj3PY5B3Q36
fztUhRwXNO29CtZLO20yWnFOkhJLhezWpU57cBL5g9ad6+G77idf9bIeXmqq8hO8SLvQNuS73XqU
bpH6pmXg94Q1fnhZV6NQwbjF+yAg13/m24o02aMP/qbAF9fOMZbDi8AY3flFzUFw18AJjlTDMsO/
RY9GVEkM0xNf/0B9yU1R8xYH+65Ok32Qy4eB30Bn5824fcd4jqCnJSIUQQBHwnR6GUuyd2/h/y2e
b8s/BH/+fX/A9PucFx69K+pt6hi2Gn8MQ4vNJeDN/ES9kdpz83BZOf1r/RJ5GFDE61xAgdfdCJgg
ROrH0/Ubj4+O+5XuFoIzKPIHEcIt3pZHfzn01adoMVNknE77iAKWRPy/p77T4kakRrjL8Q8JRnPg
/QNJeKCYto8FStc8EN/VZX4Ieu87XnxkGvQY/kQJz5xPGRiW0oajcg8qpTnOypKpfHfcs44srkWi
fzlrHtNdiR97gDGKTjZLkwNzK1VI+G/tsAQpbFeMpD6GQ7E3ehfvLJjO2iQA7TkL5idQMoI62thh
/XZwo8QbdlQ8np2fBhBRaiYQv6QphI4fkO18RcOwXZg40rbhsusASREvbp8uQBEAfE7sae507/FT
eFktbHbpQ0fciinB9bwBdlkqtpxbx55MGUq0ZILGFqd3vze4Z/QcxhmXfzugeCwZalq3Y7fEBfBg
ykfD5CAzAswc0q/1s4tzwMJXpE7gzTHjUIPe3oqJJIPnoCSmSBjA04CpZsr/G9zh4s3vKqxMrXlq
RRkbWND/8ZIGat2LrWQ0BmGlCM2z46vVzO48NFoEONjeoT5cUMUbxuBIMNppZzfTRTAZcVKekhmG
I3r2f5XKbhtBQXkZHbfbbMXfxgrMkQ39hLRFZ03hP2WJfeZ7ql8pOF+XLmpUMGBMfCFF01+DAksc
uAn4l3SpRtzrKnLWOhPnCgI6t+3fMLj6WFb0iUc2HJQNoqzxGEk+KnRe5nvPKcr2oHVSM30npwhW
sGXbtCvY0XWo1xJX++18FKdAxNcT6DFyXFrpDYe7MJrKw3VNdH3WtAGvTcWFETee8lL9/PiDsX8a
dMflFbNIhVSJ7/4+eKRhY2vOdXwpnHh2WM5sydi2p0q+RhCcW8ufxqJyHHmDtGGim+LmArIRgU10
NRSPQsR4+4N8tr3QxcIEh+UnvwPT+BOd0b0Cm1R4NBvFgMfRtSprHWuwYZQZzoOh5TLMJajehwmy
vzFvusnQb1MyaUJaRibFuAJoLqqNr3MIW/M2r9Rwg6XUhwdcPKW48jopi0/MZU5oY4E6yfbCcRPo
wVUmqM+OqwYNaP5ZV7Wv0yM8GsN8Ir+j9ZIf/Cj1Xs2snLOvHMLhvAqrGfKWa3uV53ZwqEmG1qGS
ob+4pCgBzf30VIpw+yzvCM0cWeFZaQ6QcOjPD7S4tdlYDO6Qiiabvj66gIft9iBSnDpAKktjlOSl
ftcC6+Ryan+8HpYLR+gwNH/3Vw6CohF5CIDLdUtUS5sF20n+UKisu8MXbyf4ySvTCatu4cvdwtoM
N4X7PD9ugEaT+CdwoIoC1yaJ0h4k5NiKxroUDTBWNUfrz2kHB1GZAlkA5uSCuuuXwVlnrEoteTvq
YQ2Mt93dL915Ewl2syJlrbsIhLmYdInk0JpnNpGzbv9/crr/bGhJWTtsVwTJp8TlVojTRYfpLQ7d
f+mVQGp9JPdMgisFLakNAm1qxwTFYw2ph3KvBV66teu+TOtmbeX8CM05O/0WAnOvjJ4auE5UKRwd
RbRqeXt9rZY/I2OEXLNF0v3gCLkfMgij7w0W1ywgv/7d0Of7v8j90+4Uq2rv3MSwBYb4T8mJdpe5
k1HN1aVS80DxZnGBKTG3KTBZWfeAruF5UU0t/2wzKiq60gdJ9cQ+glLjRulSKprPrGpkZQILqVD3
UrGot/Xiq55e55x8yE5N6wSNjC0tX1Xf/SFqckrRizeh6ohxqow9gomDQUltgnB6RZgiYvTGzUzZ
zRNXJqn/yRAugbUl63kv4v+gtCc/MD6JNj9LYvDu8YZIpTqPNWj4KQZRLECDIFmsL2qwt/TAjgLq
oG3f1FpdPOCBnIL3QOW8oIP/L/AeOg/yB/BiyOdNjysiHAQ5d2M3cG81VWOrHpDv/dOw8eEFLIxF
wUIVuDDL0re/b2vX7ASXrDy6lk2pfU9MlKVZh6CKeNqgfPlYO8P7Ao75aou8kR/W6KXMuqpgtd25
Bs3qw9LY5qNEHumdtpQFWOaAvBmLEfhZaIUrWXmuzp4IVUFdgpn1x90siHuJyJPJgnXE6DlSHsWj
jArRxx+Wcq7yuLMfUPMqPviS2h4Oi5G78OjXSmAFNu7Wc5Vqi5sHSURR2TdWyfQqiFc7aTgT9nz8
SCNvU0bp+ksdonpLLSb2MKMcakE3F9DFpPoa90W2JehEVxsMgkbCC54n7SdJ0EhDAC14iCAkA+Er
I5W+PxEfnA4JFBaC1+CAqQCzJRDzJzqxpwm8qANNul/qib7ydGoweFmVM2hXFnA21xwdmzEYPz/K
0Vwyu0FiPszES83T4RCOxRkVaWiP2Zhd78E/AKmJ/fKufeXzCMRCxw85fpHUy4Z4+kvjQfPF0xee
Q6/T+ncaH+8XuSIBP4IXqMNgx1GdsSlPKfqbu9HODz/+bZo+M2WXVnQkSuTXhi4dxxSQqjNu/QJX
XZBVK4k7sEfGsn1Ik0a5gWhr4fA91fCVrgEbecBY5YToSphW5yh0BQthm8tEHyt+erF8pBjg63tH
RCSMq2n4iMl5yLOajtP24sEBESgzvtEsczpG5jZHpM7ZULz/pnivLfQJ3nQMnm6E50n3Z+VQI5ZB
lI6E4ZKnk7oYLerQzpb+oQaL2eCp5Gmw0+macpUs7tO9MT+rk/3y51lIABgqFUYGnWXgrOe6rsoX
AFg/ysFEXmqJmhfIKfzGaiezRSlqn79FZaM79EQYW7vmL9zpTTbE0xNIfA/boPsmT2TlZnIThAka
Xh1CyKsin5LcBlGMAQLQOLpWVIBA1rVWII/6ggAHZziZwr+/VqJad2/aLJHywQ00EvVlainq+YmJ
hf8UX7DCH2pfi4e0BHQdRguaBCIZUlIotqKyhv5rQBxcUWVlls6TCTCbfvUHS3xRA5HCJE07T/uW
R4rU5zzAbEZ1ZgAOkcv+GO2iRdBHZPr593QDr/SMnJUDdAksHpfhH7zXn3LslHU19WybRlfUv0sb
+vE91p8dZgw/Go1dJjCt2TUWmvltb0M5fDI+McAQfvvtLhUvbPekGUBPcBUkHwSWK3/faSVeJILI
3D9fBlrpLMi82N3uHIhig7qw04xw6GLRBcCjip4TQeSB1Hv+vMu/arS/953cn2u2Yo6S9PszXRLU
NEXHmeqh+EDk8XV1T2OAJRgtvGy+ilT6j5t+lr3p8X81yPiGVaIILLVR7NnxWgEQL0cPZodIlU4v
WLaIffKRM5njDFJ6u2u/0HICPYvJeOlQXdULQBCM7bJJuG8lRjfkt1QqP9A5DyXsxhBzpr0Ah1RT
FoStLnv3H2ltumdHbpXIh1luu3sjljL0ccblSNJ0Dy48edHPW0y6v1je2vhdO8MYeFrXy8Qo7j+t
OYWPFC+QouGAN3Fx8985DA0iEUgrdgbyBAzUkERhdyT9n+AM/GboFSvr60eP7coi8z6KjvVa0xeE
LqxH/1qziynK8w//ndx487qdAEPd7+dsz3I9q/ix3+AsDN4ArAB+UM7TbW7Bkd1zX91kBFdcmVPR
JczQOQyLSCI5GSqtB16wQqrbNpnBnflwjTaIKOicP+q44U0S6ekk7VHVkxplaUHWygyQ6mFIfEUA
2MKQ/7KmB2JA5XNFUdVGIJENeMTlnfciKU62JXoAW79ds3U9Cs4EfpuhHMhj9LeVWve3pKbhR6eC
uQoXmsCZiVtnWnAU7TRCxNu0kI3AKJbPmN82klX8Kr+9cZAOdKkCVQhSULAKKTnYSD2pLG1UBQ9Z
TYGrCMBhMkLVvxzm/rtxiCW4oWx8gC+6BTskNLZJ5ZqxrlQW4TSmxx1dcU3MV4bHJ604Rvdb2fsi
j7QkXcoYeYn5RkSN0qhxsYZ4ZAy4P1SmVXIwXhW7X6puHgvRmuA4RUo2u1WXkpJGnv8eT/NcM2RU
qeA/R5E4Gvfu1r5qxVtVlkc8CL/89lGgUk0u0DRSP20aBSUqPKxdcJ4En6LYbdSQvgVa17V1qFWr
h/ifwwAfX2lwiHiU277z/A/ntEE8PMINAWhX3FJg3Er+k2c1xW2x3OSn0YrRZl/4fXBz1vzqAjrz
DtNRZ+YbNREP/klKXSeYPiK5R6+fnIG8xDe/ZPe8SyJr3lJUreSsjJz1dW2sQuFydlK9r2e3H9FM
qGsRKachsLkZ4u0yUvbEBo97xavodZiU3g5NpkACASntD9X54Jv5WFAJHvPYJQ2h4/F3k5wx5L+o
7gO+QZlRlIoXAd7bQtlCW0pi7b7u2MaxGME79fnFsR/GtfRjMsa6sth8W9e9Ne4SMmaVrbi1Abmd
bnCsbYfdsvK5BZBdrPI1ButcRvck7WB1WlwYGVxIqY6lbjxuTRXQRmnXXKpylDdVdVT/Us90FBa9
mPVTA0vSFiXzK4E82v3FugwWV16VvWXqp3OGBprLwpvrUbkdghjj1K+azjSO8YnGEtZMVIZxv5r0
AT8+QXtBcEmNumkwdw03g+FC/bSd/a0hQuN/qdD9oi2rDWZI9eDo3rSJvalqOyWE+BTKNv0ahHQv
TD7w2nE2mvhPL2mD7mQFWCTr0UO/FajzDLl97GoCUE8vZf6QPUIM1QDGcD72f5TULifrcoGqQaa4
TIBZ79aqfmSZWC0PMucyRqmp15yMO+wptKsvgCIrrGfF5EFq0OKlxC8kWAo0KBNjQN1F29Rr5FP5
1eP5GDBDbaQ3LMG06P3M9apknSjG/vXPMs3edAdH3MuWRd08SOecdhuAyz/jkcyS9ggex5BcAjIl
1xxIKLhBlW6R4sswDi4ZeYCuu8CLd3gN3edFXNXpxOvUfJzQrYF95qxOrIEXfpcviisBWTLc94MQ
x2KlqBn7jFz+iy49ddTUSlPvjkCxIBIVwNiZ7jUxLKp2y9oA2gC5OTelBgY0hxC5jnwnSTooAtIh
X84fb3O6H7VWCmqTvage+V7vG8aitAsKa9yKOlikxEXwI7LcOBYQlZnQBKKDM4AUDKtHgIezMmip
Zhq5i4e7sf6BraPM3rRdqfBiGIYwO4G37NgK4VAT9nQX6WuVdDlCS8klYcYGy3L48nUYkmTr+1Iu
twuf6fST7k9A6UIW71E9K64+9UZXKZGBsI+LTbfMHGjAoccGLwrXMW3TEk/OpZXLupQBWr6df7/W
M/YTKwmitPVjmmXgY1cgYYcRy6Bli/uv3iTeUovnmhZUNtGB96dENSYOmI/36ginVjuucHeWnDav
zYY01SBwUWcAq635M5+RakUL37UXKHgaAYNKe7r/GmbEvl9QIDtzOnKEQ9F0DN/kJhubV9Sh390h
Bp5PjJTwikdgrPoFb8edPCTssyUyE35DMPtFOrMmeQamhyOXjMQVYsTR5F6ki7KVz908HlQmBwwI
R3SAXuHHejznAvK3oJ2YKXBI8At2gQByYlSitLC0fWZfbulT/V7oeovN18SvuyfaRZ2j5tppgLKX
TKhYqnezr1PIx7q5CrPy676TpP/vy8UrXY0xjFUylw/3LR4ic7Evfjjj993a0jmUV4Xs2mbiFuHR
65HX/Kr8U+BrzimqCnShGwBJ25Lt1RUrwr4dBy8m929Rfb83KW1XZkk4q+hwIYhhD5ZAvdLovC7o
J6yr7NtIbEaJSsGcGJ5nby9LoTB97x2VyeQb42wcXA2shVLqAZVgOO8F5jUSg/CItgxRchIWsGrE
BAREz3c+CuuleVhaTTxvg5KYogL/DQ0AkAyjJac9Sq68FoboKD0dpRNBDo5OetUM/CBg+qik/Znr
Nkxb5U4dJ9DU7Tuw2S6UUL1Dajg208YEzo275VEmjNQLZr1z4mtMtZLCEy395BaN4ZOSBtX8ZDXn
hQRpJw444AVROowjVqhn7YnRIJHoxtQpilwLqGgrhu2sJioPQHGZioTxo9hPR8ql/WSGC+67yx/m
DL5YwGUXlp56QkgwyJNJQJ63zDI5D5hipjxDheXodaj/LIF18TLSXUOPDUTZo1NNO4iZkYc7AnBZ
0v4WakDbZpmeGrXHiUTxwWZvx2r6NFj1m6o0SO4KhHsg4jjb2o1esBzNDyyW+CMYb4De6rvgA2x2
g2C/pTy41PX4XK4W0eaBoaFuPaz5nMRWoWnWMiY6wVGbUCIiBKTyM6Pos3WX6jSyOLCPUpWtm8qn
sw8esypfYPhXuakk8LkOURY9+hYuveRlq9uRsXihFgqUZLghvfS+EoNB9Ze9zvQ03dgQvrxP5isU
gUjGcK6pHgxrn5ymqHujimgnHzcDkPtgUfzeCcMGX0Causop3KmYZgf19qhFaFuBbjUcuwRVZk2k
WUAfoej/OvysonCa44X6ZfVw6Z6EsedZGrtgUJikJDdLkpIXLrs3YyBQwi5y7PoEhqPy4yDPCzxj
b08zl6OK264G7mNyU8ozyNflGEYwxc9l/Z5t2BJP884cTdUqa4iPHD1CiG3nok9qGFI8BL9ALglw
GGvEA32NLqDNzZNTslAf+mXxnS0xqNu5Nep20UDYl2I5trIKgXJoZ+IBaAr7VH2RD7h+/ZuuovJr
ecqHQ9RSm/e+u/KTgg5UbbiGcelxjKdbtgQ6lYozgaOqzt1gRe+sgeV/AR7EIPtuCCbYQmACcB/R
ZoAFR9GQTx43PEs0rfS1cTRTGBfu11asCax0VqevQeJaS/0ykLsfZdVIqeaCb94i3lqlC14KHlx9
QCGXZvDTo4yZf0dhxQNAkaFyigmgmP9uatBFDjaVowwvWfxhtvgfbV9RtfJPDiRKLwgPW2Cs0Zpa
DKa7iORysSAlBJMaztCXmv/IGcIbXxV6fcMkqtzfPLxSD8fXpGZh8d6qbqECCFF7nnXt4ZxzkQew
MFqZu+Ty9tBYKzNK54AVQ57dXf+9F6unyMd2qY9DeA6c1/EwFH3P2g1DkwQuftw9d7d1H1klQ4Zg
IHnKBcInuyX4kC48Vkn6hJl3W8h1jicHXqFfKMRKCrbX2znKXOVxs9xguWofDy3QCVJoTXdUJG4Y
ZXhe1vlLY8tJLHPfmJmHvQWrODC7lddU26WSfmDmYFIcP7IkHufw0lCWBSDtllFdv1tKdPCaoxS/
YJpFS9xETG/gWDTJJgjV1ZGPWeNvRyq4AO6kDqpacDE3jE8yx720dePoKZdV/+E1Ahh/kFyQGvr2
meL3LAg7kE7YEqmUHHy5fDmRdulybIWkqzV6at/+0hQSOlJCVzyC53ec/qI2hId2XlcA8iY+iWt2
UvZhm4aMHrMf2t8Lf+w/A5jIo85lzrk6v6YyEt5wljPHKSRP33V0MitoLx/cqdU0e1W4aZigmcn6
y+NdB2AkhJjwVhX7mjN1nuAGbhwNZC80CAKDhsOG0geeirNoIRAiEUxl+pXN1O+BM21ezqsyP/om
esWfkWo3R87z5gqHFTLdZnI0gxsN/wH1oaDCabRjSmwDhSquhsPEmsFlAzXWSfqzu6WfBm3e9+iX
BGk/azU0pQfW6cVNt1+B90JadFOeTM1dF/zD0sFeyx99K2B3XwowYeZgVObaV00Uy8YRtMcMa4GG
NdIUOcUEAyVEvqR4hxWnq8XCt5vAYsDgqwqhEnnAQNs49WI0jnkPr84Q6n0DMelvSZIhA3x3yzf5
74uwjBWeIFkScMUYVRwEuLxe4ufiN3ApsfQwNpjVOUWxTMuQcPCvhL3LwEeQp4SglO+pO0r8DZ6g
TSzuxDsmmjFxly9f2UMFlKt0yVqrcsksv6yZAnJMLzOBAGCA9TKeIqV3QAPxoibSXDCRlrMYBf2B
vTrcl7r53IrWFKoschWwO59iPCr7oEMUy9b72XnSmCuMnAGuJtzrBuIg1LvSlEBvXNfVnxzaA4eM
//YI1VEBkpU5fzKtjnQ1BzMOg+rls9ZJL2KocpCWEg4e/oAvXEtNv6b9LTg0YgW5UpQxGlx8TBb1
lBryeDd8OcxbnabFTpp02UTgaNhszby58NkbE3A/Pkj1SSEcgH8UQgCqjtafxXcosi/WbWnPTU29
ncfkZWo0qYDTP/zQgj6PjAIjKmtrYweWx9Ui2HME00meFQtb2PB9EwHdhYoWPfBiFmhRqB+f/G2W
T6ZZDrzTO8o+c/2RSMYNEA5EUpUHh3ZoL/VH3UK8R9cL3KhDGDdb/m7b8zZzb01zIgwOAVSS7d4S
jO0kEckq1neYRiwaJBQ6JMntFif8Xg6fMcCvwasfmUKWeCUnYbxTvrsIgVd12WFeFI5YoOTwSSVu
MIl/saTAfhOVfjaQQCJm/5i2dHe/uSAYAlZ9C2vef2IdzYDHC4J2YcbE/nEMOzbt08BjnC80RR9u
yHYZgYPcpWZcpmU0pJxr3Ab6VEvpCK5fhVUsH02ygWgzJDNZ8lBUkFGcOMTEA+BDnZHTdVT8LENY
ngEpBJzOCEgs8tSd3jcGKwynCsn14Ek3muSZtqz7UmlN4TUtWOKPzHvjPYF1G9uUDVudjaVkvBJi
WNgKwQgIWPdrVWb5nGksYt6zfa8aE7aMPvhZ4d4SrYvo/iaqwBj7V1wCbVs/dyScSL51DDA3F5Yf
3KqqvOa/GutkSUnJ+p5WCIhD0JFtnjarezcerMKB9aenGBwlpFQmFPRj7md5K6RD3+FP4VCnJqx6
FTXMoVbHw3TaDPqyyUY327u8KXp/Ft+F2accSSirvRtYYnfjrhe7I6jsxYE1qs5gMCRO5uCNBuke
B4tLHPbDofdf6m7YZo70WbcdA+nFViluJ5LN7Ivnh7T7Cy53dV20roy3kZMod8JlEacCXWVF81yO
cKFsXj3d2rc4d/9B+q+lb8bD0DDFi92bLIGmrD37fbI6WCV5OsOkJkTCDxEpB5C/ccQa1yv7/mJS
1YOdMzJuaU4R2E1n5upF8RLlMKVgXnnuvGMrLcmsw/1uxkzNR9IFSLt2XmvnYmWw0CKGNdrepfNV
437sBBrzKGQawTR1bM0QJ5LTRin3Y4CI/kNzO9LkKzoz7W/nIRA1PCEb/AYhYwsccSzg4wdpmWl8
kSX9pgkTnWnMMEKkeQJH9LY4D/uC5b0P3cs5XDzttI/gZL1ISoII++gP5D1kjlYWfsT8xlasiMvO
GXtkb8kA0aO1s35QJNYkYmz3DopSezRxtIi3dilYcJceRcfKJnmr1x//SAQSGWk6Ox7DlpumauQv
BUHI6BVKhZEtaMFBzKSf/moxpYf3hhoSzgoYwkttyhcyyHT1F1F/iTMIMC1fvwpVA/92Q6A1hV9E
hEmHIj3nB/HGnPPCagkYb9sq72LQHvYe8t9MZs2J1XCXT6f7udSI2aPC4uNpldXa4mjbUelnQdq7
1reM4xwvlhg2+j1RNDuDh13HseONaBl1xm8BVs4r4/wag7h2nL0n4cj8xFk3E/cVP+DgCb2mlNT/
hq68qKquTdEdnvw8NJ6TeTBWrByn9I72TtipbXFQp4feEjBTAzana2wiw0ONkJic2RzLxV289rGm
f5VqHRY6t7SCrvKsVYqnPxRDnyPtU7u8A2aZFde0VWIKyTCHwVcjg8SSah/mpWIR9kWHhHszGelJ
i/4qPcLg9Yo4E35OwXBlzLyYKxljGyMx14iUX5cQ17KzsaH1+UsUaSCApghaG6F2wsOTAnWJ463l
GeSBiaC25fXFIEK82AaLLO9ADQL6TKIN8oTQREPXj78UKSqI12WDrkyg+6uktf6mOYf8qcv8ry4D
kLeZMy/ZJRQ5Ho6twJYEPjWWBsxD+3QJ+iqv64Fhc1hh+y9DpiFuPFTsxE0MHDWAh5pnAEXskWJb
sp3FWplrXJl3g+dIEbJosbk3cqJW1v1jMqpdEzifYtahYqx0Zc4bjHEHRzYkTiAluqi4ChXS+T1J
E2S9h1aSYBOZQphHLYJlyuN3oRyl7b/h7Dhnerwzd0NQOySbE5K53y2EIScppDPy8AbhOaVTjW9O
AB8eeCdWSfbqb+n6A5qkZg/PX5Y2QwqhyRJJt6plhQeM/bSmR8nkWJYuUuLDaLU5FfpVSVe8x/U/
o3LvV0RQH+iEiljTNGmEzmAL8e0kdmvdN0b6K5Fhl4Yjz6MTmv9209xa4Gkx8fs3d4r7gPDrrSqM
lLnpd/++VCxS/2aHRbLkngGNmw470XOi75V1Jk053QZ+nMY24Dhb4I1AshaCj6oztZ3nxJIjaj+J
EBxKK5qQFfmDhy5hXvXt4+Jn6inVBZ0CDDGGfND1YnXdiQvSaV9eJkmH6As2b4xPfLCdrG+33CYX
4dBOptBY+iDycRRosZbMAOpEbb7cq05tNCa7cQvczsSurlmVSLXMfZNxJV2Gkn41QvSalUAIP4SW
AiCDxZxO0tY3alZ9qaqZL8ROuY8RvFs8/BIaPaegm2naNKqJY6TBDh4YV0OwAsEttHn1SYRct40f
aa1rc7T/syrrQ2BGq+fmjoiNf7RHmBpiQ93wO5FC+FFMMfSVCBRekePCP0PGWCZ/E1+BXDxTTpfC
UpL9FJZiT8MR5TxoF7lbWD75TuCdp4H19toxTsPVyyk/7ZTlAtp7DEhR8Ue3pTIFFp/I0OwQMcyd
/S3xQb9czpYyMquRNIRtBm2u7xw9qALr94HpwsEXRDL+QtFKn+Dn8HfMpJ1I3px6PseIIxcGRNFD
2NlCq/QGSKfm4FULQ/orfFzbqOmmzqL0KAdi8rzM28gsFxSlNMmmMyVRBTwPabju5EP/FBuBDD8+
JKVM5tgqym+tKqZ92WFG5bPgvRdqWCx8X2YBHV1GKWAflfer8FQGLF1lOW/HDFkDmEejWV1S7pc/
6jxlAXrjWYfjazHT1rdFK0iqI/bsBsPW2MT+e+P7GVBi8vQyGGhyTwzNEn6Z/8twpB9siNDxrRdI
JziU/+BWwpS7r0IYzZE5xyyYTfvc6ZeiYYK1rZHYTQg7tW79qPXrSQbuAyqKhU0uQBmelwweqdgZ
UAz75TeBDozUmXE6E/IbTmQI67EXIbVrGfxESTRfPDHgTaWBgbcfdB/EcgdyK+KEn0l3kJTsZNbS
5O+SJPkHod0MQHaqxECjoATlrm60otYqDIzKixmeq1YwOL7ljvFda9ceyZTjlQjt4p+yVb4NQWgi
oIxlDKVb0n5KFgT4R9xEYsYrQLwe5GgW1UoMKd6In87bsYViWKN/ylybYO/U6ZYhvn8mL4bLNfuO
j4dQe7HvJyOEqjEzTlvdS8ea0ygA/xMPheB/aRZ01FxLs8FRS6bVj74EZO8jIajVMGSKOEHA+7lY
CnZcx14lXKopCl4LTewApEP8qC4YTTbPdn1h+32/e9VPTgcEiDZW53+Zr/naoqku+dK4uSFxNJdg
povZHepty1Bh6JyvOrVGTIS1UM2mmUjiQqNQeiIzAZDugeyBl+JSID9uDA0YfZ/NNbM934KnyOw6
lgQkPrlPV+/OqLPkh7QtSoFVl8J4WVBIjGNBmWpsPPZK3xj/3zi4GC8zrFee7Qh3OKg36UHF9P5a
NVf3Ltnm0MvexWPSSqhnzj/x5nbw3jqyOuaUXnCdiEaCiNJH7Wew0lMCzc1l10MyUlsRQyur0p3j
HIHyKMSNx3Hhb+mlhpEVVGgw3M1AafSAZQBxKkdo0d1PtjRVV9PFqS/6Ewpev5NHcqPPIH/nQKLS
pNxtDO4UPyODdSqKqO3WOHzZaKrfvgaCrCTDaXhcV6qsZLZxPGE7M+V6bbPtb61hpOtY5XAF4xYu
1mRgeAiaIKKogX8wdLKoeNQV9eU/6usorc/4WxFNyRLgd6GM0UyW2rO+uPbgt+DJcfZv6muOZQgw
pcmiqv/CYf93l9g+JWgRjZ/kjhxlsS9SheA1FEI7GgVv+SNQEQeihuFtJ5shfoEy3BopOrQubQvn
7RWVZKgOYGVgKqIUscXSzsh+XjI1Uv3tPtIecd9qBWAmqgIYiRtyrcXbUsBIFtF2cCsR12kleZGs
s12k+QSWRt6Pen9BerSsZan+FZhhu7NGU9EDgb6FWOtgoApf5wl+fjvDMA/b/4J4fmFWxn4QDngZ
Lq3uNaP5OjzeTlhbRjqhGYsIBluNIWgg1h8PsN8MAvawkP3qk6l6/XrdpR6G5OlL/ERWXTmwM7wx
jGPgAk5Br7xn9gTiQu2xdxjgNwmjRAQwn0Y3CUlMp+4iZTQ+k2iBiZruLBh1YYP/F4afVmpVoDMC
INNgrHLCEfPSF8ZdYVSCo2T5O5cky4hYRLrt7HsHn1/JCqbI/wUCFO/YoydVNdeHw003/91TG9O1
GSHAzznqXMo9/iaJBSwLaKIMat7CTv0hyOtJaD6X6JZHT8rE7KfwUHJDUOe/d+j8xTeTZSn0fcBt
Y/dBm5ZQ9qUN5EKhLyuMvptmDYaUdgRYFeiHLUezqm1d3xYIbCNRq4pOtOtV+iQ1OQMU1VNRu38o
H7QrNiDmZ8JJJ9RrCr16sHanVIg5NXnO7/rSvH5IDbHKfXHLXvMscu9+jgPaE7uSB97cCbBj6RVl
E5z+cFo2qGnwryNJ0XPxU+JbyqvOpLppxs8/UY1Sk4XLUUGlm8xEjpZ/jptkb8jfvtzCVeRe5mAo
+Cy2PutG9ThX54utqhq+IZg6mREJjHqfUrtrZIxo9tKBe7AoEOZkkCP4yGhMMuw1h3p9rjSEhCU3
FRnSkR6LnkM5TiNOORQ8n0RNciELHOzta6AD7T9RNRrRtWew/TViD2WOCQlNCO28qEdToXtgwLu+
2DDDb7cRDy95vgp8xvSjMmwtwqorKnyeeOh2baibUgmkbYzcL/0WQaX/LTrzQjRjcjHGksz53BkT
b4KRh2Xrt/lSMecJ78YHXFeSKoz8CV/s8umsoxcF4rP0QN13AGpXq1UtV/pTI4YNSmB+kvzBJssP
HlJIc3J5SVds0PWGS/srJPittGvsV5wPRkUR1EY4GpumSmkIkby+4cIryjprmiRajlsuJx4JEpBM
SX/Zbg9TJXvPGN0zbdk2uYUwF4CsS8Fjz4r2WoxyRoLARIkVA5G6GTcuwFLL1ScG8szsIZu80mRn
KS9FgGNk7XAvk3z6v3gg2jLy8lHG8POkzOSQ0A//3B6932yvGkJg0SehhfY8P8fV4y4nbqN3ZFWk
WAOOgoHgQzNrAe7kb0/tvr+YcI42idjb32B+vq+6SooDL+dJuQHhMGmjKX+oZ9lReJrK2DjqoCPB
+J7o1j2K0WX1xa2VBy29bKiIgv20+N/ddaS1nIpZLMkLct0z0n2kgtXWR/1a/pay9dFHLMaB9tCj
xWfIEH1A2/n6AUYiT8e+DlSV5PC/iUGkRULOR3LF/eUQWXA4t1AekF1MJj4Su7bA93at9sZQPtf4
eNn8uBetbGvS7IgCVqngHhscd/prs7xeDumynT2Ni6IhXWo1hbYmIf3TBggk9NKzHqWuiA6l9bLa
n64gYSDCcqJynV/Pgsv2rkuqY0n7wzJMCN+4fSRGLNe/wCIDOAlVCjLzu/S/FAf10G4CHLcD3+vB
zHfT7rpmk/5tgkgw64T8OL7eZmIjGsu9dMCWWZVyu76gzSQHUHqghqXZy4zg40K/5+g0wIX4HD30
tUTWr5a6YM1Tyf5BmdvjVaQw0TgtUSkvCSI2Mq/KEIvraioxh9JAh+cDs28gLj4T27OS7RV8rTqF
8NjWWa6McMKlzcDEUYhq1uYpcMsHKNbkjDGtAT/ELC+InQGjZotEKpD7qE9aYwbBWN/WmXwCRo3I
5OoVqBSKEdbySFv46HPWxh9xOCXzdBHlBxj7xtrNoWiWvJGEAF4Tk3rE/uYCSGwV4NDU98tekYmg
WsG2XNWLkxyAIAAGUTr/3c5E9XUzINhnI4Bauy2U2DIkwZIbs+nbB4HVRlPCpj394cmUalLZpJyg
oN/oPIozx/1O7uqCfBxWWWZLrYzU5oP4FnmgM7tepS0shtZyixz+vEK9XuUHOI1nkxReGZt2e5Cq
VEXxeWYpEt1DLASvIIvxvUMLunnoFb+1qpNMXloBLW/qgMGgL4oD1zqXO0mm2mGRDG0pLoFBgZIE
B1Qq0DVyIwL9YNOQjPeK3n//B/fHMtw0ldtTnSS0NuhMCN+H6FEWwxBeBZfEgQ8uHAyqhDqkjgwW
lV+5LU5VGE8i6aGpnFwEpitmJz1yVTAdj+4c3o3azpnuFJaUxjlacKQRaAUYVvC/K39WC6AQgyWY
8QHZLnEq+CW2rDKMk9RLDl66mBbHcbJIOL8ZBU+vjEimoNJJRGm6nqEaY7BtzPw0c8FcsYThgKFq
O0SsUUs7kHI+9i+dV9Z5e1PSMxYZOM9G8jAEzHwnNOQpnpRB2OsLPZTZPLedvKUgOV+nNGrpE273
nfRn+29wkscAXDaQjuOk2oMq8Dj6tVhyYMhXg8OH7f5h4xTNq1qsTbKUMMWd6W+8MUN8qF/Recte
u6pSGXhIidWH2DTdfmRNslhiWe+1bSex4k4JI8CJINGWpNceK+JBIoICmjbJnm/u+HXnot0sMt9i
nckrPHEHh+Wvdb1avRwGwOyEL261gsXrGAickRwq52LybrtSadf67UAaWkP4O379kivmD1GoAlcE
RjehYoxXab/DQTCm2jLo8clFkn//1Dyzzbby9qA8rxiYFXRyoxUOYkol6EJFZ4EEgEWouKc3yruO
pu+/b1yoZOA94bWKG1D4YvrgwciNm2JtCscLHLRbnOYsL7BCi34pF118YkbRYWbSDVJPvjilEmDa
VK4U6XaEQdmAhJs2FTaz0c84EHSyA8M2jGybWxXPebNJBTtyY3ButbKJCMb+UTx3SB/oxFzX65KN
2Lh/oAWiPEuPT5PIRdEAxfTunyiopIC+m9NoSuqIQ62uK2pq7PRuOYMmuVkHyFQfhD0hfHsKjmDM
bub5dU6zvSA0Tlr0gfrfJYFy7npe5wDyA+uGhquuNcy5eYi0i95FL4HfosKPB8P03Erv/w6fUG3Y
YYW1sEPlLj+lEEyd4CjrtnGQQ0+h2FpbhDbfGeaTa8kgeL0TlfGWmqDSoKCQ9/tlyLPGU6njLVXi
G2gALY8/ZAfzTmhjFUryd/1nHnTPkxwnseV4uvzcV5cEaMxEWIYk7p3I9xJ4WaDORJ8YXCWaF6BY
o5lq7Srad6ZYqQWdOlFtLTDRvg1pLHA7eX+/G+7OLtmATYWTKbDMPRDluoKT8n4hZGyjpRIITOjP
8UPLGAJ1MOGMed/GgWCAA/hu9t5SCQoX86ooO/GOhAaO/4/hBpBKhLmmGwin9DDX+f+lVq5tnBvi
Tackhocn3FwTh34RDN50vi1GdOu0/kP9kQApwkGSvEkufDAHGG37rfbQBeh/dkp4hhXAYu5ItjpC
1htKl/MyGOwrB8qI1agHhIWVacUvGa3acVVDaE/iaZg3e3naBNPPFr61tVR6CuMcK/a2HRxHwyny
2iFzm+p1l1q7+Rbgx6cOLdJes388maEyWxA7upTR/Xwgd9/VTib13734SWksQPwnHz5+jtQfX/Kl
zj9GOuBIQiJzbmdhXIWSs5TsjOn7EoW6v5YaY7MC25z6AxfzOi6pDh+hNZzk8iyOgPjs8gKb34ti
c85EkindLNIiURdnWhebT9ok57jBLVUHfT3NsF1564t0zOpWPbmy2e46M4GlFPNmvE7wYxFKAV1p
aebfyxSuO41XCWKfPuJDJVIzl3bFth97E006qiDg1Le+5lGefxnT16W/p6CYqlEewcMRDJ/wCrz9
17PEiTzypOzGqWnoKa4xlfzj/OLOmz6okpUxEZQve2aTAdAob/PRXgKDw0qpmhYYDaNon/S9OAhY
EwbYBbKJmVdniifXKUu1xDKHoG4o3DdxAhwJJu4AQQlVGA204d7ld9o3QDUPAiRoqZzfh/SKwWKi
J5xA2z/7OS2tStZ7FjIMY1q0nKzi6TK3d8LPWE6JP1lxiklHZhLXCEy5bOurqj9tAE/vTjFjuJMH
cwvp1XrwULIDCBWJpscWcI61Y26iog5MstRkc268dxlJDdzsdo50eL69SAIntmhVt+COxafhFIOb
N5thNDUhDQvvSJsQq+zHHO98H5yyu3GW8eJNZAbg63UX+WveYN7xgW3y+i4VW3uQ6wwxbNx6EuRp
wh9EessL2RhmMh97rLcEdl49fGKKPkR9XWyc/DGtKn9eERbu0NhawZTckdOUQhEmgwGOEY2P+n15
77lDBlmxIvSe3jjZpBueC8SqVDjPQnC9vh5fqJarBX4TDv1N0T7vgvuwti+0WuwVxdefu698BlHY
G5Q1JaOwbuU52PfAemnm16Mrs6phfCLFemAlGQcPNY9wcJopg+4uyOB3wjT/4J7ic46jYLlFGRdA
8O+scwRBGleLV/5QLTSZXrU/AJvBLKJ/I09AvIFzfLGLTDCFPSgVMNaasgpV3uizsw9fy+VYVSVl
8LtCxu7RF/HVno5QxIXtHbKLyIgSMvSsNQD+fkepfSAEvqaQCNgSV5bAaN9HMZ/pzMABl9o5Ch++
UPiz+8nGY123upHy11SGdJTPwAz/MYKrZvb+3DziJh7saBXDJIOtGqkWtgRI+Of8scqUUdlpFSSM
K+ol/QWj1qsvIOJs3TRAbhoGoiAjgtz661bfgbMIls7TpWd8/c4SgN1l/cePKtzk6KcRg+aMiz5k
HXRUEOkH3PKjIRs8JicezKewQ1/bNT5lBfdPd/lTLIECjHLLsVLAkfIXsi50WRKIItn1IBn9hBXE
cc5F+f4WIZUN0TpvFvW51YerxnThJu5MB4d8nlK/RufrQeZHE3kQFjRvXUcc0iywmpH66CwSkXEl
xnOceWM5RRu4GnCULU7jvd1BNvP6S31PtvFVFJqDG42wUh1ZoFWv7Hg5Zcfae9hxfOiLuaZmoNQb
zL0Rn2VdIaR3mtYDXr4RoQbEw/eSDNGxmJsL6bGrRcxf0E61gO6USfNlDGVtYb9f946QMAAsowtK
8SmRjoD7Ruhvkh7arytnsHTq+mpOKEzqpiJ+1ZGx1aVPVmTTgrch6t4n1imbGJer1Tmm+KCJdJMk
qpjwTrRIxm/n8Yw8QiYCVVNs3825frS9QiFoxeRaQ8CYUM1Zwz8FICtCusYJ3WaYlHFMHpi4cUap
uQruK3KwvyOWqnrOcndBG5gJIvR+eWmxpU6ZTPsHqBEX934xVf2hfx58p2DUswPemkgrLvkH2z1K
OCFJl/nxGqxsIOF5h9/LHiVbGoYLblsXe1zdrzFZ6i7QoybuhyxWQ+DptwCQYG6cAjU/ejlKmMjX
NFokuQQba3YMF/TBY41XnzZrcN4HXfTa2ApaiLOSLZ9gjbI0TQggEi7h0QUzAae0QhG+Vdzs4Sfi
2enRDvTo6ybrqhjPeMsmlPUP5zU6Be/fTbZaDwv/yymek12r33xdCNKyeZFGaJHxtXYhvWbMRJ3f
v/7MZs2Dc90HANJPgUJDHUT77loaeWhiVPe0Q4RSL1ftY8Z6OWA2ipgGzfB17yHXptrz8o3RdZPR
TKv0w6mUG36V24nh9jA3Ih5NJNDEQbEDNGvaUT7d2CiSIBJ3hZSIpRes4ydmGqOqY/4mF02hUjJp
Es0oAknlFXg2RrwHc3GjsHYru/7Tzet+TiLDPmfA3kOvlrGHfCNe53GPE/5UwiwMbGgFhYpZezvd
Y40ntUHaiENKEWitiRZ5VwHp0V+oMaKl46tuvBF2mUFAePelQc97n475up2xFo4Q0cba/Hjvrby3
dlE3q/0gefFsi6a4n00T7m0J4PWRMwlGul/v1bRvFBJCaKvJ4IuB95CAwIIP8AWQMA5SL5jkmIjF
2h7TswSS78oqWJqGrBJJgF0I/Jmk56ErZZKE24ajTGymekf8WdtZAZZdxAE50eIDdK9K5Sw9n0UO
CuhmzrvGtZ5zo5YCJ2ERknTn0bMKTqrpFZRJwRt9P0/DyOwVArDL4SHyryDmvUHi23xmjMN2YS4v
Y6CMDjIwf2Patm1yI7YGkTBxUKI2IwkQneUZW2hWqvdjnUlTwiBc4h/GaFIN34DCMxtwsR1zTLej
JtI+GOdZ36+oNx+NpC0y0YbYFgBZSWjeh+noTgck9pRVcvQczquSIfQLN3uEP/TPItJHP4Xm0JcG
fZtXUwlbpZtOg5VuOu2PangO8vhMA/BHelgtBrTc20VcGw+QD1gmKkxuANmM9b/kAf8fNn+SxT7d
Ch/NYNr+vWak4p+xgLgVgYwFdCvNdcGu+G870ocpQ3VRZ2K2a/POXZlS5BBhwlnK9DH8s8OjR1Du
st/iQ8yFZ1DcXkoTPkipUQXw0huZZAK0uZ0kJ8df5cR9CU1LlY4yTKN1MRGmqM/W+4df0ulnRbd+
BzyskRBEfOtbhUNNMfThNIIezchODadUi5B9ywYUR3VlR7mzpWXH2u5YvTVuFfKKsGTHbRqwjHfh
8KGJ7DFsHswu29eW4+KDNqbsDFptWxRFkTCdSH7BnDBQkLvpmAD6hQS1uZGNWfQlPpy4yEZtTNin
f9N1v8fh+gxnshwRMMzyUrqjL+s54XfkRMgWV8dELbStVQhZcUxmqDrqbk3ljC9f/C+Ro1IA3oZV
OX9pf1Wi97xw/hM2h9R2hVSQ+Y1AbtIy22qX9T/GZdEp0NF+JggvEgRd1jZbYWRZlZC0D/pmA6/W
inoRHqw+nS2VKJiQu2KVlw7i5LikRP3S7dup/vqCVxKPiADOSn1kdzxVlLqXuX9VZUnnLnLqMKwe
9cFeuq9HiajastE0cDFhgXAUF7RUcHkKSNyvMZOvPHC1LFOGRB46qsNzX5QccFiUeRW8BdDxoTLX
3sF3WGtTsUuXSQuudHZ12vqRFRf5+tlivdY4t8OCvW1PULN3V18ZUJJsNx1S3veD5/wqJdDgu5Ge
Qopgqtc1i7CePuCelv3E3TsXN+OVgQwWkFm3/s4lWakKGra9LHb+hs3vbiKjFlF0L65IL0WHt+1q
/xl1BBRwK7gQwXUaY3Bj+lx/uKCrkYVUFW7UIVm9LkMJrXlsDKrjT0OQcTKbIBkv5pNS/b4/pPF5
QfSb5Iw4vSUearzrQ63vftlQzuLkzKgXBgBf0ctS1g2aHZaBmGuT9tDt/N3M2iNh9DTwH7n6TnsZ
xjdQq1zUww1zDsVTNsWzHsvPV2TQ2hcspYJgJ2ErHRqZ0Rrl1n/YolHk+6v67K9p1dmvSsmO8pzA
kjdwvIcrh274iCIB7Tlq8PcgV5QQrafyVTWXr0rNmSOgCGn7nqyr+Ie+RWNoUei0grPFOX0IeI5E
aZ0g6PwW2tT/dL+URhwWT5iNBEGwG9LlGmCFJFujQ1dD/gj67AiV8sqLk+620fiVtKSD/gZpm+b0
QfW6T04+sn68I/sHCVIXQCyADhgTFaE5qDBvWweJb13NjWemdeFZ7fO3yFODf0kyKS5xiVH4YBH5
ortcMbYgjuiw0q52L1Eiz9IggDZ3BBqXkLoCje4mFoJDprA8L5FaG9mFV8bJa7xT2RX0GfR9V4YD
NckNiE9TKowTkyOdK5QZJSgR8TdA4JhujJlkZif9mIAu5XD65tHhOekQwJ1jDrTbycKj+JIBHNK0
yGOv4eoWsJ4OwqB7LpkLIuo29A0ELS5fLxP5b4oC9D6yIHGjA6qUTDKBu1RT733C/sVeA6ZxaaSF
PaJY2evhhz9xCrgLYJRALbiPCd7WgHg5WMPvmjc0yeIyggxNquyK3tck2mEZYNeq8mfsSO8fmdCB
yxmrVksUKntiXuYTReudnLsEhKG+dJRtVVeLL0PStpulsDIfADYwf49PAJ2PhWqSh5yKnI5gnUQ2
uN07LhHXPgIqW01LhFzKuf+cV8nLjte4OmuGi9Jk5uErCw4jej4Xyib59Q1HY8XZ54zBbcT+LfFg
kfbHngDAVZJIU9fNS3Jp3RTexLFoWwcqANhqIZzylwSaB4pTN4A05wQ3xBkhYhAEVK++3XSW5tBm
SOcyKMWdUCUCx+jjWcYVkZOrcxzxOyMC0HPNaNwsR2g/9LWEHASuCT+35CtPaztYDAKL8g3kdBAN
NymKlzZuRNrfGy66f/O48hsIfuPor2n46+hXm7YKbDmFi/kr19v4Ff/w0/gNqwQMRkFk3AKx7diN
JgpoVrG8/8r3NAC3v7WMl+eucVWwf5CE/zSReKJlm16RLXq/TyTbbveotF2DpB8dSB5f3o1jYUi1
cVIIZqQLuQFVaFaICqz9QKqFv1lUek/euYdrs1CKKPP3Q31j2CMMx9/VYR6dSfAyvPJGwxfszOlR
JhoEAlmDfpgnQYNU6O5OiLwZl89MqDu2tT6eXRrZFfSLnWA35ytpmVQC689ZCKVsM5RgFyjUQeQ5
PnRj5UdNaSp6ID2u1NOoMr+WEjvC1jVCipiPnXQWc7OmrS7806jbMnbw+AKgXfEXpIoRFBHoYAlW
h5aHWiasMT0atXNbS27xB9Yzk2roBTuCGDLiYxiXxkkMCz/9QH9/FFDE3QcqIn1+/fmRJ6iJqpmD
ZDLsQ9smb20KrJX3oiIkrZDJfPWwuq3k7WI0rg2gGcLBX0Xe5vcWZxl7qUZcongYHQX30bV+NHmW
9Du3VJayxMKeYSofjzAzMTpnjkkirZSE2BueMVlRoZnkvdkZhb0XLPHiXe606yLDYi7aSWbz43lW
3G9IeWtwImE9PNQky5kMs3BlqfY3l0ICFL5u9yWDjQzLZ9ikH9v3K0vkiNJCogg7RNLXIgqBWgw1
NtWOglmx8hEM3gLLy1U8NcfNJCHNNPPPa3Vk3tAejnfsRsEHA3zGKu4j1AOI1e6M5Ovcn2aFDh2p
2cq2aE1JA5LRz6XF2NKvCRs7rI8VewsVIRH6bCrNQWbw/3KtfpjbpfwjZqFkJDlZLN54q8nwDwxw
ZmNqaj6xhhjiz/ozIsTd4BeHJUiBgyzAvB6u5K/DdDbbafmvOklw9KDUyvdv8AWl4cAyijOppKrE
onVseuQJd5ct7rHjPu/ZeyWWzYUQZpUUV7y2r17mpFfGXifwIKqjl+NlqTjXM23zXbMYcqAXn9T9
tIiBeW5be8BkskMq8rxInPKEQXrg0SkZAovRLHYoEoPSdrVUhBlavWpbHrkcoAB6smJevx+Avmu6
rZPCn3hZT5UX5PLWkmtfLwKoqu9A0mbwLouiE7IJAp0xRW+9WZGW8dD426oG3P6fFs3+nqO3NU8R
56J0mWqewcOp1OqftD/3iQ5miFvJrrGUOZ45d2JOBKEeTvk4XHxso0Hju4THwOqPaC+7mnb4VKBd
oLnmFzOjvcsEuTyxCjd6/T5TfeBke7eyBpYo9XqOmV6atC/oIE1KVPCP5tZTDFzzWYnO+KObfAzu
Bqx7jGCc7noKGU1kG+aDQ6njSwmiUuf+brD4RVC5aMx5iIIarAwOs/fZ5GrVAp5RQW09FbbWzYJm
CUpD4zUWMdkWxtu2YyAXG5bcFXN1jAS+02wLblcydh1xojD1/iN6uzVvh5mZrA4HkCoPKL0w5QvD
B1Ws8fMzttEUI4t7YYosdc6W/0X3hJkw2QkzSQB+S9MCpHehDslJM03QpGY5JNKiXICY2G/LbfLl
Num9CObu+CUklOcw7lyFOoBYKEkZUa0pvTk3t5M1t9rweJkc0GSbNlBO/CNe5oEn38ik+01tcXJG
6rJsgI6NBv+yCv56EmfCiww2uyIsTR74vCLIaPsse3cdcnpybFlX6uMCEt0lRqDO0lrrV0CdDnJc
SbtnNjc1h18vi920IpjvfvtyKLww6EMUBwJOhhOeuXeczA+45tMXh7QHec+c+05EUVIc454x3rly
zXEE7MwMvkpDdZ6xYpXohlzIcUoidK13lBlhxkjSSnj1V+wXDzTkLgBZjBzlx5bZ4dlPrN0c5+u6
8FGLOpDiv2ypyqkPU87zstOMaX0GhffIzXD5zfCdYL5F+kr/q9+jcdw6dfnZz4clF7ulta+EZH+A
vW7Z0ia9q67H2YhOX2sTGDIoFDtiC4DjsIsc5IUuFSFnbH0JbQisYTgb0D1yYVfcnoiRsb+oPQEk
lDxBK9u9yz47p04Ca3O74zPW6Hf2UqRKWBj1V5CpoU2zocMJ3q1TlZytRa8vgQnR7UdCauMke5qG
1PkJ7+3BGkq8UV0BpwLn9tGgqiD659o6eMNa0mRLbraY4AH+siIjaGC25bp9PXgMdnGrPrncsEsh
ZU3kKk5iwkN8jozVpl30gADe/MdYaBFCj4CjAkmM3dg6HE7VUngXI5zuDE8oTTHddQHitr5mEiNm
Q+hUnx8xN6sed0GYKQIH79NyUAGde4S/snWO6PQd6U054Vw8fhOqI3TWL8Xi1lTuklMthkz+9y5R
lg9DDWZ/Rb81jV1dbIFpjqO4wMyZ0bLP0jVwMgO39FgAJRZ6Sf1ssY1P7xtSr/c5cimQfrVsmxZ+
k8FJLlU3CRm+RLS+rQl0JXytjzRMdu2aw3fCIc/5fqp1YRyaKmzyAgB07jw22fnVAp+TlWiI/d8c
KaN0s3jaKKNIZUaXL21q5OQS4Im9H00qelTqutmKHbZe7yMn59bBZ+2dN+yVLICb0eiLCLxK5bjx
NiGLKUPIfj0hWCnnuF9CI2O9bsITL30YMOFt0Qd/QRL5XjKQKpAwz53+20Kv0FA4lSxJmMAAOf0p
96ekGffsGyX7RWWCY1cxsetoGXYExaw8LVjYWtNqHbXHXTeAV5pEwhhNNRjHK8DcpqcfGutW5oKq
zKdi+KrGeoX5/ZKMLoCf3WLpX6I51Yd501qiSC1MJzpFOzNUpC/IMvG/INnumgJ1p54tkvMnsmfR
AlyZNYdU6gYo3vXtROj9SWGSG1/NyBeVCEHCyaw44s2DJUZeX9zojgP4dGsXdeD2elJrcj98LRtW
oh87azJI0FLCO7Ld3XAFwZjYNeeAN+1tsyaUDqMKwI/0MDMORXJwU4GZlRH4UowUZeM4VWxG1+mp
BcrjE5HgnoapAznJH66bLK8z3Y7nHU1g94iAQWMAHoMg8reBzs+VK2g3MJtzZBl0p2gqKX5sp69L
Pjim8P2dzPjrTYG2DPcvFobCxZ/mGNiZV7WRLgOobbV/zxi045jk5udP68KluRbsUJaST/c1wfvk
qtyKokjKWSSRFBvfS7Ds2+tD9EAl7Ssv6vdBZbJ7W9dz1VnTXPNLaLWJmrsjhjS22f/PQoBSiz3X
cObUK0DmTNftLTRy8nGENR9i6CsL6d12FLr4Byx/JOx4W1E88oW3qOl+ZaO9VwE22LtGj2gwSp5Q
vBiTiF5vE/7h8SeCFlp2Lktv4IE/Vu5TYutdtBKXiYx2KLmnBKoNiYc0ze0An6SCQQHlTsECBjSv
7gHG9n39xzSbqmk2JnA3JUi0WXa8/B156JuD1SAgpDZD43UQwD9QvesGFo8omwZpyrgxFwSamCrh
93l2NGSJFKz33jk7lpCwBl886fzcpyrtPTAtDA8wPUTCHLfS7dT0NFZ+VIilqvqt5JPRR8q5S0fz
C78hD8eOKWo0uELTO0gxlddb5i4swShXfphCXzYDulbcDePlp2p1gRjZUWa0U+xdINGhFi8KbtAZ
5gcE+0Pv8cHIpNoZRl13Bl2AxV13jxKf4ClYEOId14x37QdcVO8Kglr5tyPlafOPZN5PiXhasTQ3
TbAyn6yHlH/9vWHO4i6TQB17366IisPlXsHlD3S3u7Vav9rZxyGhFPCHS621nFcx0E1L+npxNO7Y
1LF32JZf1Rk8mZPEzZ7kZeYzQ+qEUxYcim6H9VCPjaAcMY7aoec/+K+rp5Yx14BHQcGDUFFEGsmf
y7dp52Ptt93qrWyRIbLdbuFyAcN4dZHqd3BtHndh2QNgu0oOIqpIC20qt86iUrMSxcgMzjWtBGG2
J93Tr2hhQvrE2Z3VZE58ULZIhJuUx6hZprWOt8QMYkpxagcAx3bAtjrOfbxX9LvdIRaJcuAI57dJ
xJAW2LBZ7vwE4I8P0ToC6g5ZIPvMnHjuqjb1yAYvWb9abQ6NmOkNa7S5H26G+MxnGZArGKTr33EZ
05U/kE5B5uZAgH9P590Ab8Hc1GLYUv75yHXZTyDAoQozqP9onKLm6jOYRABKEtR9fGH+7DKLcO0q
Cf66p2JS07sl1os4D8KNurMpd1MXNmFXBMPhkFMb+wANsuIodpxLSM7rr10V6YlUKf5v7+kQebOu
EoIh/Mx+4aUPa+OmxnQD3f6M2ISkKzOQwwjq2D+RJji9SsQD/ygU3tYSchxMr20+XXGGuJmQ5UmR
IIQbrS87TijDKlzSqoj4wZmXQVV3xygfFIDhZWhbHzkRZ4rlcq8RgP97mV/agWH2JOhQojHHtYWY
mfzDBeYeTzj3dZ4Qkz0fabfTG7k9hbAzKpgIGLV18j+ZzhHO5LRyo2tYENXRXOcyWBKvLZLvHDWV
e/kQYC1d+kSAAP9G6W4k97LyvrqHZrbLnYFZSkNIdILo+5mHZP4lxHLo07FghjrSYFo7m9letynb
T2TmZDqvCLUffHYSTP6yX6UG/FdhAHMi84/0HKyo0slHgm/icRI1DCIV3/C720cK+pEKMD4F1XWq
2pgib0D8x2kaamZWnKQa9qKd61KAQjQAA/ZQIkiw3M5kCdh0g57t5wrAlOEg6tNR1j877fd+mPrE
KYiIF+aD65j66roqygmLQ10+jaotNQWy2jaRuutUFQct0O7BkpKoaCPWTeJA+RAQ0sQgURz+GTgo
uG8o4Clol+eVG7jGkRyadcr4O15iaPmSX0vjAONtR9mPgVVbUodkKfY3RLbA/m7cQ1PvQ5osbJfO
vmYtbLOmjXDobMsgy2qNGx5dPWHYqcFvdLAnp0YRWdggrEiw6RUjEHfno4t8sDQFgyfa+U9qBcYO
Bg8hsoh7CYaNkAzNEXZHnz+rvUIFt5aWiVJKFt8q5YYUdEr+ZbLwSSxOq+fBmMB3+ji+9l+TUz0p
QBSYNl5yW8pEN29yVOGgG0hOLZtH83AxN1cK6SMtKx9Z8V0yU0Uan7RfONhWFi5XMLRhTpp2qjsz
FI01DdLKGltU2DxbDUBD71oNgZR1ngyX5d5m6ExX5HaMgCkK1vF01eC/SpsdanLQOzOB5u8SNMyv
pSulwykhcdvyeQXU2sBBGozCdPBeKAvJBn7HFMQgzzdRLRriM5J8EufS4KBxU3VGUrfHw9iXVyeE
NChnZN8hnL4bQtRheMPmd6777InYlLlHTwtm+jBRcCO4jemSFIZLOWo/XSQJfXMSnFmI9ZQj0ZP0
qhGDv1C8Rnjm21dogYzTOVFzebTBgU4bLpogd2EKst0R0N6TfvArOGlLeRSgYOG3t0CGTzwEJfnv
/3rjziU9vN6epRblwEe7ZOkvDFI975QXb7lA2J05drInmP2MR42MFPr1JJPNTLA74cjzTHz8OR0X
3CUj/NzfzpOGkJq2hWeugFezN7F2LQm++c0mXJa4m1+gB/40V1r8X9ErhyxmT4Kj5jHhtjn80u/7
i1fMWzPg/k0TVYqNEggPG2OwLXy5nSoJeK9s+6muKuB01wsLjUvfgdsiKRGBLbyRvSS5Na/TY0ll
zKTvAw3QpIBOBtkhozAqTCxuDGuDelWlIN26K6aQHxNGvL6qZIfRBNTTJU+ZmWhnKqIsDCGjMy0L
eiN1i+hgZc42RU2p/wa6H2nR1xRelKtjiCOI9SKfxZjTM8KLB+lI4C8l0mWa8WemTEs6Qb5KYCSc
kdaZoWwwnI5/adfoQcXc4e8xSgFA1FSKiC9Kl7g7OH7b4gHGNpvBa7H5TlG2oitI8zxZsW+FsooV
Ee2gzATka3vvkqn37A8iMVmJpnJ8RrQbjTvHT9UKYlu1dwrbhmwOLTjaR0RFVUqL/0uQHTowuvt7
ScDNvQa1JkJv9WfIi9lapS4gq0jG+H/iJrvY4qi0OUUuxffCv6Vz/1c5yO9nDgqsBLP6hrYMj6F1
Hw72+a46nCt9lAcBmGZATR+x1HPk+VKBuKOvO15f4ILI0nwinBK8zr63Lx0yy4sY3NADAgfuAus7
5Qzj3Qb03oB86z0MW211xxP6zoMmr85+YTUnDPyqjc0NWlyylDZtlQHw9njDroazTiWHglxUTdU+
l8N2AtDl3oDtPtLWHjskQa+yIxMYQq7wO70x2TlXOBsSsvYKlzG+sh4AxFVvFavPG51dKre8ML32
37AHvtrfwkl4lyOvqrO93WetcptnqwNTyAFKdTEcPRkqsX/O2iEnxQ3wcoDHs+ziwXeSLVv01vt9
Yxsgp6mEmD71HKt+7Auf/x9EnANQavRlxmNmZohL8y07IDCuaeTfpPAehkBIcrZK6xH8Ets6qYOu
GVq3fz7x8Y06nYiZQ3JPlXS1rtyeY8MtcGJKWfHJij+8B+ycKY13056yWpMv1f3JQjivpduCaJxU
Mjs7s3vOpH7QsOjUXpQhNnDhPpbM/kFHcp8Vg/e4HAVdJa6+kDXHtMkLGOd+wml9+ysxjhz2HIyb
y+V++0NfUF+GbnJespimo0FYizbd4SeRqO7obpemQkK9MZfVfU+S8Hx2KJTQ7JB6q2osSsEOpUyx
/9uZAO6D2uioiK0y9LwddAwaKIjI3qD/4BeV8TXyPraVrH6Ju5D8fIdpmJWb9tL3yhKLWljSUWry
XR51Tf/LkvoIfMdHqjFfx0gVdIILGLOSRwvu4A1nRwi08ZIlRE6yfIiLaI1ViXh63kas8EbOob0H
H153BwSXj3MwKfrP4D9i+ozg0ln7keMScqbZWhLqA58Blp/i1xO5WLL1Qimdo8LCpfydmeKTi9wt
/RKtHPLgKJxYTduxh2iaiptdUiRyUym4js5sKIjX8D0LaNwmc9EdwZW+g6raKWbIjvW9tQwKKuyM
EJC3mztmPtn2OEbQTrO32e0PBKxb4qjxjxWBU7RRtmN4ecSAInYchJOK9GfXtuqWk5JHUbL8qknF
VIhrJYO83Pqiu5fzBXQpTMqrNvIsqKSlwVz7fsae9/W28MPRuSerJfMj8kn72QPeuiMESnfRj5hd
e9QyLA2eotSQV8HdgDq5iD+gYD2gctaus2UWWZyKOZNgW4oeOfENtcVq3SzD7Snz2V9RSp64xfEu
U+SyEgyIyKAvm1utWcSDyXyBI5zKBZ2TLfHTE+xGz2UmJfLJXUTKHdwr99/uuKjynFmj/FRaBWsu
V3m3VQIZsxnu+BNNYuwgkYwh9v4qYBRRWyS2NZV7gjI8+gmbfNr+SweQBH8RoPO6BsFemENQbovg
ZMzIwZ4rJj1CpJQ96hD1RrMe8rJI0fz6AunNuH48q0W4vcNESBkSpM2DsB3+iHNJiOiiVIf8d2bS
iGut8rNkD57q30KC1dEHHwNzg+6pkJITlBZbn8XkAPmR+x1JzRt3MIVOFHnmcmwbNRXtoZHBgT2e
R19N8vITd/FSU6CQRVryaCuBfaNAgTukPtMC193JkA2xJpPd5yoHVJQWXmqjOSvWQg3z1dxpfLgT
m5OOjSTKB3iXRs5j62ADxTqIL4jAdJlwe8bFWYUJm49jFzg6hnsmwIiiiF0sZe3WUyu4rN1XF3kx
QLDnUDdRWgbaaJmmiICxbvijmedZeMgCSMe+UdoY3W0zdn4vb6r2Q3hIG0IBz8Z+LkWfTHaOnbpZ
QTHmu3PvdlGliWbMdp7+nliLErwr3TbkP+nrxbwqliRzfD/Af+WzouPIagmW4Vm9jEhJ+xs1CLgS
pJErC0S/zWQI6j57Au7S9iopvJPpj8CMrYc0Gr8kGyVZTgFIyF9gnJWEdi/gO8HDEa2vL20XvORQ
ANR0UoF0IMHNSS1Ymi1T4/4Aq98vUMAEZEe0jdXLbgcOng/no+icJptm86gVDOZJSjrURunSohLH
YqmMC+pl9eP4ADGghDRv4rkn4TbYj7o7wF2/nPJ/3l6v2IUpfKjhMobOsHeDO57dmG3eGnuyzI1j
U6T9iPM4Ndl90sOlMoRG/IAuz0LDDtSHURvaMRhk5/6EV0UIZOkHxzjUpGBXnVBGNqvJSBfSgqq2
Sccy+IIy0jcCb1HJ1uNL2CNGMdomo18qKewtRofzxp6fyMZHtrniyps6FKaZDdSVlZonGZ/scCua
IRinPX0aGpO/hZMqS0C4Myq0YYOoTB6trU/52mWgVLf2z9Nb0qhcfQTSGGmTQyqdd+0iR+lhNlPN
MxqqeGywSZbgX4haVO4ojc//OdzrUm5HytORpBwh+xVlvbkresbHQTtucCF1IS4FCWo2mg0zipkU
Y5uHIs2V9tZdT2IC+Xp4WysK34YKs474On3+gSgvbR3IxZc4+hES+nlyRdkYYdNBQPqDWYtPerK0
YuqEab0Lu+Ipd/+8ID3Ngvm/r5SNu5hJrMlkSDqcE4l/WHEly8Oretpk86BKghHA/D0/gjT3Bhg1
2iHw4sfOe4Gqf+fgD6BRpUrs/U1Ebzup3dD6c/lliNiGYtJazbYntomDBTuVrNCofOi6sw5dAdNG
l5ZHM96UcaPVx2tt+xkuq3CbADB14Chy4dkSewK1IwkzMSO3ZyT1MfN/Emy52nNy39qkNAZh1Iix
lxVZ1rDd6RlYvLlWxBnYdcw5Lf8nvtZRD+dz6DpIzxclaKF+7w8UDDIiJVl4p04jkwZTl/Ajjq2w
5JxwD8LFuyzKM+Mr22jBiROMv/DaQHpS8Dqynt6unUgy75XThOl6RGIYJS+1idRJlXFkFrYK2Pws
zdG4Li0f0hAQZnbZQX+ZGw/yoIoL6twmE4G58rIWbJhaQSPmjklYoR4fPMMGfJpH9lj+MDCmVEjw
BiTz2bY1rfMxFRNGsTP29/NPF6P+QXewXXiAM4QTYVj8ZKDWYBUZ0hhVop0tpsaVrF9lK+rUrNk0
E5Y7vaSHLAZG/Shrs7IKM3AQlK84IeS37TibwvZTdZb9ZPX99QrRPLGCFPMh7UsPSnAcDdw7Tue6
YzDcY9rTEhbWTSbFtgPrMQqeTfhpJnb4MbMlXYbxtItag1z5FEhNUbSihqYWlwR1XE89D3fvBzWF
WkH18djxUR0fWZBE/NN9PuI7DETBE6aqQAf1Zle1lWAEMYRilCTS/K93u2yT03pNKh7sJCPYvJr5
Vh+x11I3IhgyVWKiN9kNLVXRQaMZdUGvKxMmSvpZkk2RTgsqt3sR1iiL6q8Mg1yu5hTYBObPpBob
bN77i3HGJx2PjcKtNx2iMHYMPUAeLfx/LqjnLABVu/5c6SloJEsCTWKzZKOYPMApZlMlVP7snyoc
ED60ffI4wjpVerBuj07gKt73+TW0oGO+tnzfQVWM1drEbm9HH7JaRQHhUF6W7Z5LqUpypoYY0OLL
0Mq+/2wGL+2U4Xr/Z+WzjAILdapMpoNbwI1Upe8SzgHKn8WWJh3KHaD5dSlCytRw6q3MLjkgB/wq
rx1ih59WxdmqfWKLGqP3ZIzNdDCY1218FFnBIqGkqeV0QsKVBsqNn/qiRvs7PDhlxRvYL9athPU5
RehX5lu9BLTeYzO3PYy2tmBwE/wK/Tz2mlmzUiOTcvxoDbG65Vo+rG0cH3UCHKvteZSIjJ+tiKyl
xsH39dhTrCXPFWJwTaT8lItITcZ+i/uDjaD/6FIqigBgP/cljPZTkx82sAsnrc5cdPg13WpiDh0O
YNIaCeHQIS5IOhZQoqse6EQLBRzyqd/6QaEO4GC1j+Z/4KBEaT04fxy0tgkxfKbwA7Zawtt3/foW
+h7xuD0vUZXyf5vWHg/ZyexfgVkwUVoLRF7f1hw/MWp1o8skfpl9bWjBVxpkDcKNxD9FQPbqGwGl
wScs37c+8oJfIuGC7pnRz/0p3a/wcBiPWA3t3t2lQaSJMojnBRAlOGtkS1Z80UgylECZ5EAtPYd2
a2oa/QFIYTeACAXNQ7MF6wgaozIc/pCi5wa5ZAA+hiclrNVn1ahHvi5sMHOFBNFJ8vNhdGmWJtZn
fGkTwpMoP1jEmZvhKN40jFMqWz0rxaKOnq7ecDWEHXCrT3YPh3+DTcryVpKSmGZVU35Koh9XBRGV
nZq3edUUF4Rtyi204DTU5Egkyk6q1QK2Jiwol+Rpe0v/06RYcnXgY2aGk/o//530qQa5Y1D4VMLx
wDxBDs4dZOV3EDbtA2cCxFXO2kajwb2OTDf5wBr4boPMmmIs1cVk0RGFy8cBmAdfYg8dsb1QLvoD
Nid+Xa3HRiEx/YuqfiE0jb2DXGz/4HISCwq2xqABFZGx44voV88DxpGos0wqb1IEeAPo704bloSI
5F8q+8ejfsAvP52mQaMDS7koCx63LY5isb9bLHcdOr8L8AiotD5pVK/TiF6F2fD0TGIAfwgZQZXD
Z364UfkKS7BIKwffpfnoHVMGAkhP3SJI4LkwVfeFHLlyQWlxGhLSSfego82XFer5QdNhlqHWDMX8
tHK/1Vj2Lew7SgX7JVlkbeQgK4OGdGsQvdszOdA3U9jVi4mJZZRD98mQxH5PS1VY3cJf2gDBn3ZT
pc4rwFzHEHNtF/z51PtQ11ysZJoJxe5VOJVtcvm6jK9YKHdrqXp83LMpVhxwBpyAHFRFyF3VGCcZ
Vp20HHWgwAh1m3u0uEH9Y++lGAxYUdb6WHSe7qj7lhwSd8f03LXJGNi0/2jxNkM5Wn8LBjZ8XfIL
vrTZzcYVjJjC7nTLdwkXg9QwGXRJ5CUVNCZx9soHPDHfr71QajwwBAiaJ9J9ZlqbyrPr0o9ve+KE
4PjknUTIq5LluMAGOWi4Zs9qT8zpZFYZpjdSjbn0ZonffxjQfRd5YhKelnkY2oaWBS/tR2h4PuAo
zfqQmHMZU00yV5qBwr4RHPYZ0vjLtn30PK71zmdVnEuo5W4cQAhjwgJK5cHASgCz+e5wPt/ue+9u
Obil0f/9aHrhfLWdU6reUo7DPPJRM+xsETJ+/adEAeN/8nBqQ6pyA8/Zz6I79InhWDtv039oDVzO
kjZDaPe1B9x9+cz7+ihsjwWbYd55rF40B/sSEJT252qBih/rmCllWvtBx9hvkxbyIE80F+evu4eU
xFFl/s3qGy0WVeiZCEVsHBi83D0/GTScvS4bFNeA9wCgNc0/NWkmhBjnn/7PSbpTMV9DeSjQkSOe
zJQey31Xkxa/xyV/jOTQNjUuUyDd4u7yvnOghGTW8HN7PQvP145ZHslWE3xMCwHuYfrl22dRL/Lz
cLgZwIKVFWZune2JoSDj6fI4yauKB5a1/OCC1nOlN3OHZdjy+5XIjOTQxwxsvcdAr8yUEBgL0sMd
L0YNBKRO4tYJOJw/eCBeNzkBa+zKZ3xEq5Ex1I4MqwBD0K2QaO7Kv31L94F44hOiUsdiZfCvLx2m
HZnsvgzPPciz2aq0Tcq0K8S0GFs3+jpnaPeIa6jdjruDpf4wMMEkRYL6EJDSkObvP4obbzJSy7s2
/Xvz/ltkCguBV8QRMRmzzwMUD3eKTfbzs+M03kwgoWAB9VQ98oUVdgRFOp6INSwYK6AkUaqpdCQS
0YGloyoU9kooMrs9lDc7lROodIuciAlxSNCyq/XuAmbSXAaEXnJ0qaMbgFctjqXzpaccWeiSBK+g
Oonz31elhzRrm2Vq+nI3BMAPk+kBlYPPdQQA/JOT7yYQHDVt5yae7brH+3Vl9uWPc08hJaHbMRCc
pnHSQ3MU84iwEzh07XMmikCnpkAHfldsQuuWEiKOSbsVWupqyjEVxQKtH7wXayynCC/CIfWi3Z8B
WQtJ3e/cUOOpPD6URSxhCBmEI8SCpVOYj7gZw/jLO23n7FLQ1n+6VWiAsRgwxceao+Ah2X9H8wUG
dYw6ssFuZS7kIJYxgbDFIwQTc/7i/ov3nW6U7MmiLqQIxNN5shYXKLQnCM82ThgCcVDINb6NOpjR
aXQ23DbaJNFXmczBdsD6TkoTrLGOeDwxvM14xqZ9cA0r/N7pRJkQ1Chwds5HSg6t0REChh3oB1lH
cChc9hH06pDsjdfcHVbN/ncOiGIurx6SHfy1d3RhaMkILVHeUgY7QL99Ux4WQqUC+iz5aLwvwq4b
OGpnU8AJMeiKWKDKuao46qxEiozFxzOelPRzFsN53CnyDW7d0rm//p8lIrAZ1eqzXsJ1UHEhM2yc
E8BmcHK8AU8UZNY+nurDU/vxUMViea2epUOePtKsQh9q/n7I3srQWU0LYIxPl/lft1WJ6vq1Lsv/
O4sqOgTDrZMouyPknqTpZklO6dDGagyBfW4lecOEVCN6jIREoHvGkK6XV/yNahegJatYnaCNGp0O
4uP8J1YZLa5+1q1V8Z/pWtT9X3VGEkKSdWJVPFq127jOnVc0rv5u9q1zKF1zvAiyoAjAsta5H/0z
Qas2Xws26W1PP7EPiGtqnEcsOQE9qpTRCi8CbLw3c2zb3+dvc/nxeef5RM7XankEWIAJBmFv5GaN
p2RHibeGkCGODiHHMh0AM2ASZoICy5KByhdCBvI2+MhbNfqDder7D48tC7WjTLNYlLCiLU0BMNv4
7AR0r1aAuntp7zy+8QdZJYoNExcKKYeJmw8Rzdxy8uW3GQUQ/NtmbwR4rsjUu9zceDFJTz0Nbt6+
At5B3l+n7j8zc4Xc0PO0ZbAlZqNvk3ac0zkHrwTOgxywjzTpy0erjJZsQLjFArGXXWxS+A9o29DQ
hIBpKfHACthnWUj+zXt8DUrcp+Tt9t2KKLjrMwac/89FlLjqHbgiG75DEKj82SzPNaujhxXNOS6s
MWkj3WJsMnhVuUaE2m6eSTf02D+kaRR+630sNWZwfFDL385fxyLiDYnbEoWE7Pjj90nfmcJkj9yQ
fIWhjmixTo+fUYDqGuWlu9WYlTdzJvto50yTrM58c1LvYO863deJ14YFR/8fv6HzefeyEgoMmKQU
WetBlq9PUTYFJHS6qN+3XzVxpb1y9KFUtp5w6aBvr4d53PY5MUPUY1pg2cdLNbJ/lnFOC2avb8jB
BMRtKOR5+SzuarpZK29AD14WXYp9qu4iOoZC5hXhN60ENUitfTHSzQvgLWuZb7usOvxWD1BJMF34
JAP+FUqPfBaCbVUp0c+atWXTdEZST+KKKamQMdwW5fJj0YYqd7dsBoP4EtnTjMsMZ4SAWdzy8DJs
4oc+jhPx+9LzVryoqCxsL45r7nkWoG0jlvye1Io17pL3H1oNET2smEgu8cRsZDkVPLudxyzhfk1r
Rt7A3TVjBLZbMS+5taii20+j+wT7BTigpTqPp71+psNL2FN7g1R9I/rGFT+6p4yLEfDzNYXigqcX
ZYR4al2SBYn6cA3OnCIg4wylQ14L6NdGgQFPMoqU02T7aTlqnx06P7kLlX13pILTIzruHCEDiE1j
+UbeGnVxcCdK262JgoM3gweXLZiUiFkhUieKpMUY+DL/rgfVFgAekzrY8VrYselu5PEtCokWzOr3
a2qfEZmZS4BCsSeCZukZobnufch3BFS+E6RZepKSm6UTsMPtDzD5azVMNTobroURyRI0FnpXp0F9
Pdj/zg1Ow2vuK2NtmAalmE3QfgUFj1P2M0TAbWZr8WcotJUzEwFQxEIeYPJ240ep4ad1b0B1nn0C
Op+Zem+9AAKvPvNwAFkAOYrvd/oBhACXeXXNm+ks0bZFLXFaJrHd9I/IibejEOZKJVetTTlTsDdJ
2VE0Y/8psZ5mHqVbUaITn+uDLO/BBFtnulL76tu3qGF37csSmbpW3L/qS9LkQZ+wo87DNH7oTuv9
1mS1FtuT0xv7vZHgziliKA0dSnBZNeTs9oTRwIQi+oKU6gksoxjkXq67tr75/KiDDCAfXUhL3whf
kkJ4O3LfBleAetI37AC+gJntu0veoy9Qm43R/CfN8mJfbYqlkP3Pk0QYQEt6ZwZHFePYVHKBqI8c
xMQ575HaOEmE/YTeEH3P68nwrOpUUBjwo9uUR3ct7mYqgzig21aoNwG7cZAvueDig1CnYeu1nYXo
jZR0RgIt27T2pUID6x7rpITxZ3O7BXyFylcMcw4nHPB0WHOF/RLOgbEehyFw4MKycVVEe4FR0xYp
QkxBi05nlC+KmFZQR/r6xhqijJ8a1wbMRL9o3t/UEsABVjriFIEu239D81Wx310/WDTGgwB4mgQK
m0Br+RbJP7pXbP33U2p6adTaEcwys5rBmRgCq7nPhnqZUpJpMfDwN/6kcCdyFjDxkhnlSBgIiFgI
3sFVN7V8mHBYDTfSsBQ7LU/ArhdB9WR7lycWVwltnRqNphyjIu7cvGaM18YcnHDG6wxBGNwMrxqq
cdtor23b19IdP4NpdrYxZ+dHVZHn8VgMU+o0qW99hXoSFDrlcvzvCF0QOtwDN756D5310JHkXw2o
4nwWrCBwZQg8h4l3DHTtOzyuMJtvkWNO48m/ImS070Bg3fYBfrgrIEZLkLXW95hnLuQDnsuj8tax
9f6f9mw8pEbTzVx/1bTbu6ns/nC70y9VVXymfcuyZ/RaPTYvIUqWQhxtoQAlcVmCHoZLfDthTGKG
9iik3z2rQElaov/cTjTBHVdkDdzt9Up8tnJ8DvM9kkULVo35qWyWUG2b47pLk8uzdd/8FFeOXsfJ
9yRDBpU7l2qLY3nraP+e8wR+rL0djZMC2uZYgRJ21FOK0uQewXiIer5WydCeP+Koo4zscUo+1sgQ
zRIXD02wxBsAx+ZAPlDx86Lsxd77IRsJ0XmelDERHY7kTr+p0iEUZ6MdXYU6pNIA/6zZ+l4I3IAd
QOIgdVnmnSU9g6w5H4rLN4vStLsSNUKGyMJz2Y5DLAlnOpwtA2rg32RXDoeMPZ4u8HY1Ta+JH9f2
OTmBNQgEySY/UevV/HG7vXs4mTmOoK0D4YMXVIoxXbh5MyJIxECG/krxVKsJDWtp5y6DdVjlRfS2
cHcIfoToElEn6HZ1S9bCo0pWDWs+w7nBNpgvXK+msxD5pftw+w10HwbbKClSmWKb5b+1600Zq/3c
VZmyZ6W0yhrFu3X2zzKlg8E4c7j1ZpGHYyoog0ru8cUMKQj7C6+JeOMYyHhZtdLfnTXbNHVSRiDz
YCEfSHFSaAQlCMmJiUAx/PTOd6ryn3oV2fhAUT7NkbXW7o5iVP5XOyAqjEom20PX3tqbzd5MgqNW
d2XngtdwYyBTci3buSSG+Lk1NZaSB4WSIPkbpKdhGboY1qG7ya4xGSenDOo86OyiqsVG0iCCnIUW
Y46UsAZrBhyX8o3mcPkD17S8QDERBOUfkfGxACW88t+6E84tHnP+P07lIJqHg0XHwj79XcdBtY5v
sIh/flf/iI7uhG6rQZzjUcmjYtg2xlyWRsjreME5cxWZ1plGgyKrYP2vf4Ag5sEmeTv0arL/feZ8
nfwrTBC23KafCaFb6dpiEWDhGyae4/hryEsahoir5WYBvifHb/s66YRhu7jqoXKM/s+cEyBkQqio
9TlOI/Fhpm27VL3lUtrCvsi7m59BTb0De4kzZ0oLumM1vu3/zfn48w+np6wqIqCBXY96Dg2+0Zi4
gIlnyq1Q9+bZkenRmgf21BnZnYwIL9xUKC5r6CtVOCWo+aBhoMbwocJFdMmFZ+bOhmw8qQdUCyUL
emH/196psQgNLWaO99n+Trfg0HsqVPATuUW69ow4ypgFQFQwNIimea7I7e4mT7JQA0CoID0rwJBO
KHAV4DRzJ4Ad539gDbZIEbma0lE+jbPIA8J0u4O9Z4aNz2OD76j2yHW9HR0CQ2AjT7YvcRlXrewl
5S7cBG7z0qCEkMk4R3WbFrNUtn8y6VZUcdDICiwSvHagp0ZQQH9P2a3BbhwdOptJJs6Cv6bZ7Rsi
V2B7yQ7Ap4Yh75k+zA8xmM9AqPAKTogOxR6a15W5Xkx24tMzxheauXrWjGUHV8N/Hq7cIpvDi6gu
UvI8KbptSbGJM+8VVQRjqUERpAbuGT47jScZIBrkKeKUN+EElCr1UN3MGqqpD2P10jOFFtW3OySE
PrucWckj9g7vup7M3l9GgtJW740VWlQqJUgXE4vm9tIGkHbSeuD+Ny51hWYHTomIrmC8QJkyZm3Y
h9/9GzXd+YZNBGW51Mu5PoHIW3tDW0iK277kdTyV8jv20ve/ssUlclLqtbE5W2AkqDto3uXu+vIs
IDvhLJu5z1UjiijTbp6FMB/t8UprRqBP6Q5/IwkCF0KLEgi8hpO2hryy1BUG1MtnzZRkP2cCxOtp
M79mXuGpa982ZpMCLqBhWnrpFStnvyVJSfE4uRhNX+lJzsDWT98Y097zeCpm5kW7my/0cluwg6ei
UbBg6oNj4QgsKP8JHvZLHxG8MA1tdSPkk5BSJGmQ5leQ9+bXAthhDKGG/Y5f8k7D/UzfJMB2aN34
/GmkuuFWbjniK6ZCGUgiaZoA0HH+VrvbGliA/eoTtXbHCLAc6OFYpRSkcWDGtfO57AoMJwt3ehU3
/4cTnKbNOdVLab9AbNXtr9ENwQdKNZgxHafK7y0FbueiWfxwNUAKP51SkAxBnkiOq1L3KnoAdH4E
8KbXBOgU23qseVh9+D+lt2+0CAHm6nLm1MJqsWnfYSIM/lcTwV18+FQQKhmiaM4g7yp/orRQSppI
3ZAF9fBWbHCZ84Niwg3arsoofGpWYSuZrUVI1QDdPLV74ufABjc4DOh7GL51sXGRkgFdz0esKzys
WTxvKc+l2iILcEj46mPoWXOZ5VXcAUWQqQTHGIhrluQGPCwafwr3LxfTS3YM+nZLBWmz6ZLe6/eD
XWj4lHgL08IA0kg5HhHU90WGEWQK1bLAcLLwdU3DO0ve3Dzto1WaMZq1uJZinS4OBeqlAQuKtjCl
6q6cQw7bfavJwUW7bXZ2XHQ9QuuQA6xWPCIIda91ghe5dNcGf//N0XkHpQopL2zT3uqvoWlyEHak
a0AVRPI3OlwDzLTzm/ROv849JXmNh7C/kTztQddjjZqtSZOgvWWdhFI4N7Sn8+D3rLA8mA1HukB+
5J1k6rbih8L/nfGqT27sCJJoQl8ZXAleDO6CoiPt3tLRJAL/gssUU5tmpmnyGhE+rnqNFafWzidr
dkqr5bgoRD/QQ9o4tSC6AILMY8a2bqdL6AMpDDmeg2zdgEGv4lzYdDf1Kz8TqMEVXdIqb9AgQl5n
In4HO5gnXHAK+p5flL/o47S9X7yOrOIUWPNCgxVfXdZgfZ8uvzXyzDhMTIQHjeE6hedal0cCXEdH
JhsVK9xKXqJKcyIfjBtP1KcZSXqrfCXorP4WnOylp0yOH7ygrvu6UrY7XDdI99arxG4rbY45EtU9
Fuj7rN/YVPD9aJgUa4w1xLLxaFyw4BGxjYexn7oAzAGVj31iWHId5glQa5CUAPYP/YfRCwgklej3
HYNjTxC0O56K9DAVrEd/CHgjf5X730dURhRPoNHbhpjDj6YzvUsfN3y0hhm70OZwgoRKLF+qO6ur
fyn34nacLUB6FCLe19Q3Q+rk06cg/mzmsPapJcASLeHwmG/q+Crtb/ceRXKms39Gfk+ZmMIrsdtp
CO59xp8a61N8ilD65GtkdSDTJls6S4ccmLmT1yUtrMt8TM5vRxiXezjHwJTrgQdq71KZYi8DS3CU
3n7hYXNE21XBbVJj/OEDEZ/aoh6afkWRdrCfOPHmQeUzT9bTxKja3gWkpe4Dp8osRWO9Cd9fcmbr
PG0dwozrosWgjWfq9G3qf2zgJcCdRY0s73LxMS4tQ0snhL8XrULhdtzRyDehXo7zrGmr4DnqrBUh
NINsYfu80tT1ljQQn5gbKb+XB9bF13a3qjw4BjswzjZnkRAqpfbh5NpgO7M5FwbzLYxLVg6GBPvV
1IKhRczUaiIUOhBht1KDS8/9Xv165AVXctcfSvuW/ivzS7E0Mv3OCiazckbPWE2tk4+2a6Cj8Xov
qqgykxOmxVFl/z5Brmlfw8GZDh6QF1X7+BYFxZXXpzlIcjpA08OQzebj4Zj3XdqegGDmI32N8ePQ
agt+EBpMnLI6k/eEvpJwAJ/ZxxY0K+F2PhZ3nqUQ1ivmRCv8hvuaQxTMU7rnXMiNaqsxUq/vlXSc
rpxrMPW8ZLFKfezgi1JIIrwqJYgL+6l346YGukcr3Alrxg4h/Fkoq/5VHzZS11fm3pgzgbdykmgD
k/gRXhzoFsucbrHXA+CRJDz0XK3gzUOTVH1sOz1DTOODvVsOveY3jsOBHlKV3eVxwIU/wbTMdHJc
ywj03lmkgTedv7nlTdaqC1IiZuAQKezoRpblg8rRt21jToE/6IV5NOE3aZr2ac18mdiXPPtubVDC
x8USsbn9VBctO8PS2oU+TH6Cr+kD4uTihEZCoM7CfhIUV7XRfcBvgHRhzH2j13RJi5CC3UffmFVd
4wyFRHynbkB6e0h6q5AT5R1PDKK5KF/7EWISDKKcxpo8KAd+Vav13no9jyR3lxmfDCpJrpHALd+R
hSc1HU3z6Ss6p/+YKro2qUdo+z3S/1OQm8EQaTKFaYQANOmrYE6BcKsofzMlNueXd/aEN94KNYzQ
CFqO56uoc7yMznU8s1SYZcFc+ZB3JqwgHVnFX7ZTbLeHpokKJ8ESnE1dImRc7thyvFWs2maR03v1
zRGMP6Fo2uIYgtMHquxAyWJeH8/8dcVmZdBHjUmWhW2gvpINbGm9NI5d9MfqnPd5i3AtYvP3hC92
rYc26pGSpUqt3YZJjHbT8P3TtkU9z8tWXGp60j5Dmbd5FGM+jv6sQ6V95/Z9eTYHJVUvITcRL84Z
x/MQPirT0R6fiEqigL7hTEIKXhXG+KpIFJkK7HiydVT1gNvNwjhS/Vzfrfk8XHo7P6F8FiyNltiw
xOuP9SyaUcHaM2EhE1pBRMtlLEysiMjI/xsjiQl7SKjfI0//XYjJVNCnvnB/Jf9luUPtSQT6DO4c
QevcdjWNq+pQ6uv7/p3c2nURLPLwqfNjFK1dk5RXeUCUyZudhhVo7C0wDDtmfsHvt1FLSQgA/V9n
dkGaR/u5rumLaWked205zMdMAUCci2UuGyqPseUFpNUoipra/rg6FQtyvQFuTIXMq2hI91pGe3Xo
YuPCyQ3LQentdNL3ent+6lAdI297mWJ9d9Vme1k/J6tS7ipON0t4ffop95PDW4wKuIZmnhZOWy8h
x+nkKY5WjaJGIDq1VhShjJ/c0uIEo9ON6XeN+sCbpW/wABamsK7R5EEbnFD8is9iz0+1ou2BVB/y
AJqszzZI8Wc5GpSukX7ZlwRl5BUOsjOaztuOUDr3UjNsN8u6PXCwtXXdj474pFVOMzoozuioKm4Q
hn/pzpd2zjkz3XZkj5gX91K0sFhBES/Bp33VQblnfCTIxT53eqBAhqbebfUnU/BNB9o7T45C2NNX
Sxb9PrNWc1yrczOn8qnlWnz/iImF0Aa0HAdsyg6+FlxZTvBDGaGutuCsRBwiQsxv0xhRuFuzuPCk
vuaQ5OB/JU+/m5MVGNxgk6XEBNWOCmZPaTVDM7v6KcKtBkwPyS2gn8GW2p7tKupe1J8mPCDLvKih
bhT8K4z5khMBW2U5w2HZ5lQhs2ALslwKIbgcQiA/O9TagTs4D3b0RcJafRkjT5XXQrD6EGJvpnPD
cdXgjn8tfOa6pgTSYffCJhxTyDmZnN5xqWPK7FcIearvM9VzyNwvz98PfV8OXUoNgeZux+nBg4O6
nYrNc5TaQSSpQYFuXRDijQ8wNz4rmmzr5yLrTLCgKU7zf2CZv8ZlaQTekNkvYjWi+kVW9zMOgxZs
8hSCTsObndZgvFs/wbOlr8SmB1TWCla7VnNtrhvshvoMI4tN6CNy4cZoWsiRD7jwOhn/V8twcIox
L+43DaCFLro1pWq8B0uPLQqaP9LGMabq/ns5BnIWfO4rpvJsZ6y3WNG4qCyw1yEETvwIQHfcwnYK
b+fZpCd7VaxSO9ev3+1M2aF9rE3g3LM5u6ycApWXVeP+V1sr5v4h7JKC/6j3HwbOi3r0yqXdHGs+
pZolu3ClTfAaB312R4cuz4cB824xhhYvz5qO4IBgdMcH1AflL66b93j/xb4+8mVTd5nc8WlOM3JN
VRbz9LZAsEOhRIM/+jeT8pegzqbYuOWjH5+yjN4GloBPwyln1TbffsXgW6DzHYX8uILcFDIsUgt8
zgmNpSU0OwA975Z3ea87uphmZvrXXhTLh8nQOOezCcynTybWNLmmxnC28ynIGNkWbQa4Hz1Acas/
f1jzf9qP2Y6+9bEKsSk826ITAf1NHUWvShJyRX1i25iyVyzGIj82EncfIIUZjKDEba66F1He29ZU
SA+lQfVFSJy8RMcnAjUADoSavOr1vo/+1vdSK83RNivZHJ6lq6nkxpBTLsnJnN/zR3XOwbD/ayma
ynIO6RRRirEkxNCtiFESWS3vBPt/Y4qmWUqjGuOOJVNUC/mysrSsC+IUc3lOkBGWagMSDpj0bKpf
hNZRPuEpF1eX2sGKwGDIgqL8nFSkp2ebXE8XEv4SFK6gHLbIeYMWzntZSXmPEeCv/6ZOmarEb8V+
zP/a+nGhd7u97WLz4rFCPxVLI25SfyusalL+FXbGB3p2fRKvItXMSKUZLEr9agzk6lc+V6LEVB95
1n8WDQiHNquiICsEk9wGydAymsGRFqdBUgXmWMLCJPy5SULDJ+OhTHjGiK7HDzXB5vWJk4EeHkdT
0U4fpB9w4LzspZvTUHHgjb/Uo3g9sbHeA8wb0HjSZvQNO80UvXKUzEu2OxNFBHZZ1+96Ac/NunkB
XmBRdj86XD5CHBmGNSUl5F9LKfR5poRx02NbWDS4mSy/TAotu9d5gH8gWseea3kF8brmgkrWDQla
lOdoNQg6Y/eXFB95hGkfGZSNy9SdJ0BlNh/lZp+I8qvzMSLNoWly+hb/jF+DqnxalvMHTSaykrsD
EHH/FoiYLP1zMh9FL5MZjPxBqjMRoVpqZpGyxLglbHn5W8WwcZju6VNiUL/VkHwbWVIeMv5Sjr+2
Hb8qvmFMev/zgxKbd+ypS/uE/wqRIdbkId7GBKmww4RaFD47SeLCNqzMZEDdZcvqoo06kdM73LK1
9/AU+RtHILyIQq9yUB8ut+nS7FjWQiY3wt3JOE1+sIdYfvKMMG1Dwa6hUzupxLRiceQRqlcFaIso
bwgl2PaPcb09s3ukF4e/bIOL0Ss0wlLOpj+PSJu9Ktyj1xzEN1uLWOXV+LsxONaDaiN05PBLvrGM
QNf+tZ34EwVV+vEakdu64fT9TPi2z0TRA5ImVwuvdr9qQ/T05Slelb8h6c8UrBNVv3Q3ZgpeE7EX
FQqbo5dQEU3+mm4bdnxBDGcGwekoru37goKBsZrsL8L84gPkbUlEpCD1g5kf3g7uDcemLtIwv3hk
+1a2bbP5QZX4YgjrBXfN21cPnfKdYrERfRPecNEx3foDseoZdxKU1e+MZo3x3qw3Ym8gtTvwt24V
RgS96fKugfrOBI7aT97VqCfgj8czmXA+gyluOzY37yy/zimoCUyCZqUsI0WUNTkOmCXB4/UPOcVc
cCYapl+18weJs9kbdyC9eG1rzBgtokhlbKdf/5tyIxnACQwBAItY+GucN4I1VpKjcOl9woqMGLuG
juSMTTXt4tMFoQNduKfW4WmANUM7jUWF+5I1bzR2kwTWMGtNPwlk/fK1gIY+T4a3RxMDcMZ/X0qd
LVg7UtzXJJF/JRtkjTTpa20H0JY+fjFNB7vaR2i3ukccRkd3UJlLWaRJnDrq4VXyVgTbh2LBdvHp
QhXxmxLqGrnE+5hNta8afDLWbSWzrMAz+HQk7SDsR7bL5adKd/gVBOtSyLYnGVH3wiFFBznrIdTn
fh/wYLKvZLDbfZteSaFhxPZ3V17XWNDRVijPcwfQG3Joc54q3NOAdeaixsDly8ceWdJpsSWTg6Yh
M9zQ7GcrWuxmGo/ZxhpVpQ+D9PgwIjX6eWfQf2yBQ3nNh46d9GpMbMItc+stmm23/BzETf9TxlQe
6C0pjgTaqyWzYkZqTtwaQeL3WMoGIEJlJpo1HaB/eesOejCuZep0Ul+YMjj5303U9reoE4zrMW5M
/J5IhMhbPQjKC+tdiv61WHrXE1W7EziOA/77z1cuA/D9Mte9K0tv7pjWi465/NcZfvWTvN/OSmeM
Uu2p94xI2EhYaLjPTd5NvQ48yQEPnHhSEd09Y3PlpIelPknbdo6buJGTNKTJAxrAuPQUSNTfKkeJ
BT6QAOb/mkgkrSNMBkW4sfWnnF7IlbqTndllc6eqwsg2prMIsJ6TepdLtUDnHTu1dIVjzIfyBeNe
SmygX1vMBMxrF3O1OGHR3QWj3rAjjol2jo6TnH90grSjMLiwvdIuaVDMVfqlK/bljEKLmQtVQs9a
LPg2MS3GA1kh4SGiHL37g2rNBvAxrNdZdFIQ4ww74nYiqioYwBaeBhjuvy9R5GHW5xf8X0VtIMLF
r9GQROZ2w2e/wMP2sqjWwdvoppDnazwhchbXtqD5AVSh427L1V8zcvfME8O0XMKUlgBxLvbTmQPm
mwT7xhJnhlugbl3CpaF9cwlKf28K7QocWv6ungppE34ks0I9UQrT0eA5GvOObx4dxxlfXVd1cExP
1yACFzA0n/2tAKtVgllNxKuJF2JvFlr+x8JzfTkBPAwIVxSPbiIn7VDbmR8z33PS6XJ4BTiebO+8
kAdxvP0BB2ekdXidbGEUmCW3HsMKdR9j5UP4gaUiKcqf7uw+y1nPU3wFCgBDwsyrM2hvXk2EOQh5
0AlB4HHLLzAkS93994xrPHvQimnPT7Lgjl+4JFwBx19v+KFq+FOogns0kYJmcB9JTEfqF7tzn0V4
LjLHkViRTst7b8xjaAU8CwgUWA6WVl8SACd0gS0DHEnjHzFv/sESxQiw4lEKrz1IP/bZtsknrkoO
ssWSUowtWakh9QqK0r443Gt44d0Cp/PAvhZKqq9NJmBBq5ehpefh/IbQDAb2s7n3jKGNmzkFTRar
hzWVIgKSzReRfEKdz5K4Zo0rFyMWR5DYgj9iVa7Zdhw+599wV8HQu26Sv2TjivvUD1FEwjoK887+
wytyBbHcZVS5S2OY6BYsHsKSOD0CpdC4M10GAr4l3mPRFx9wyHJxrAHId+LmgKboDz0/hA30ESAR
U9PYAGBCAqu384M0k4knr58rBDCWA8pJJZC4UJd0agzCUGvMNOQxqEQvaypj9A1Oe4m/sVzaQlBp
HJJc34LBCS3rFaI7EAUjGGgIgn6pFZJQOcV5q/BjmnQllsmLT9TntNI3lYuriJXUTl2Aw3Y8hKn5
7Hxl18DXiexRZ/HvZEARLlqLQVb1COlUNnSR72TlGLMYTclsLjVbqShl9f/i0f3p9e3tHTOR9ayK
z7SIUQbr8LpgUMcdOczcFd4bI7B+7GsyQElBFNjJn6hhCqNxW1p+IImjvwKaCH2WfFeJsppV8hqg
nbkjAf8JmFGzFJrjttgAcQR5B8fkJ0jf53ncfdiG/YSWtmXL5isPcjOYwhipKlB56JReODJMmpzq
WzkS3HR0ASvKIbQiCwmT0ul2WtIStNvXUiWQDF6nQc+pl3yHLF+5Z8olCOVEq4JA6a+5Ph4FBt4M
cc2T8TNes8RWFZAUcuGzwqw5L2LBCI32QccoB4ZKLIajt3K18ZvKDPJ2PY4hkJlIegkyMzaWOmAy
hYhrnS0103j7MD1SniWWr3A1SUhFgaT5c+l2/+GJ2vQLkeYtaLguAS7tm8sBA6J+oG+6YTThl0eQ
V6E+t6q+t37/qjJzUu2A/yJCCZ86qMnHsVr1BXL+xzT6DW8J+rn9wGJAfual7LgAOSSXTdO+qAWQ
vFW3gfG/W6B71yA0QTjw+W/qknxlvPUq7SowOFiJE5IgCHsakLEULQw3NyJFGZMOBb2BOZwaceVj
/5mqJSwCSABcBaRP1Z/aPRxZvA3H51B1P9LKeMZfdfe7bkfZbP4l+5oB8qpdGmCYS79IFkPCxxTr
/bzUYIrPZiy0iw1fOwzbtLsBd8FXinwZkBTxP9+J3W6Jm5+2NyLWloqkZc16OTiyNhYZ3kG9nIrE
AFhu3nPyn/xKDIFX3U8sSx6ngZQXfoFsvyfqZcw+XEgl4g2Qlf4+zNOCoYQZxNhtF+ue3aOJKeAo
N23m7YBPLHuFiJoZw9OT4CWipSAA+6RIai2krLNvTJRtPhTCLSOLHv6kvHxrtEZ8dlU5gYb09Gs8
eUGAJpO7JMatwUHzFIdBJDI1AbWfjCDqnJkrxOgmwJDM+uNZJC6XI7TpICmAHs7i2jYgs5nfwnLj
xl37KrJowoaVdW6WGwf0TTSGUUaVZJyURHYrw2iw7XjPX7RPwU8JWWBi3dGNjz9pxQwg4SnQOzwP
XsD3tcd4BcAZDBPRxyMR1nS2HftZRhyD2ERnxZAvHT3AAD0Rv0pUg2lGrlQD5bhHw3Q9bRMCeU5/
ibD9sYiirleumHahOz34+n5UyoXVTuF0iZlK3FrPC9A35g4XUccMkYRADZL4ag3rq8ftZCJxkeJv
0t7OpnQ1nuNm3ryP8TNgDaIMYxvxIuNitUeRWS9h7tn6eWuKqMMqVIGXhqslX/L9BxC8yEIGPNiZ
pQar/7jONcdWNGGkNfYsNTXQ2R3m6y7eBunyx0F4qq4UyVyJzckxI24jJBU7kKeRobNXElJJz1E/
NytfrCgjyUa7GqzdnLc2xJHwAJPwF6poUXJi48dKGI5EskawR5Of08PUu8lc/jiEdqJnyD9WY2R8
pvN0ZlGPTyFs1V4Mc+M4WLDBCLyRpzcogFO9ty6RacCQAM5gzdg6jWLOPYbm1Q1HO5Xp+ASIVxGr
MSg75pZVAFftixqKaFDdIpluTxiot3zxHEVdle+XXX+hZgGAy3pEQYK1FN/u6E+ShA5aLuzZEZvp
pUFqO80piljgmbNjx2+ZVu2RYtLgvKbeg+dvw7+RZ+hDBGhhmMQzaQ7aGQ1xBN4KRQSSDm4xYXKj
wyniNJcAFjFLuBIIqNge0kNU8rdtrb9b7dUHHYIUPeeNq4rkC6pYpKPTK+PqXYOJguBJRTv6mVFj
ELpgLQnUfbGsY/adL+kYintdM9v7bnYt4J0fC2R1jhtacX8eSrCMr49Yipbpa9zYyWIQj4YNvPjx
kOn2RzrGLf4wYoYJdbfECJrJpezkeycibB4o14XXPM08yQ0+GD09A+p89u3ZZbPGK5SqE4PZQIZc
/ia+WhMsDSGi0qoBH6oldXC4YAPN2IxN/JyISwDaypW8a8zHFRkHcMExCN3Bqy9RghHDqTY4P3GM
AP7/mlW3qbZ16CPU5mo1Qd9tMWwDAjfOkAWfBUEYYgjkk7zTuooRdvHL3aCVFU6ws5fbTFZpUlYX
RnKJy3P3NGOzFt5BJjoT3tAyIEc0ZOYiH+0JFVvzOWxkNExmS7R9sTSV/AmbS9SWC8Rayh8glU/+
YGWTRsA2ZlX3XSN3kLDdHeB+nuGHSasaZWZRiSgGpQ0iZENZK6rIwwjxs/68Gq3hXVzYbPuKHNv+
X/SVVRZXpExC2gdWJWkKnvaqFz90nxlLlCJUwbsYrUPaWDcMGVboDDjMrJQpmi3bmXM4xnFEOwsj
cKM6OU34rrbwm2zJIsDcUiFfUNsCTqpSRrNXBxAjOP7JRRWezoZL5fI6Xhe2NbSMDS3q6JBTNGB6
etJoAX2/UNRbi2AlMwWaYX/vENzHfAq3vEXgdKsCNF2D2nSm3xIYm8E3BOGjWkJ8VhYTT9+XEWEh
UnMs1r4ZbCxegowc5rTh3rNKQosbEJQFL24lqGPCWvpiLvY8pCc+wiLl5LB4wEtJN5v+PLhE0xV/
arQHRcZI5A+AyXBU82rFSMu1Kh5Yzog5m9ZiKkgHAUbeY5Q59cahc+b03Fx/+cFVSaf8tSBffnWf
EbIDrNXXhPfN7IHBxDD10IsDKnwJpIn2/jMCIyk8nyn5LrxWYRbrJQz7t7D0BmuOFqaF+Wn4vQRJ
8plDV7RrF/3n7QSntTsW1tFJ7EqOQqIHyLOtEkiAMhPNyWx9qGA9roSMqpUGYHOah7HRCG7VNUKB
nhfRyaoWAOAnFLIj/x16mH41I0YLD6CciHfmbqg1Ovo9corMm60dacFq/XiHAzjJ9siMSkXRbB57
s2zWtMz08Az3ioYHbAjtfzD4+p8sVuD6Mfa0spYBCz1Pd88hZFR0JTin+JLSWRUoeeBdygumP1D+
zTPZ1n408j/VvcdSXkDpKzVSDaUx/EK3Isn6sFtU+OQe2EACW7NCwDkmqgCe/n2dkIiGSKJ9OCB9
mlUI5wsx7FZchBIofyEZlcVjkin1HHgh+H9hPIousnqu5DPebCeramgr7IN6PUclrc50Sx/dFmxm
Shd9uF6L/Uq9VYZJ6ilhsg4dZD1hO5FwN0TrwNJceoMfSxSJ6QahnLUgiYxTMdTYUssfhJ/TAssL
C3yfZLS6iXxn6dsletuq9F02BxlypY4qzuZJAfox3uUtuIXYhqHMXIF7d4IyuYgum704EooKpxyF
a25LaNMPy2AcJ0HW6WYVbxyHMFajbsN8l0AZUwqKsvde0+E3Nvbp3hjI0stHdu1ZyKvRCkTbBNw8
dxtNjYsaBd2H1ij6A/pOPmjM//f21emg8PXe4yGG5Tr2pRNqvlm44mD3E2RUsbgE/Xl0nnyTVejd
EymP0cPCoryq1zzR5LtKakuiUoytjDDbBTVMsDVONvdJy/6yi48xZu8Mj0fs6IAq/Bjm/cxEFxlF
cCmlzKWyn4ty9SczS7voJmaef8Y5cPNvRXvwZHbSlQpv5PdSfvo5tTA2XIFhvOKX35kUF65E+wFZ
W2w8e1jtP16iBY4wa44x4ITyOQ46K+x50fSmlfo1adcKhWJdf9bjszUAdrzOSXVhQZV9uyupbs9j
bKjyyoEXhbo1yv3+mB+mJ514CKwcvv4AhIDiFBFfzKXyAYNrADUJS0phhyXmZIb0g/Yiy4e74JLZ
ZnYOOhKoUVHif8m8CMR+XffaB2zyxV+KX18RAgxqPgSTJv5prmKcZ6iEEN2xhl4z1YgP5kNfknW+
gAFL/Sfem1zkSqB9U1tfiyC05cezQwZlu13febIRHmHMMxrvOT0viNCKajpsLV6RkQC49/X+xmLC
9Fiw09g+qbNdWUgrawon2B3LXHxbTKCx6icQK+qdSN4uiUsMAPKZbIn3Pz+z5CxWI6kG5/wL8irG
I0MsmYpA4CMY/M0OeREUybqwnsvO535HI6X1G79whlKbdsq9tWah4v59b2XcspS4ijl7PnZ/pIS3
N/vwtbU6ufzVBzZ5uqA40gZHVtBheupQyFhb5BQJ9VlKcIh4LVaZogsM+AaygAIKNlcaoBTcFvwl
jYD+NF28HEUnTy+0A84obpMLccCiUAmDwVj4OYv2JlNxsQxXYnneyfs7kgUPm3+k9ECdZVt2HDkT
fdAezktlQwtx1YEsAdaPAVbc1uwX0ntWIiPwTWmu3HamnjS0khPmgOiheAGNtmhaKJzifsd+BWuR
3b3roSRTwZpHTXsi3xKW3bFdSubZQahLw6+qmRZP72UAZR70g03rYgk8Iu5m/fMHhz/eknsM4VB4
qKsA6tjY0PHThsvXQmQmtQZ1vGhnpHPMsprU+8IhgPPEkU3YKuC01JabB6Q+bkoMQa+Fqqvznnoz
fdN284imaH6zTYPVkhm1tQOD5KPC8+LsXqXMMS4wC4DlD9p9cqzRGLf17qlhy5cP42FcWBe99ooD
Y51DFf7L995dzRMCzInxqTX7oep/ryQIsAW+hC3gMIOrfOqPO/nvuP6k/M7gp6jSWfNg1K34e6Pi
HgYZlo4WxZQDyc+Bu+B0WM3kNaO30XFwUezXLw2Yf5AjIWxFut4TQalBURhEHA7Ja48nM4lyeKoF
e68KHs3e2JeIywNuUa6IjSXzaYt0nIMIB1KI3VdGFAdiy+hyX1UsmHm/tf3h2sgk4M0n2/sT+lRd
vfpe3vL5jB569DVTKv/Ky/oqQMFxuSs/wgZ/Uiiios90OQsG97j2RDCuK5g30rSC/aGl555jWa6T
Gu8cQBTSjxKbx/XIM6t16ZPLTsqQ1XpSj5L/mfDYG+KS8LW8tjGYmyxdYBtVh+ddD+FshKVpXhjo
IC+z6D6eqtszkY/CPfhr2nVBQj2OdvWAtXlCmBpG94oa06aopSyEJ6dxPmJHgQ+AY0HMeCJnIBhe
F37JSUHP/6enhqaKbOPyfUM+TQQ8l06kulQ6f86knUFSRVm5huDr0w0dmUbk80fIx1okS1Tn+e/N
CllxVowhd9eafC1QW+1Al8BURkf1kZFiPB93NLF322gaX1n7M4zT9oPh0/nHg+DrIse+zAXyrvel
cVkKLM2Hr0jZKMJuzBk9cBu+VLXDDHhgjnMxE6Rl48PS5ClU8rHpCupoFpu31Kz21shbXigZZebU
ne1yuPCSui/COBT/5aW9UMABQafAGBJuXP8Zjv/JORiFTAOOqS3qY1e/40k0Hut0SL+zekl5pDLI
6EF+eMtmcrHiRx2duNMg3E+CnpS1e0vpcHR3QWcVaMdamErevRqUBae1NERteXatCp2X9WkA53d/
ruxycdtqbIltyMdBHrYGgW/bxnt3BHgJJP1apxj6ojoPN5/Kns+j5K3AbjIpMDHnBGfQP/PIpLgW
vHUKZSbSsQfrt+AOowaZQCr/Wwfox8awKvuBTIkt4mKBxCiIHSzsNScE62A04DvZYaitDZjcpQ9B
WKiX2w+sVHzSBw1cr1AC+NhtEZGQW/gD9hwTQSKuoMe5UdQhPSSfEugH5T9mL1HSk1jj9EUWAvmu
VlJnjQ/uRB5dH8wgloj18OqFjNG1RzhstdwBYmBxBCLkhUmfKrzf5L8z1Idm/PumRP+CzZKDO63T
bt0Y9NA82Q4JF2rhYhXsXFJ083/O/iTSep05qCYny9D74sEx1tebw9jOEzKBWa0S19QGOVEx+lpc
Iahjw+EeZFh5+QvMRJlrNNOeL+VHhdw1Wtq++rXJ9556n0YYfbjR4W2iFhIbLkFTluiTh9ukTvg9
F3b3wE308XEi8QBdtihM3z9WuU9CCSoMvqYELEzxfPCuNNOZFky+pjzrijH9VCvk9xE0e4e9A7TQ
s3f5AlkiMUscishRIJv32zOQ2KBCJvZBv9DUnrFbRwg7peGBwTmy+bpZfYa9/RGT4rnTZ/Iha2CU
f62An5agq80fL9qti9wLXp5WEQmOZJnbpWU5iR53w/2dJ16itGNxY73iex8f69acvtxGBq4QGzm6
GVVmSaHhTCNQMFwoILM2eUp7Tq/e97/r+WBlGGhcUPq+/n1dQUUnOUzJG2LRBu6mILjXHdHsCVWM
EFBdtVKrZ9tjw9a4jOvH9MdrL8OP6RsGvReok55r7Q+LicsmgB9WsknJ0IUqVnFFJEdGeLlOWo/h
cICHfymV/jYVtwsIoliqgEbQAV8pfFUaHrJITqRo38JrHDiyOJI4nsHFsE2h5XJCfxfdlWEHDaE1
M/vvGtqIZMMDcQPpR2V3J9oB2XrnOfJiqUAx/Xv2E8s43NSG/flfqXxx9K4ena5FDArz8xtwAZqZ
KBftk5064YPIQe/TB6BfJhvwOWLxhK67yOjyYD1UhG/lKWXRKZlHSCh1ZumQH5g6+neywupWuKlg
Wm9JwrE9M0rBNLi2uu11tys7F+7AdGMYGsZZydhdjH2LAwSj3K0x2dTMBuguVQ3t4nkSlWvz8ndu
i+wRpJr0DiWEciwq5SLQ+CWWhfUILMC3sO4y+MASebK/n582ukzWf69CE6a0ubaFPwAxydXs2iS4
naa6MSmzTwB6cX4X/W90GqHBx4hutQNFohz7TuuSNJg+Cf7fhJZcCeEspjKu1vtaqsDUkx6XDawB
dZRye8zaTahQdYE37EAxJPDhFbO0YpoxpwtGR9xrWD30l8Vibp9+uBmRzd1fTWtQUOhQsxnBIMaL
h/Qd3QYXJQYy9F1TdYIqIugZdcM19xM/5QGKOwkPZv2UjDU2TUbCIMfpP1lqMh3Aj9x4nxBQiKYv
er8qgSEnNpLBRr6YlnEY3P+EkkfHOJk8mqKCTDHvYHpGMBAEsHXknAK9YWEMVVWoL+V107C1Lip1
S7Qf+JeEAkMX7FlWyT4ItlXHIUpIDJ44oVuhFL1G47WenXnjb6xerkp5h0y6bM02U7ONmdGNR/tJ
0V1zeMyyMdVlR20MbP2q3eJp0rFJQLILOV9d3VWSgD9tJaZai/k4L/mr1rWxnCmonggseYECslxw
JvGe9KmBi4s90T/Sjz/ZJF4mw9iLbIi6/IjW91kjUyi7hpfSnRQIObOCdhRJAHg0JCORkmrcUqNb
NQ1EOFGSRm5biIIUu3Sf543bZIEnMsuG02OfdRgUi56yw+lq+XxXWqNJohO1FqOKn69sfol+mYHr
1D2VZ/Gk6Sk+oNlaFFaKY1G7PG1LAEeed3MDEYxzN12LOmB+7Ybs3xm223mRS3mhStx+7wmJ7Cwf
lgslZfEq76IXRXKfQomrk9suTx8tb1wVNCGbi4NXuXNplWwpUShE7enSTfp8ZzvYNb6emn7VxA4b
wGn8+zQm4alCjgZcuEIScTQGPGKIdMVH73TOg6/4lFIYs+CQV26uEUSk34EPlNwoQp1gUPCd6AXE
qbkIwbZhZkm5ZSFDAJjYJHY3jN0IfYCO59vvbwFEdSR8EoQkw60uLCCddsHjuYfRhPpd99KIZYJ4
rpMzICUHgr3ESjeIh6PKu/iiBVDeb/PwYF9DsXjsuizJ7AJfHQ2o+btg5C4D40SK9E56RnKuYvDk
CRzbMBslRBfBePj+xOmo7Ac1zC5v/JOl6NGIqazSLwDwqI2P8G5yUs+10Ot+BAwU3BaWYb9CWooV
KtlEnngC6HuIF0BJJlEadD+Am1tPk3giUix8OvMzbZBYp+ukni8MePpJCKdqj4pxzCk/iGqwGUJD
sywTyXPj6I5dMBmWgnA7jidZ/300mfyDGpEL1KpytAwfuN3LDGNobM6BFDhORKkUb5ruy3iY5I0Z
IhBWMb7FXF5kSInjEFJMa/e+Q58V2OiL6Aeo1HhW8mR3Ijm+OEkXU6OVkwcanOgb2giV3BYChKF8
hEM5+KvJi+Hyc/QkhQxYdWzzx0iKzOGZ7pg1jdjFJkLFpo2Flj6a6Cndwq7Y0z6PeW+fIqWQUl6n
PIs49d1AG0BDeYboIHMFh/KrsGwt2zcYGHXFCIuZ612XxCOGwgP9++D4JQD/2O7V6aRKNtSYddIh
afy0A0gZfalu4i4VjplALYUvCpThfz0pxZy7zBlF3IOOuP6/tthhSqxaxQA8g1DDCK9uJ8+m74aK
yQNejoi7rbd4kvdZw7U8oW2rhDUCrrqicy/7NscPe2z1tP2KzNFN5ca1K3VEMdv4aUJZQ1epQc7y
mxz7/8/Dhe9v6KnRYIZulkZGRT/1n/l4ZvEawYwEqPPp5x9UG0FGEzKwOGChakfNf3Gx/QkGtwVs
JK5iWfdiYW0TLoom2nYI+836FQaC/UjyN5I2sQNVemvnjFTd4Tkx4WA1NVHKlm2RcHahhsYK0b+9
h1y2wXcsABYOQlUG8TXADTQu/19XqyxaaLlOU0TLcPQ8NAxoU9+5QUJqzxEtiaSxie0wf2b9hQj3
QSRDdoDdH6oAB411Y6cp/bCxi9rmcUNcX9pin6/s5qCLn/h8bF3P7pl0QYl48At7GQKUp9Rc27JE
QSuYB5n5AkGFERPK6hqCfdCwBLGVcli3LCMgGjDAj65+A+HE5MVWnRsRRIqwRVytTo7U3t4Yx8rw
4r5lQBw/VslhoZFl5poQ4jEp+S7n4hY17w54qoEola7+/ocQp6R/OGmsVRzfeBmDerodhpntJv9p
q2xhM2U+Q0xF8+S6nmpioam8M6ZVI6sszCguxgo/WDLbqHRqRvYRONB6RKX+f5NzYlKXGaUUlNyF
AlPzzwlMqn1NvRgcCYgv0dn6q89iyWO5KYX8zJ/FQpwksM9uaItJe5bXvxBwPGgn/Nqns/swos5c
FrLfntS8fIWlBi6+F8fTw3UhBT7srmtqG223yRlLvJPqwT09ngld8ronoaptltG8ZYfvPT8csC33
dAT/DJgkUXa9IfDgu7Vxmod5KQ4FcK6cUmdMYsZgdhzmIvzElgko4f6IlA4gHqYvJXw0xeT8r7DD
DvERSdmA7WGXvcRGXrT0u21R40VIs1TiNh5D8pp446j1ZdPU9O9InMTHraRX8/FjMgC4er+PDK3p
9tDrR/Nu4w+uasVaf/lfc2dRMc8quZif4yctdc3P56ZxZdOL0uQ4x2b4/7ypNPcFJ6SYlVbhFHDd
zxGdp5l7+QKPEkifPgthRG6uu7fbsXn28a16Ot8+z0ec95qH3lYkKyYAvHF7pascKA6fvmwSED7I
Un3wIraxmb4BvvEeue7RlaFb5iXThMolGw2/1ENSNKk1ZyNTet1GgRSKbuUZeM7fWUsiU9zMGzyJ
SFVZEVpkyX/MpUS5IsIKX30Af7/CcWeqD2RFTNZn0EI798wUyB6AW+BqRWuQSdKlw8AuVpZWElmQ
dsdzfA55ZuQOOpSO3M6JSuO7QrBMcoz9Jp4gMrFJhV7gQCIZnMo2OEaWLcJ06nL6+LFgZpVFPQju
n24GBzZqqdxX0WFbSy1uognrv9cEGqJrsxAK3UwRujaTttAS1koi/kOgWAvN/NA1UY0r2rDnChmc
yLDSxM97DvS5qVlm/k3vDloo6tshO1hVtBTYu3RibIH1YUOz7FqICD4JPD/DWQnaYChvCMnUkllB
fReky4G8up0ZGm2OzZePliEGlr4QESzoNFI+8QiCM+o7pDg+/SJkDnUrRYnG9SgBmyfH4Ixp3q7e
/DJhfNzRB2tFoFDDhVLD8YA3xiySE6ovRIPek8nS0GWEDj01xhBWNEGH0L/wpd6k7ibqS58NPFJv
Srw4kcWJrWRqo+EyUJrzPzxdshqnkQOcf5b0gmVoup5YpD9sa2jgadwSfUs3i5Xb3VFxugm8NfRa
WqPsO0Yj/FYETkIGxuHtAkvVhoaN7aN7f2lW4qvl05frPQWpbOgT0PUyepwrxsbSU1AJXSs1XlSw
01uSTgF/t95t7f0LfgDXMPPF8lMtMb/ExT457EPqeu9yUiyF9QIaKxQ7goKtGV/Tln39MAgLbrT3
Yc9XR35rfSmzxfij9YPCSHdpxpd5LDT8aTnD98OsGXchzF/Yz4bvXdn2cY3rGe14X/t1qAVLA9gk
dTAB1tuQVEIwl8sc7i8Lmam+yuC39O3uR11wSu6lP5B6ock+aZfSEwptM+yEpHnZ4Z1SOR7qqoQ+
xvL4z3HExODjOSCHZpGKdgii5R90G56bKg3G4qRi8Ss3pkP/dCofORdtON/sJpwKNrlXd6TZy57n
v3ZCOd1DdMHaxkw25UK8ZJzudiMxSXIdG3AIl03KWj9uHdYyWLF61wykm5wMn0Zh3OyCqib36D17
zKQpi9SMg8uqTTy+lll60gxyStXmZgCsMFm4LsoC72+DFW0DpqWqud+hJLviD6OOC1ExsjdIoA1N
cmt5ZfvuUqrPRF+ze8bWsCh7hLjyhHrUmWLvLdw9nz0Bn4sjOxV3e2/DrLzRmiorvcdNxYrb8+U8
MoxYbo6KajK7ffAFHR5JK7jT2P+3zcOfi6AQNe5AqdhgEGAuIn+trEkwbDPg/aYSDsn/7K4qRWNi
u42ebDG5CJERfN81esvl3rT5QvaQPof1KcjtjsoYN+AlXWkSEHlF3Fzb5coe2DdkWPTSNwI/y9ll
GywN8hRwCR0R20PihL6QHg53BpxnCL2tLGwLmtky4/Ik1m9XNoce4rjDKteacFZ+LFaZfqAyHaay
PSKcHApA6BnMn+YWbYuuiVTtUtALn60H5hsbJDNWdk76SGGnV2ilXSQkimK9BhzZGH7e0KLY0Rok
JefBBeY910DUsgxPCRbs9K5aDfTJO7O9SibDUBY9zFFqajASjhXAgkh5tnYykkbrLFIDSeYYYA9C
/Ul3i/c6TxVlMMHLqK1WTy6TBwsfH1oD002Dnl+x2o2599VSABc1dZDraiI19QWrMrHwasHQ6tdT
UWfR56d79YcE//cLNUoqoLpe1a8t1msJme98258g25hLP6u/wpPrVsgyDofB35tf/ZcHLnkQjW/p
6TuejngNO46XNWQs5tFRaqyoaU38AnPOWtFfI4fRaJNFTTLRDH8+X52sgi+YP3emRyiEGkQjh3zc
nzsWnJrf+ZdKHBphS/8WcXT72LAbXQHZ1BYvyS4eAOPyiUN/5It8daytN3lrzBlT2hd302HwKYWK
KNmRtWGN5XthtIteTBIAAak5l3kfGF+WaVx05cOiIRMi4595knpL1Adu/MlTMGiQxNajtuKnGq0C
zhuLFbjV5TJzZklcw7cUL0HKlSsL83D1TbdLBi4yUjZt/sSg7L40f10xVB9vu/tNHbmCCG0Lynii
5oWID/r2Yg6amV3xT2l/Yu4AbTWKiIe/Ci8DN1AnSiRKUK2uZs2245OwQuMPe4OR70EfhX4ibcB7
Ujqi0JgxH3eQSFrFhEpR+TLLIW1iP/JpgrkcRUd7GMD77E/tI0lzTgHg27D6HgD0VYDTyNE30Ews
2MP6x9cNnIXrfXjmg1ggJ0h5sWQipowJ92gOyGLK6DiyvHgdktcRLi86bve6KwHDotX2K2T/G+m0
OE9baM75/pVwLwWG1x9sSyJAOU7slC7Y1cLoRKw5Ot9ASpgm2ZdPQXZ5QUHiKTy/bCDWf6nbQmWG
vlPOQjgwuldlDrr6xS8JctuvhSzI5v59O/ynAFdC6kS5Xdw2qCawn0hZtIyFFAdYgLd0vx/5EMKF
zHO2TlsUkLQHqCR2iKr4ettYrkULSrex55/R8Y6sdzl4C72VtFmUkdP15Gsv7fXVnZAkUWqCg6Fd
hPynK3BehJpgkVPRrUYBhM0GFlR4Vu7s92/3xkYxD6iPI1V24/1ajqDZ/EMluKVlQsDlcZ5PiDVP
/5PbPL5c5VujIk2YOw5H9M/E9nFKWbNWmYFGYE1pkU6Zc3F+8LRyPuHFRK2f5AQBIf/qEhSkkwYQ
KwboJOGWknayqdeVV0oN1EWRiDqZ8nmUJXbnpFXf61WkIytCgWBUCYYTLA+vuA6xEPequ1WEOkZ5
lQNeMh8tUXd5si9A4tIxAnMM52FX+mOl1GyAa8Sv8U7a9kh23VjVXqulbFKsy77oqe7JkWlZazCW
sT5AfgNhtobW8uqD5GcwxgQGS1dD1EtCqhqcVWmhSI5G4Dl72GpT0Bdshd6a7LhS4yBGjkHcFEmk
q1RUjeNYx64NXEgDyuC3P3Slpj1J2otWevzxmnc8fLKT9tQ+Idw75w04rqMIg4yr8/8Ex3YMBpPF
JeGBoBbJM4qqw74CJ8fgie45xwpWWazCgqVezCLSKi/DPemi4Qno8KMm7gYU5HN+uvul/lBs+RUo
ZTFLozGlof6MvC1XLprF/NlYO8RacxfoxgHpvy9Boceg27QfAH6TBX7b4LdFOaAyVyUju+BjSTRX
UErVgejowAp4ZhH5a8yZlEnOrKxWH+UHdZffAfW6tko/OO03NC8ni6JEGK6+dTqs2ZlDr+Rl/mMt
PT1/eBM8OAqJQXbFIw5TuwkeiBbglKr/5L7HXdGjikfQDuq9x/1nTD2GcQ8C2IdhzSbGApgeqruL
YyHF7iw9qObzdek+E8NN9iJDmow3F7EOSbVNWKohEqZ2kKHLDPk0qr22RTZ3x+gF6pLhQEY51LaD
tHTGQCViDwcOKS/vKOSDRIeluX/YLQJEHTp3OG1A91gL6jDBeun+TKRk2U8X0lna98WUPSg30t98
uv9g2bASPoLY80/TW1dtFQxL+zQnola1FpxLQa1leQUMJUbPhBFv54fiBq1yEIr/sTjxtSr6U4lE
uD+AT5tww7fpEMzIJozqxbn3h4lV1p7gaKKq2u8xNrt2wtStnhcIFchHPZCmmw/lmilO9mPbUOhS
XIEefQmzmqaDZd4my630V4KgaSrciBx3kLiGeAPRajzU49KOYYrGXfKEHh074Sr1ZV+ge9AzzXo+
6bpofInIr/Pm2nayUW1mozz018Php4DHZmPOT7xPmFsbNVwOYx+tn63kWwj0ZBndsN58P8yXbUig
Hy7nXM6q5gD//P5U8Gn1d5sjAPZWuaV9vvu07SkOUIRgjjO9aVcVf9Ds5OeeXaW4/MiG3UXFzI19
BuB2/MlsD0EJcxwZfPuTei0PFgXXLrnRbLoFU2icTK8+w48PFdwZWjsul6zhEWRp3Q7D7G+0Gk0T
NNj+UNvofoX1xGBpUMFt2aTxNFoAXGr6w3JCVj1UORHfLdX9FNKd2O2AJwAVg7BL7I4ktzhwhDCo
obMR2b58QlAhrwnC8mSvhrwJ1/kE97nnyyI4Etgp4JQLw6/loL87imrhlcbFeyUkR9yYyADs6s2B
vyItTP1N0nUW8sq8yKSI1GggwChLE2r8NeDKG5C3EWGcMeJvjTOgutUkJEBPM4BRDIw9sdKlVWSH
EZKK/0MVM+GkEfNUxUnfhZtT1iFeCE4a9HFoFk2Fn8pwO4HQiYmvjwkpTHkY5GCMYMgeLVky+EI2
7li40MNDwqBHsWIs5C1WYAbIMmNf+ZT4NO2+guDn2dfcbWSvDMKlrOV0x16D9RLzdiVlFzpe9hIF
3Sr1qg/XlrXx8Lmj1OMU/p6eNkZX+2xRDTlJmBfVgBIa7mgjz7DjVtlN6gUvyNyE1E5RR2h3FNdP
6VyRmz2eJhvkFInNdHNwwov9Wrr//XEJMHMPotLpqMzlWDwMUTbOhqH4OqBTd9197n2BXT5zCBtV
BIO4+DsPJtC6KvodAdArhLC8zTgTaqck09puCReMRLt3socCixNDn8ekOqiQu2cyl6vGE3jtibkA
xaZ2lz0qHPq7iGYPJlLCYxT8X0a3A+AN+CNQCyfuxm1upci4zjU11YxZfOAlhFw2t2yQSlh32onc
t+BimsCo2kZ2r7pLnCJCpD18kjTED/+/yjoUvjQ1JVcPyaHkF75c+80aln9Oi5+U8WqMV5pHjSry
n4U1wUL8tJJFe1HsVRB7tHV00aSXgrkskI7U+efU3d2/t1QyNVh3N5pYOz30ks96Fu5ACJTrbEc9
9cWaQLXInStkBN97nN3VkdZGzJXGhYBKM1nufWSdnIXBQkIlb/lnNzDNHt+CiAvV9esQzh16IYd+
nmtzrefAy1e7+NdzI9aML5db96I66o85Wfk7MtL4m+NC8sEpC9B9v5NayJW44cwE8UdBO6LYiz49
UF+4ny842NOfKYf0qO7Zht3ZT44VkEBqh7t/JXwruTbhKQxBo0s/jbMQ4e2Y5RjV0vxatchkHZQa
KBjcX6gby9MDFiSyMRbgSgIoX4yntddyyfMlV/lxrXB9rqpy4YC6dNgMYymLQj2qmdpd/6K1NTI0
kiBizba0qvXrRWI11mfzMfmbJu3SHTHMYT3W7VcTSPU0Sxy3Z1KZJNhJjUknSiiotlLZ99k2xL2J
oOLputJNOj0d7pQYj7ManLNk4aBlKkigT1xx4PqzWndpH5YN0VoGnzDAfvbJ3cDAJDl5iuQ8B3YO
RMPunTbSi9wU+0E3aZgva74NAkajAaVYFxmKZaUUVOpqCuRjyoswNVh8fJji2MEozhoEUP1q3v9+
H4xxndOXIFChTVdekYCxilMc8NnqqUeEZ2v36dTwb039eaYmiaitLaH/4Ph4E3xhWepHK7e/snfe
QINIimBSJ6HbCayjJwBJsm8mtrGTfmVka8NLCdoxcjGqehRSjlIlUEsMoXOa5G/MUPqWJaPsFI2g
Z2Hmy3gAVVDS/G4PIlVzuEJZG+vOwUz+jqXFGIiSjIbt80voMrubOrpsftbdBh9tmFpCqD1/O9KH
Fvwg4wI28BQADjsUH6gR9pMn5qvAPvS8BG3CAO1tVWFooWNGEqg2IdhoBmGCbKDMyvCZgrqza6ud
x7mzsFNKxMHNTvCS5d035aHjHBy6Z6Fs+FhxmqgS/kX6aJ21QOKV85EaLamTu72+gLeM8Q3lcZRv
gDfH1DNaYaYQ6vlIUlLbBoxe2LSaP3ayrCcAeR5C+hr3jB2RLju0AT5XehFHGFgKw3j16s+bbdbj
EkONoJygE2uZFgLcVLwbgfV9AjRTJfx7ENtxS5YBxK7YFq7v3hsD1n0jAFTnihYsZ8oDsw24C1cQ
HSimRM0OJ46nNIJYmFBa7GZ89W8wAYhMfd3+5HTzatqOoRuqoXFUkVNCrjmm8QmtseTIJ1ZalMVl
+5V12qX2TmJqdP/ARYLXWqVE88ZCfnRJaDVfDUcaOHDmQ/1A+4uIxUwe6T5YThqq0astUSRUhktB
DhyxW/bValN9lKZL+iMlyvTV6Ttlp0P9BZ52VKksyd8lBm+MOwqe7HnUQ9fxX8m0bp+cEaU2HKyM
iaay0hwT6WcNrB3hmPnHiUFdC2jfFlIS28zCY6xqxz34u0fCUP+ZJDx5JHWvouWY3o598oSjUsWt
0OMuXL7SL15AMQoDQEHM8vk42SLJPzvH3Wb18bObMvyE4is+m3HlH2nRYQO4bpVLty5Uef+sXNoq
vpn+uZqECcKW8k/0Kh7aeUbMBmTOWaS+o+eMVEhWBd58j1rBUnoXCk6v/oQksVzKlbqdC+0yYXqr
Xa29Ur/mXcFQL5KGC36x1z3HuDF3frM3XIKWBpk+O1Qxh6Vve7s2yev4l0RT3tUMLtfWnd5WxeM5
tvTa1488OVfo0Qb96vj5KG6Nnbyu49iLBZKCzXwkme8svsWOa8uAWTOlpQ/cyKzIC3bzlkhZxbGy
G9x89dIzvvUxLa8y/CstFnmFE7afVDHv0N4HB9Br2tFHeHAlxwWNYFVrEH0ciQKiBCkPt6hntpn5
AFykWEvcdkJdDZtPCDhMjoPIOA8Fj127zexXBVtMv3PhLUQjEPwkTxxXV+SzlyimfWt4Fm/wINAs
1EbSajBYhB+sQOfcUuQTe7NEhd7oX4BGKAMnrj73bsRsPQfKXnO9MFnVsV1KI6Q5gRjBOnonPi+1
EWE3OacbLRiTU0SuIKmj+Toxc/Fhh5KyOq0KE2MLBm+nQuvbxT8VOjeYqHY5NbINEsYzADCAuNbr
eV4bOL7SZiLnBc3JidhR1q5K+viC+3gQg4SY2LQ+mPSg0XMrJb6Re25zRYRfsN4QPr6oLnIyfQk7
4n7FBk+eIjPhafeStxLxwlJDCJKKR6QMmvAp/jWd/w5QI1YtINbhIS85trjxsei8JI3OoVqoAxWE
CwT2+teYtM4a7EY780L2ZIuYVYJHHDogx1aw3DVLjHMymNkWQmK4ctefw7+HGIud6NoURAPlY+Xj
MyYnbKxEEH87ZyLJ4J8qayuh9OdkmB0v7QBSAcJYlsqz/oRWGbMC6bbZCQHgdwtW+UaSU2/yQalV
maWjXaQ48SrxqkgARmUsxF1+zN+FjVcSmb1yM6YmYMbdXUGjl+/28cbElf2dz48edukOvxsDxYUK
IM78iGNiWyclkTgoI6rljUbbMP8mj7AqQCz+Tc0kRG0fIBXgaFq6ooVDElDJkqdkhAk9tTifBP0r
7wz46tod+P6+OnlOacCzQnnjG49nsukZX33uFASwZav7JNzXT8SifB4O/y7Ga7yC3FmNg59xwK2D
d6+BnBUtdKp8yLY+V/tLusI1A7te4I/wEJFoooNXUqOdQ5YvB3uOJopxs7sD71U2uVNRk/poPOD+
UpxLLvhAwqfUEiE35/y10dIcRKt9JKU3M9ppVOB6BQF5B1ImFNI5gaxvVZTBWL298d6F2E9xjjkZ
L5FOKaRQIs13pNk5IYnHW199N4KJdyiRuSNZYH+wcOsG/9TyDhF9OKpVLTuV0QxaG20VfZswJnL6
aMB65kBnDqGJQDA7h+HEqoX6fs43csZCowlsEhpx35+8R2eJ3xv35wZemfcEQkVDvm4D+9RAOLUd
Im7LGKf5uFIbZOhWO3no/foyB46+qj6TBopoPgC7F3UwW3EER8thI2FAxH9fXhF5eZ+zzwuLlf8u
LgReeNlXhaU0Pwn6LM/eoZlSNzUDrKqkxHNCpH6Z4l2dXQeBNYRK9vY4pp/bWuLZDAG9O4NqKly7
7JvYDscMV8Zflk5/1o0Q9+VzVu6mrxypEwODrPB7bCq1DLSkF3NMkLwaxdzbqC3c5GSzpNzIeBOI
HTD+CIsqaEmDzr9uLnc6HKJac7Z3P5L3DH+QuAaTxl3TM/oGr7I3lSVu68lUoYXLomtXJp4xRTvI
0xQb/hNy/JzPlIf+99/Hu71tAsh/pLKPdLNIAe/P/HVtzjZI4cVBZlQvmnyK6R88gIcglTU3ohx4
HecXwLfYOwpfjwVy0bJCBuuTu/FbVa9JJYQvCkUGNdQNdfTL9d1sOTVfIxXK62wF/qjAaqmS4x+O
LmnbbyTscFxtLNJahqBYKa7LaIJ9I47ndfGqLZaecH6ylblWuLwIYnhdtZ6MXxyUvPsqMfKCPSDd
DGDcc9y/OXm9Wv0oZrKtzqXa0qDdNkGPCN1AJePkI5nmPRIU7KHB+ctUWad5Qhx00T917q8D/+IV
Wpm52y4FJJIX1BLaOR+nC3WFuBMg0wirDfKS7eiTy4oJjfTyF159lRjHEmRhoMFjSljZRXUnX2h7
p4DfQOD7tXKtX5ZqRxMATfXva27ErJGgjfkCi39oIVgGg2QvHbqIlI37oByCtXQz9rwav7jN3AbQ
hWnS9UjXec7XpgpmGZj4eY6MXE0uVHDZT5OTQhw6ohzH4RUW2tfgm39kFuCwqMyGgfB39ovtjjOz
IwMs/u6NOvw5wOUI/bPhQBOLJtTNSOyokjRh+4Pf7rIPI1aP9kNUjlXhfD86td2ed/jiq5YvGURH
MUzadaT+SQBAJGXHgmGR5H5DVa6LlON99ZhDsPB9DSmDtNm9q7wz7GMBj0zDtoaIc8Qwpc5Ye9LB
tvlRd6X54N8QtSoG3Mg5askGyhOmLolXC/v9NkUuiVwo+0PryEdeIgRSd5YaDijUuKI8rH3VBPyN
opuN/Rxp//kIUdx87wQO+UHaVejqSmtm2zKruPoJq/jUMdP4Q5JjABGw1qdfgoGTLl1hLEI1HgQu
GYeGA4zGO/HxTfm8wy5lf2jx0eE5ct1ajDj0waKI8lcHiiA9e3ziEdo8NvyKFTuYiWPJTT6jewYE
EJxtzZz1ejtnomNQvnxV6nnTZt0H5FjkPUTQBSPxWDUSIibavTCU618ZZ4tsKX6HRGIry5AutO5G
btiVh6NdguGTa/HsCrgfODm7A3z+khCHYlVZFXkbk2pa92235/AtP187LGNPqLIgN+j0qBV4LyAB
Y1F0opwAKdWLwU1kg3wJndqoFC8CeqzrhahXzSNjVmE2c4BHZBVGx04qxIWYWPTUxP7jH8//bIZ7
QKqu3uTZUvnZuR+uMSz5FKqg+rslvWpyCPZfB4sCkM20Fn6aJWBHOCTadtNu4ue474WfSU3/XR/Y
DXth14STf4CwyDDMtC3zLPo4cXqA/5ZXsFN+Z+dPWODQQI9lKlQyVQAEtnYb7JHAnc/Pcwqw6nX6
ggfxqRsdixkSXsi/ogy1h6LaNI1j3k8focGJBP8vzbw/NtqVe1fCOtdQNGLTbNioD0fO1CaEIWr3
CVJzOJj70yfbS4d+vnz9S0CL7RGduvGcL+Lh/8JhmrP4yDRy6X2RsWSogTSOb7eoVniGGQbcE2To
3J4ryXdZLKAxQpIPzOAC/vpsXkpf9RrbzuU0vbreGeZnLJgaBjTjpBknkZocmTB2S+/8vWsAPbAy
3hlXRjtnlxcT6FVSvmP9o2NqkG7d6T22Z6b5omuEtzdet+yHl48Iq4Us3S8p2vavy4EIk8RhJF9s
3iUF0aAYRrNRUkFHslWyILHxIs50je/Nbqm+lNwhjH8MvFGPhLTiJ7pAgkkn/Dcz6eJrM2LEOiDX
1VDpO2nhA32FvRkrrkEq4Wmk2Xt/80zcW5LIRQPErmyuilBao+P7C1K8jMi5/a4ta7qL2GkaR48M
leJFta/cjcfG9WfJZaWCgFcqNHCtiIO2cNEdOywCh9p2VGlmFh3+zVdf0UWlfTc6i/S059G6fGyb
vOp8UUu45VZGtzaF9z56mwNfdOtDru68RiY2wN8c+QC+qCCyWy7OftPTV+iSO59mWU74ruoqzQvU
TkMAveEb7ZBgO60yZzSB1v7BFuLpRWd+dpHKCImrf9WbOLhm5d16fqRizjKVzD8qTUEP4HGS45a7
Jk3dkQoruVTei1KS9Bq9UcNfNNdNHAubsKA2GDlI3RVT6NJFMfc9EFgMxR4WjcA2Uv25gxRjBFHi
sbYUdg9HLySxiNFzTbtRrGswTv2fhRojLsyYTMsLA2PkrjOYv4ow4JkrxuT2X0NoYszgUop1/WpY
xSzaXQyKe6ofhUkS/OJ7Cf1eAV+uPyAumCUAZFdirP12TH7lZ99Q6VgUAWNAiv65lV9x+dqQhzJU
camDEQWvr+YwjnzC5ZXZYNVSHHLe9xmNk4upBiJFtDF5OrjUnDsKrDy+1CZ+pQFPlvqPzmAEsZzY
tH6uxIUNJRkVF2q7DXCo3ATPuamrYycY4d1KxgVS32wrh4r0r09EZfZkuOKpttZw1zNS4Qy4FIcz
9l1gHrpPq+y76r7J9WffKkKMtMyQGMIEhFZssZoGCZZ1rPheFVlWHKbvNRBapyY/YFgkqXvTLGlq
xxaXuP8zOELSmuGWjkHHTCe5H3swpQ5RimSsl+MF0UZdTC/hbqWAK/ZSZz2hFj1C3gzoBYVzbmx6
cPl3/SAeEMs1iypj37mkW8wdMfwxsKs6Epsx1QvDpQZGQzp2TIFIugKqFyXOVP5f1cOpcLusq7q/
2E32to7sxswQww+FjdnDD/x8tkYrAyyP4VH0wjJiGynEpT4WNC9wt2BL1UPuY3QZXfnptE4dtmrh
P5ul66LkAu56btsrAbkAsEKgZ0iSy10pbLUyg3RUBQX9YADmFqRUsMwFPV2lYMz+EIEG7klmnSdM
P70U0LCFXFhcCJtklyl2xNCLUpKNMzNGSqiHymw/pkHzqM2Ls17tisdGCY4YB1scpmdkrv5TDkh/
j0U9n+X2M6slZsic9iphHAwIMpr9VE91Hvaormsp8QMpZb2MnVJWH5wkVmHTip4gYmX3Dmmj1i+d
r71DCta5g4d+r8+NIOZz+Wbm55aMYPe5isysz/yshnz7vjH1hLTwLjneBj3rzN+BMJOsb+VNHuJB
En3hGIz2NX5N5QJX2xz42kIjZNeVJQ8316qO50jwhU+nTk1sWytO5cqXJzZ28bbx2SlzbmsIOLyi
mDXeuQUSn1P0wxsgOe+IvVG6ZumnVl3a3Sj9cSUpW+chACYUWsrCnyXUl1laIb1G+glbRRYJJJA3
FssCamDqDDol7P/0P8oUhHsUCbaLfYxp4yGzHisSlKo0eQRRrndqN71wDsDiuH2RIJzyZjQ2xCcl
qL+59wxrHTE4iuQgqEMrnDrexEEIE5qJLuv8/nz1z2RTFe+etorMFyK5D1vE5R4TrBpUOow8mRKX
nbpbH2FMijmFlPTVIr8IjiioDadrtDCEn/h8JK3ty5/TpjzTvENKiw9GuUDadxR+FM25LPDT3bYm
jNsjaAuYG54aa/L0h5De/DBjobKfT/JzQW2R2vA0YniE5QYsyb1iPQ1zwcjgOdmA3Kn6B+uoqzaK
fAqvhkQVQGN3Qp7DswDpZx9zkr3a8QIMHgK7nDtQnHV6k+U6f6X8D1psAGDBPk0nFn5GRSZY3NIx
JLknyTeRYko0ziPUIyEgVH7ZZdZfhAU+3Y2mpxnfRUHuCKgj1PWczFuQ5q7W5dp3ZvWVH6ZUoIT7
llFURV5om1g36INJI2seiYEq05IFtHDdiQzaHHwRTGUPr1cq51Zkg+W2cd96FX5Disg3+ZnwVIDX
SIMw/k9dKMiGjTJTWzzIiJFIDJbbhdu4uugyYCbh680H1VUCSrPVIrYBUANN1NUdYLOm2NaO7BKK
Be4LUVrIqWppYkA8AQ0fHdD0n8vukckKPJx1ei6KYUrfMYHHWbiWJmqyke5pwbLcJzpMa1qtFML9
ecTBpo1i9+xilTJZXMugRjlYqo+P5mapeT/lZw0VIFn+QkfdiHPkzmsoXDrSSnGdvCW2Hy2Qdk6I
4L4cNzCM0YtDtM0oQD0RVZMhoOZtOMoauW64bdxYXF3mgiA0vF8UhwOjbhFazwsmPI3F1JG4D3vT
qmqlMdk+yBQVxwbOpgYdUrlKeDhCrhdPJNy3HUg28XgBHKMdYgSpqWmzK5c38yChWU6Z5IXr+UVF
Y+6wuwfc7HCp+BVCG57D1PinjkYJReZcUMT2s1q1HqE05EQdGAKAtViGl9PDuIjDtlC5sGV1GTpF
NDj5v6jrJQX/o9jtr96+M6y0Cxx+xCoWrVWUo3lXke4mK4g6v3oxQkQR5Afbhv4DSrW4+xtwIDnr
9yXo97wLK0nkNh6SI8pIFSHCFbT+bcropbuMEozHsoNCTzaK/ic3ZMLsD1K96fEgwHmxfnhcJy1C
dnb/A6MjX3PAomG8Ve/+vV4ZEWOoAHKVKuHyv6uucsCEEquN1xWVYAHn6DyKaz/0+3hQpt0LlPnE
vf8NQswbKY7ZExV/wL2ruCXJ9zY3IAUYPaV09uYVx+PSA1SqL3PFfv7Ip9N/dCx9flqonSeHBxZ+
aiPRUWhc8b0AsRZqzeo1twO/EbQe9NIvcK7IgpNzrXv5slIYEorRpc/3WC5cZGnS3U3Ezd4tEkQp
A/+haFbQpseEIcQdyW2jxK8ElToAct3NO9gBg2kjcooOMMPXMRw1uH4YejdXCyZ78wqfLvNcZPcz
q+d8HteOg7yXsQMI7guln5My2zfLCC7V09CAXtGALPGlKwxY6erOMMVP1PC8nN3PZ+8gZG4rFArU
Pn+C32Z/VdPDiS/SYhguCAJ2J108AphTyjwhEuTtwr3kLkEW6k2WHx0G+ppUVSYH27GKnZ4DYrk3
X7XHyxABKjX9cAaMyGcJ7vnif9cNYCcjXeKDafAlw93+yvWhpN0RClOGiqPWeRTMFDr7kk+14cTG
PXmhH71zOzH+rHEX6Fohbp8k7KQqMml2FzhZc5DMpeCdB5JXaKLoDdVTjLw5A4ZdW7xg84uXZmJr
40p4JlsezNt7JUfxRBnPhwPBq71Mx9NLmnotrx80VjoO0WPLLkSVQjzmSiCyQvl66b0dPL2dw8Uh
7BIsr6JYbe4pUN8OxD/KXyv6hh7PUcaKn1qlLbpwzR4XJVsRn+nLRPLZ3N4Tkk0vdTC4UpOGmJDb
+zUy76ANjwptKT/ykrs0sI8OHMOl2ZYpKZxiVzLNeUMq5DCUZ2dY+QdX6b6Y22xpzNneYs7PehxJ
ZhbtGxH6OBBGSfIPcZ3dW//PK53WAbfnFp4rAid2gSywDdJTLq8V9R0XVtI/vMoZUCa75ea9BhT5
1/Qxiew83Lkh3t1HvdEt4bflWRSrki9uw94ACjzPegNaK2qQzMjasQZ+axB5sUWdBLhs8XGO3Ebh
C0SsreATnn5vNxIlmOP7ir5Ml6+gaOQs6HML0+BwL5eqNcpbbqhPF7I2vRRv4PVSP6Sc6njoD7XI
MUjgu6Jnvzrd4DNTB4nuZJZspFt/PWkkG5BGXrxcs9HR1sYcbuCuS6Nz808wspOGQKBK7OJgr+9X
bS21hgw3Ne7cH0DAI2D3eO2M4RR0etdvChTdEogrPDe7bnjRMIbO/WCnSVM7e8lMoxOPeZRMp5iT
RT9Z/Jr1M/FVQFPFVC2tnefy+BUXAUKsv+3kvfwDs6cBPFv2tfDzGAdAc7sfmrOCIGPHDxg4nIFV
1m5drf9NXtIp4SJNFygoHsnaF3gneWzWSlTKn60kSA13nm3/joY2dAIAjP1+yoLxTu78wDa1pFsw
b8z+iWnww7XBj3mt8bFo8gZkkkxN8bSDHVgIVqG2YGWzEqkPEPg9oDtcmDLmIkDA8KORffm4lXKz
HLztDub6w6uRZ6P0SRihy7zP0ywaSRcVq7/z43gSwo/+WoG+mwtQexp+OVIM9Po6KLRzoBgUnJbE
u64uj2Qux1MigR0amM+DDhF0SirwlHs5HNPjbAN7XbwytH1GPTux5+l7iuhgJfjlmQhq+8GWKVfU
T5In1aM/BoqU7zn8JXXei/htmFiGWvf91hdjyMCYXgEXpKsKUqNhxNwopzL6nSkqoHQtx/urWNkz
f5Tm95u9nGl3AZYQtAsrJL5jtI4JQazqWDezK63OwO/Hq7on4ynHwvAPlsdOBpEXo1U2BBC8J+QB
l3euwmMZSQHc6Y1ThwA3ewpYpu/p4tkNtWJhte4WohImpDes+ts6Y9nZy0TTOlGxb2FbBI2g6wa2
7XtHYNTQy5UqM/0iIMx8E5dLQIxsrzy8xPxgrOwUoG7hFTktS/wjnBICrRbVOhTwNX1l6N9TepB5
Y+Y9qyGvaL4/OlZAinYpust1VH5m+nUW2ukIWJC7hFSNBdEXJ6uMveQ8Zkgp5a6WlZgoFYXJH7U4
4JaQWODhxF/l/Tog3RZT/NcHGfg7HChHwC4QfkY+d/aWFySta1xvY+BK4TnDRN3UhXG2XY8RS7+/
ZOqK8LhTbko9rZhZFrijfzUquEBdc8qlmKTgSCwVjcEXBQeuZ+cvani7k5dquP2hhfgMk0zTbgI6
RctA/AaBUkfR2R6jnpQJFEvWXW7Fvo4ei8P57LpmEHv4vzaopXU1foHtEGFpkzzioNzcKBPW+ydx
WJawcB5Ueg/Bv2MdE9ojOLPE19JBF8CjObhQi/zFdCtj22mhbLnBSYTnOJJ4l+Liv4b4fH60eDTB
TffLvK3agEtsRCxt+x3aeLtAW47CG/jS7ua1hXZq44C5KJf6cQDaR06oUwuhBP7br6DtZTIyTJr5
miy0AAc5ediuUDdLAFt2ZE7kohgkUUEj4VDojDEhrd45UKbAbED9cqbdpQNuQ89XLgWly7fO0UQF
vQom5bhMZ1yvVGNfzdxQkBs23D9RjzCLcvrn2twBbDxBau3bYg+Dygba8Yock6ZpyLXMioLKeP9O
Is+3KPn9aLiQmmJPW8CHjPAw4no4AjCl6UAF4Z8snBiqKEDzG/BpNnI9ohiFBuiwn8ZaTQNGA4gX
5Sq4wfCd6gvD7uSUGjbayoUQn6nYu3nn7UV+jCZK+tNqj7wInM2YK+eo9s11GD4I23pUkf5icRv1
GeL3nmHaiXdP6WI5uI602soDvtDuAGzMgAMbBQMNAVRNe5ckR1NPN6Hsn/v7bdJ3sNj2P+j21MhF
vQTYyKRnwzPoLV8ZfVDLwUfiUhhlLoJ3m0PJzW2GINVNi26vnmxkzboGC9PY/ajtS/Mw/0gF01tJ
UrTr29UAPSrF4P2lw6jwOOnbMpIt0xVBjt3sFhycx+bgc8yKHsXrzpzvvo1960e5dAUkacqnus1Y
nxkO+vlzjwyckwGYdYwWgIusoy8lPpkLIVAzHf+rMV8sE9CikiMNAywt/cib6FRF2Xi5fKDG6BPe
Rf/D/bLVHN2xqgAtFsuXyvSOSGrhzMn7IVCyekr8+Ftwgok6VEnaqJP1/YEvASKhsQsUQxzEL/IP
TYsRXQuqJwGpUvEedBaiH7/60GCOPhe6V/1ONXlN1GFrykHzAidfDJ4t0OlXDM2mYq5MQCt3I9HQ
t9dEcKeZpgnkqztSdI7zCvZ5FOlt99ElRBn9I1qqjuXeerEo0stfCvtCDJcAtdw5CjsYpr4yVNU2
jyd5hCu4dyGS34LNv/EorBjKVvZ1H6Nnw5NUZQcxoPdSkJq+lqRr3b8LrYK99TTNPVDABqNfFShc
6uF7yQoSBqiRaruaf0ISD2aArRXBsUPqL1fEdNgXpJxHEf+HK/dJUDwikPvDJAqNFXZcLzaHIdlV
75JngBTqjKLK1iE6CV7nY5Pbq7GfJAtmJWYh7JsjS8Wk4yjeaq3Stzw4GA5duHfRbt9xhAmXRdjA
LNsxHRDE+F5IqXTtYR911aOcd/wUmKLZxiNVv0JytMJS2U9tgDPykN0s9syo2OAEWLNMBrW010rj
bgig19Tczi9gd8kcW+sgQhAd/lbMwSplTIJiSlYiuNL3ZwzigXuz6b6hBbx8Drdkkqu6nCejCB1g
x1cPpnuAJmFcQkuI0pcb/ADbskAYSFmH3vkQscUQkTfiT/Pffit5+pgt/xNdh87nFqemSLWfKuWt
5QW4N5mO5WtVnRT6eonhkcyOh3unp6OSuUBg5ALao731rPS2aYA8C0Tw+aJDG9FZK6xrHmLllBUN
SpQ/oiFi1iMX6hwrtzPMQEfuhRP4XtDhtTOpF7Q12YgJgo0WdpYJqyq7mL6thQIT8fTAFVzxH2fE
9sxA0kg3jrDPnz7MRn22N0+iY9XqTWuiVmCC22Jq5LfHv54RpJlFnk+aDcd4uIeew5cyTkPryGCa
qP4LBjMh+4WIE/v650ifg+gbUAYC0SUVNvYySlIsqjUcu+cF7kIArf2R03abkPs7DKmXAaoXMhTI
8qltiw4Fza4qSemal5nSIkJXpt2XUZHzN0u/2SPvckjOI/5IgAHnHH0C4XyhpLdiB0tmMDxhyxSg
sarwuE5iLvBQPK8KzxK2PYbVTvCV+PgfO7sqqHjO8twX5GYVjPZthRD6eVUdd5Bf0uVduI1k/qiv
9ybTE+JVB9ITmoUD34s5i9ltyK/1uNTNni53c4zey//im0eFJzrCbUG813kz4Lv0d3XMGFGZ/kyy
Sel5iLvRE0U0y4Uph2+CdKentCniMX7NMBCVzuIKeLiryo5c7y/3GTreijI/N4gWndoSu+oZMOsD
RHHSYkFhm115idoY+2R/AUYhOfjMtCVx+S2NPdC9WdsoXX/I2vL2m30aRu66zLrCDIbi2ubN50ef
TNT8rHjGkOPaiGwu4SN/9DUVDZXpZDS9LnkPB203T1DivuDfu+Wd3dPBLF4tzBJl1ojFGmM9ifc/
ojPvy7uIgtU2WCUQWCcs7WCMJK6Vs5n2Dn0eV+q0EOyrMCpcbFCIUezVwuClwJa3cGYZ5zF3+8u7
vmRXD1/y0r0OiaGquSBN5PO4D2AWyiFRHgnKxUg3CT6lDBXwmMiqqgDnLMffx27iE59rvr8eEUg2
El2Ufmieq+hOk04IzLAtPcVEsQICGV/G2QTGewBkkXB7jHoU8nbormY/DOP9/0a/R7GhjpOlppvf
gCaG8WThXIyuKve5Jm1ca2DTrqjJgUyG0qJ1AMLOlyZ4Odprb+zpvZZBLPtFZG7YrG1NzbadGOr+
As5GiqyU1TsqxR/AuwnIFsetll/UIJzv9+AVZjjPrad16uZgC1IBRmrAh6eeJB0LaN9UKH0uI+4k
Ix2wxUEEXUTc8VjKYrBMSePdZj+aLEUb/bLXZ43XRw+At10Y+lJKCF9m+X1pUDptKwVJaj/Zv8jR
LKgG9ne2JoicnYvcu93DkgcWGAe8Rgid3zzwDk9RBpmGXGg8w2DrKCsb1mPk6cfkCdLZTPXZxp3N
9FlPo5T3ahUx8uJHS5UVH81OSPgdYgeQp/NAgvHC8+McnU9lO5l09N9Q3sdRsKPUL9uaNgSVigKT
9vey2BKnSPtiI7at0TicS0yLvWvAoJQemoTPEmggUjKSD2t+1cBsUSzVXosQxeRGhF4rSzchi9ZG
2zHBUMGQ+uNKTSorAP66uOv8tLJh/A421OEcaju7JsZI2NI1WexSZCKwEbQwQln4Cg5LxEOFeq1i
8yU8d2+r58UvamEkXOy4FxJUylQpUu+xWlFUKbqUSaDbv8lmTIaljUZ6a7iH0uZCF19lxdHMXhRO
wqL7XyuIzCye1FynhBjm8b5lsk0melzmJp6BHzF3r7tcYLAcZZEv7hcgVvg6Zm2UKaxW5dJ4mIYH
0UCBJUjuFSoqeTgsxrAHxA4WNxbesqyLu07+rJdq+ice1xnejRbDGZuiJ36S1W07v3s/gO7LjPZN
DT+8PcUPIs+TnHUbNHZHqLAc+to1a0HTI6bMAEOazj824ea+hc4Mt94KREdKolqxNUTQa7VSqvAC
o6e0MYnWtg18tAw2/p5ka3LmplAs/tRgXVLNb9NwCv0AEnqUwhQWwDX3zwKTNDr0p/l1H7CMniZZ
nrkIRqcmUXn8O5YphqupHnc/IrTPBQhq4dXvR+QXudAQzbOOuWa/kwMXlUeokDUZw3KLA1zxshW5
QPWZ3QAcZAHXk8ApaDZW4OTZlOXxn2ZUt02d9fvn7kSGI6DU288yiVmh7oIB7w2fVLGqbjDCZ0hQ
lzVZBpfu3BDCSxhEYCOoUyQJlNQFNeNvFcDL+vmKfGSVbH/RRIBpNn+02x27TqCKUGJ8wvxNKjRm
UGFjCUsPy63qb8Tn2407k+7/Im1Ug9qhkpsA80pO0bmiKV3yPoRwaaAq6+1IWZ0T5i713vs7fx10
A+k2dT6Wr9ysKC+aAev/Zrfrdyg5f3MR7w73jYiml4B60uf+9d3JbyyqcxH3g6a8nNoIQnFNmFsY
cKScwBaedSZSWaFRW0x5NGpkWOV3+rjWvfZGA/1ktO+g3YYWepz3i9q/KCpMYZR49G0EVfq9hfQK
sGodeQ2I3IG/l/xvXhLrK++H/RD6djiWvIen1ZoqfYu6nWnSg7H1TlbN1l5C6YQuoUSBpu0Xwtk/
kLFSQ1d8NiHMZEvEsJk/m/ksOUwlTarb5IB5fuQ4dKvvNQkNwV/vOW/htbbKujMdVdkGFigmYRYh
iCD1K+hAXFneiq6rPj72Jfo++MMOkr38YsuQkqh/+HFIQB3MrgZj218mYWhXgyVUEw/pp0oi6+FG
D29kevuIzelETYvRXkemOn37Y54Tai4twGc2Pbc8Tqw3nj3SWqX+V1MY+emKHpmvjKn6qq3o0MC9
xYw3Aw0tKNaLU3kEiZFZOzQp8HEv1kpPU76OM118nw21KmtDRIcJjjpAs3itMMnFR1YrBG8vkQZm
081SdO6tzudrVzoQ97WKhvSd7RjTxgPjAc7U7H/nUZ+KKQoHnAYSXGq7au7xVBpZmeKZgLAZsVtG
xOxq2/hoFLVCKX6ayhZohrEYK/2gFAxr0BJt3iA7bWfx+JyJl0pnuTOMydtUWsA+3fZl5NZm2r9C
aHGaslZIYIOKQXclQoFRXXptPmqFGfcT6QpHrTONA4xfsv3b4XU5cLAFz4xF3JBEYobED4E+od/p
TkbVyimZXdDXdF8/KixhVsu/qj7Ih7SYLZQULF2kCCnFaocVVqHyC+O2lHY5eKbBp8aTcNcLu9mr
UC8awAC20npo8feFsXxsXqTjUsoGURFX7IZcmnJYv7frVyqY+yO7Hxz61nOjzBkhpw/54VV0IuW5
QHERK21zYui1fxMJKYemaR6tcCTz0XhhR+DVil+G1vy07uYg3gDkCBFDHWQTE2vFoUTETC+YN/QT
fNkM22seBpVQihuST4QNT+m8NseFFoHCMCUk6fz/XgzQGrsk/ZTnJ6fIY5cNsHZKMq3LVJ7/lhFC
7BgrC4J4hVqnOMZ2aVSjN+xeSYxvF9DIPAj0TqcKhP+R3Z4Yig90dFYNIA1tc5is6tEkJr7rG65I
4TZaOhggideoE7Jp1f+wwn+EL9TdzbF2txWY0bYggxXUO2nj3II+9TSdyCxOZPZeie3Xxld8iKCD
lRPlXVeU4HgMm+5j47RUZZ+GWoCOLYXFE3jZE6XCTQBmWtCiSTHe3x+9cKa4ODv6Vxqyu3t275wO
9OMuPwYOtgib8b9Gj3+sp1KzfuO82TUiKwRR4Srtcn/+NqpcfFvNOpEclChH0xzrVrHhC9nVUcML
o49KHlybKQl5gOIeNpxNsx2CKsZmBfIKrvKrP8zLcDIPnQda32znuOeYocsa+I3hgsVbxEfsMnZe
iFW+thBhLiI3yVtmj4t27jdGy5U9PkqY99wMfrqg5W6ILJHJXULZV0KbD3KO5VsddIC9az+dMOwC
rsexbWnmZf/CDptcPwBjlp97yGo1L5KfWNic3tNz7Z9Zcx1zcifURUKIE4BKwTjSvDUp8hQq/Qyc
4+ZeLX/zdDaVQ35COVGxyZshHC8ozFoLCgFZWWPiqODzqHxzdYLLyXoWTZEoWOPV3MBThxOD5Dp2
qto/jJNbh8ShDLrY90QrwyXcaCEP4kUpa2YsgzycBLo+3saYT8hF9gMTW1izBK/gl/qSYyWa8JXq
2avTwllPoKp8NuUpF8JX6hm3VqhQ83cdo6SGOENVquF76LiMPja6EoU9Pe4FJvAgsBiWJe1DsPDU
rVMxJhXw/FWhoOZu1avIqyv0H1+3HoXiuKAdp8CvyY3kV5XieH7th9tTc04erHJLPNHA1gjw20je
VdJCSvQZadc7dLr2uBY6gqiXHX1UjhBpYnAWyy7qrpBzQF5WyaVGLtWyq2t6xkPDh0MIcL7KLMEc
2XK95IEuz0as+ZqQfKSWsr1Ghcas/tPfjiOVfNxI7cOs8Jx51WvmLG2shW4fpiZLHpKwLKHTzNMA
zJTu6BL7vAAAZnZBdf2SDAfNrC5QWZIYPsUqKR2t1iWxzU3UcEDoOvEwoQNevvH/eOUUKWipj1qT
BPnyvsw0Rc3olGnqJONs2CsuXqlkaEG3zZIplZZSzd+2WFKSMyouN7ILao+Ui9ZkXImZbSt1sD43
PQWOADkB6aO+VM6dt9oEsungb1iOuRn7df2dDksZfJ6zLcana/rQU0bzZEKXi6b/cbPQNFJ0eYHW
CFmuFyGRwT+PuGhq8UdjSPcy4Y9mpOrzVbydeG8Rp0hco8F/pqAYFfx0F3sKybaq3olrZ0auaCvU
l/PYW2wL7sq8tIkurrgWiBw5nQq+gunUhOifEFMDZR5msUCgvLEWdM6Zhv85vvMjTzEW17J2T5ru
bX51f/U3efrW8bFiIhydm3pBTij+kal3jzD9kJ1vQvv3MiOIZFEKu56GCK8xOLYd6ZhuexutV7nL
+nKT76slewe2MYQkvH5rhm222+Md7YVAnVDGxQdRIQlW5QWUAzOeadUHCtt6mK82u8KYJQ94pItW
SzXzssEf+ov1ISSuXZJgZZ/UsnY3MI0XK3kheoyewW2U9o3m7J1lrZ+nHlbTi56COq/m4USAfGQM
pC6De35lXaVztoCJrfx1me0DPbFe8spHA8u96yLbWPNbK/v7d/q8r2OTf8RiWvvV9fyHFGs210R6
Mda5c7GhdnFY6SM1jEA3rH+AtBhrN8BLeSkqedNt0Ue3lTfF6Ck+7/jvc/Bf+D9zBKRQz6E8OCqz
k4yfcSOlPTdwaDEdvL/s5MPhN3tWO2XdCdftsgwqjouSSzEx5s+w8Os2jpfu7mdz8GSHmXQIWh8T
kAsaXsgedUs/5Syqk+LVIbyTytu+LS7E2LSt1BOW9thF7698Dr+sDiGc0OkYR+sA5/5oAnyoezXp
xteJFY6qAhErEXkGjmw/Me1f+/KHdbDfryPT0RoUK/rTvyXj/2ubyVwy1fVnUI9DBAY1QzlfQT8U
5rsT4vG8KNbOF4PRKu1LtzW7O10TAHgQcbqu8RLF/AQdp9bnb6ZnGVkiGeYU8KVUDYCouicSRHZ6
rXXjknW99WXiG+Oropj/LuEYszU2wm1NPzNK8+qtaKd5LM0plk9aC7gORHEaMiocnhNrUd8G/mRG
j7aV7sWYtztN8NNnEKXNYGr+9/jAJWBI5dcrQQ0jcLriKDapbks+Kj3sAw/kNeKPMCafDEDDZzrN
o7ecxthw8EBg1Y1EqmaQLFIIv2v8TvyMIsoRogM7Y1eRIzvmHqL5Uw0EC52cncdwj1SZiwfnXfrL
pST+m1TKgvJQPwyzBBUBSJj+RZ7PoC+c3yE1JsNsNcxg4sGnF6isHkyoq9cChR1LIbJlG6I3YK+K
XhZKGbngWEI3F7oC7AgTxyxaDj8ex+ltpO5/eX7825QFYc48mHF7hpImIaWC8X6sFyHPpPXKnMwt
SbW4EXMbhjlHvxSed3ezef/Hx8W+SaVS0MvMOg8m7EChsT88stIjT1Xr6Hhjgau62QasTEXxhffY
Mj2uh/KQUmUv+atOeKVn3i4H8FZ+swmPM5ipF1LYhuR2Yp8/njTP8gfRCjNC5SSKXQg51Ah1pTy3
RMbJXNdRz/cgvSbNz3drazYZ9uoIBexZ0YkfZECqWlmE2mEiGCPytS4Osetbz2EpiTGh0ocpTNLG
OrvBFCZKZK+Uv+Y/TvW1luBW7ytjzApTeNngzWNWykXFIHBEHL6gfAijUVr81DfrRtICFeG9Shvy
Ja7AkwqqDilomv1Jb6ReLKvYCXrKufqYPQ/ftifOkwiE3s3IHwr87Nf1HF+jT0IGeup4nmHO+nY0
6BGMQo5qQOpwrzFgvbCWQkDIeEU5FE9yFY40z+xEj0OKVcUr6VB9h6JfjOHLm5yMgzpAyEkt3Xh3
hwB8F/HEStoPDs/qzkf61LoGdmuYf2QTke/CeC7aN8IEm/+p7K9K8ekozuY4Fh+xnxRi0ymWc+jp
N9EsmrMikDQrASXUR5Ay5lsDFq9DFGjGtrwDC7JKrPVgMEt3IaPWrXI5TGf5SoJKjSEUDevl76w6
Ic1+oFFNC5oBMpBrUr550Lg2R+xhiVK+tWBRtYhEMQ/KEr49ARZ6rrunII2PiHYk6q2rDzlS/Ngh
54yTuYCULPxZqZ695NYcb5CIfyNzDd5Stpwhi3/yvM4v2ECoKQbf/cx20xocLNgHMczCv/7cj/qU
sGfNXmejLF5ku3hPwUIOEdF3ZMhM6kCQMnokRpG0FgQ9hoRMXi6t5Ry4uaiXMe4sMFqKzI7XFEnT
L+nkjtIEsB4G09/gYuvElhnwR6x1q3T7lU1lnZKUzoiz9FKU/8yD4URPFJxJk8ctXQJkgsYHCgmW
wSUNgIU5L+eh4gj3Q+1HIlYXcX/9+VHBjRjN3qOkc7eivudYS5HdxRnLrP9PBnotGc+tmzoUsrVK
waUs8VlwxMr6cz3XZRhpB8sWBlP4EYXXPnfBY12VmWgWraucQfAdtDjvoOzcW/7Vyjc/XW9CnHdC
rUYn9iVLZa9lJrp5O11Xh1jbLbVKHcYD8wBIjcO0tNZOPPdOwDiw+RW2F1ZswoG7DrXZhrTvfLk/
v7Dfgd+U5gu/OaBFAq0njal4cfcq+gukYWkvViIBA1PRoRsI1oEiddhVhV+MCY5PhVF61R9SIjz9
pSaud4rLSPq9PRVenrL74bIBOk0FfpMKg8T3mR7xFtkejb7Y5sueRLRKFRchmQ6padBgvOUQINhb
DYKmbLeZoHKtmmmAcxx8FK/MwulP5mEz3rwrbgXD3tycy+d5L2nPJSB2ZiU52FqhR6jvwbPKY2Ln
FaVH4rSh2bhP16wv0eUK+0ZgQs6yv1wpptL/cAiHne52VAtj1V0ZT9mRLhXhmNFtKFB6Cg0G+xYQ
FEkqpDjh90ZwO6nmfMwZ3/EYqH4zDbPdAFwDcVwBO9e3ARwqQJR5Eq0N/nDaSKbbdAHvwYvIY22+
uRVf9M993m1RA8TN+lwmNwWsWHGYQroknepRceH6beo31PmEgJUaP42aXUYAHhPx/bY7hg+/G5MN
2ef/JnXU0diBTOPcvYBKQkzfu1CONk14PcQygfgQJ0rbqk2zNS/Q93L3Q+E3H/QHTeuK7DidetPX
nsKyQbD6MljmV+CndM7xdFqZ9W/AFd39tOoUZCWSD9lv0u0YUuoW/0bfXrZi/4h9OKMkdcCV80eI
WSP16M21kYqDnLVUp7GCFdxPFOzK9xy4bfSViQfGles8ReiBrvewpgUJ0K92XpsbwgURSoE+Fq3G
XMpOaZMPTv1kgh2nQKTsqPvz8WiTZz5L0rnucL1R0aMldG+IF5IAg5dZaoRZSowkVLdLox2JwNee
S4zsYR0N7q/8SpnnBANDY70Wi3rdiO9Pytnl9VMVbzYzuyO+Aj0GgAsN+55/EaN2n+uTdYIGe5Sn
+sw0oacGAYc2cuJ1pSkCw4D5iI20jYOnO7KU9/x5GM1Og+fppQgy4Vp1P6+EEvWsatXgbfObLves
uJiTxQYyK/j4WMuDLLdq6wFqrjvSDMqWzQYQy+29cv8WugpeuzfFFN+/EY3D89Lay89J/Anf/pn6
eiLnZU42AYaWavueVXtq70la5NvIC7Qb4Yo2tcdj8jcUZVFDyPpsz8mUrsomVaPj0eUgqtKts5KZ
XNudxFb8j4XBtmDMrLOlY3IWUlR/Lg1TKKmyUjgATox6ehDkoLHoOd7WbCmdpf8iM777uSZN4nBY
XmTI/+yu20ajrxTc7HA3le3CEfkCGhF1NnW8Zwt39Fk8JqaY2mgQv0I6+MQsVTpS0I4XeSDDzGdL
Wj/b9Nt33IDmBJeU4jNNbYAKapIvz1adav6Yrh28IwgHJwG1OIgiA78bfSgi5HgGNK4NTWOpEL5O
pNPxd+eYscSHeMRtCe2Q+cuTUeAbOVyxJ6DfLJrT+lt1DjKJa1vrAhaPLwHUrdjcd7inrmbaOYIe
hsgd4st7Akt2hd+R1KmiqvkHsOo59EC+CxSuEF2Q60mxSDqfcGzFWroVeFUVfRJcNa9g+hP0vfgh
X1OahB7aMmZ4ITEfOvMrxAbySh/zS1p4hfayTX9bMnNtHX4PGQo6yiPyNsYKz4WO/E7NDuR753MU
KJmSUn1eh7EhjWSBPnwnuOOd71YH1C6E4f/EjVyZnRUOnI4ZBUOldNUOJCJslHXvNZFr8XPrgqNg
MEp26KkvKlQC5A8/ZcDTREhYMyLxTpqMuVDerkCF1bi0adE60grjmQN87tuqmBMLK+lJLKWJ4V4s
C96IeEFgcZ3WR4CN8YBVvqu8EXt3Wo73/JGYYnZc5XpuNEvFuPfCZ+aJYkgLQJPum7DW9y7whR//
66aREwPskQdU6RIpKgAhoUg6imTNIqKNNEM+4M2tiyOz5RD09HTJ7bJJlCCli4ORPGv43i99Fd5i
VVj60VYkJeo3G7/NTDFnnGlOHSdd1D4o/jEqC1Ux8HtqLWbkIN4Uq+B+l1M7jjMvBubKw493nSeD
RtX1lqnyF5BGkmCwr0uwxR9md7DpiWPXAgpnzxwRSBz8YQSVqZ1kdNhGeY7no8mgtIqxm1M/0lc6
ZpRKMY/atxr5MAtlUCZwLJ8mcONTxM0bnZ/YnVYrRanUSZz1xYBavLTQKmFE6cz9sxHdayJAc8nY
Drxn/TGOn5Fu9EMu/7Orm/KZtcyCPAEJDIjeDeWbNvvOimMa6V9bU0lPErvQW6L8+/y41BerSXJ2
aZ8I+FfJJjigZQ7I3DjOo6d6R42Gw8XAHTbIenUVqkEMy3Bh9KWuNyUbMOvFI+oZn/pzBCIj97l6
luAWd1tphYNmLYd/nvVEKY83UKlKZSUKVx3BvcTE9ihDENiHHnAhUl/PtVpN9C5nELM3aTEm+CXZ
SDWhqcq0JTptMp0xdKLkb5l8/W4czpZhKJ2Q8ONIvqYiZa8QfdpkYj+O18wl4jHsoqZNzYeZwIk0
e+BXM/aVls+lW6yXY6iWmPm7LXPpEq0U7Y/U1DAOKypWPwGq1iLyNBcVhx2xJ0m3kiOu0nU+8v1R
26W2sLC8i+OOkA+NLPvN+j3TFw3w2h5QHI1+ZW8WBPh7iUYzTSDNz0JpDkEA7P/dQYeXWXxk8pPB
Ox+sTXT1Ev/5colSjW1gAAEcSFUi5u4xjZl1wmkIgjbW+Mg0oJipwWh2XgRrzM2tKWlgheP3+R1N
B8bzeVk/XyT9PdCLRKtI6Cb3umoYZDSA9vUraoh5yJIuUtFxKBOdyhmgdJx++dFbM9ThRoalGLMv
Y90nvmTf9WSlXd+NcClSXU44kOfCdehgEpq2fOKzn4PHiE+HzeCg4ftuHznReM7tQzNu5Ku49asL
2C+vo9K3wqcFJhfPEVeMYQJFPhUVJBS+/13Ou52QwKB+RSch1Wnl+gjoVqju8zcZFqqkQrwSR7dY
pbvOy1xne7JekdKnD3ufv0w+WMYWO79yQ8jb0AuR0yyzDGXAZD79h02cny0BcwcHEELahfc7MgKb
oTXqoNWt/kAJJii0dUqnKfBHvr7YlazAm3j4kIxGK9sDNCV8xu+ZrPiDNbScqkCjK9OsGtKrtf2N
7hKQaG38pkkRiU7fnPpWHJ47UousuQDtvE6GA+oIKAGTDm+fDQvauGTv3pCQReuUbwjyjNSnoWaW
AECShNvgWR7aAobcXxRoenUnTI0iaGpZ0ye8XCMP4l94VeVJVsogCpLDA0A1a4Pw0rxoUYNK6h13
JF81EITpXBONRVxwcGqiJD2XWgLabtMkU83e7GiI6mrtpyBpNNH3WmpxR31pmYqIz9bYV3ZKc41L
C/N1bVQueBxGdeYqlSZxa9XRlJada/xuaKEQy+6xpTzhMmmu3+tITQdIGCQxDSw/G/W3xs/34GRP
lUqoSQwXWs2pdkybzHeHPV+ZTfbHHD+UqvmCPaA1jg+OeWHeeGquFMdOdY+WE3B3Rfa0orrVRI08
ULOgxCQXrTR5Mce4owBCQh9yPgSKjkJxquC7ikF14VZKckiKkfbO+51pSjeagQZ4tpw5M0+Eou3g
3VReLQK8qR0AGY5wJVpS+6Lqf0WILFDWHwJyInNFNYTyyFA1roPkNWjnKkXl/Cq+5bGjrxg7VbgP
0p9X+lBxduT3uiJjil/lXtkfVw6rhAb34d9E+IOrjyGvE/Ir6k9PxrkujV9b07JDYfUvHYGs7jvK
u1xZKCjBDS+0Ojwi3cpOrQ8G7MVTtKNKyeLaC/Oyy3o5K7Km9Tjh34i7ARo4MDH+oz4762EyIm8T
Bzuqfu1anqNcWSYO8WcFSpBw8W+7dN28pF48YgDo6bXak5KunkQvAAeuAJJSqtGf03epPpCy3JGk
A6NXwMNMCXrqdEkaDGPIq1rcrFIM9tFSXsLpH+XrMeHFT+Rqo2sVzYM1Pj6dZGuquNtp2FWoapnZ
GtfU8CZoi7bJfErs7BWw9ZP+Z8Ouk6DCExfTs9IR87LvwDBsnDN4SfBcf+F3qpbj0VKymG7SaeKY
mPdTFHw0I41Hg1zDjuMxNU/MTv3FXhnq+j1rkkqTDt7gAiwVlkktP+i0OhYugRIibJTZH5Y6NiKU
IGB+ZtPWr+PIUy0LcyXzAkRIcdZmm2xYHdT3+2sGUZ3xN+vwqzaJj1SPDAjD2VUqqHuu057VxcnV
o1yl0/NFtcO/HyJd+6RygpwO3PrTLcc/+nvQCgTJWFzIpkHt/jvNRX7PYDDyI/ZevMQALp2qBuTo
A0tkXFntLzMw0pIvdDB6fCBWilpiiXaBlGhVbhb+YKBkwqarkmma2rHzt85MyhzEytGYpcxCoEym
+faTZz1AOKLwmLYagQ0QrwKMII8XiXDIrfpFSLYwjWLC/b6kvvsKpFEC3vodfW3ChQd0OHQYgqHt
vH4Z8FjrtDAKf4stqlOpp3ZfQ6gMX8alW80o2lO5wmbiCzchZGniIuuNy6lj8I3sjwHBfpQkXjj3
LhBnJy2heUzA5TOBLbgVEHLoYJA5xORP7GIBHyWN6Ps3/rd/9FsEL+rZeRhgW5njDdAhYoQbPW9j
d+0OoYGv8EM5FH5iGJIzUc2J3aQqgQu9qRwuK9Ap5r0gk7kUosyM05cxbETLRCu0y4Kz6I4sfJF7
mKEjn4kVaSUV0oLgjXyv+WJNuYYTLYg/a0UIocDNGc0+DYDhhChfsZVUd+XD1tOrsmRsUDIy5f7b
9P41vSH37WgMl0YYwnvWiUnryvtVbzfSHb7lNjZcSkpq2i42jJFO3GW+i6tRMDVzcIF4Vu+XkmPJ
oyQ2Ow3r/043GGfgBXm6d2gVfSH6doGNB/DHaSXnRGIKnvLTIk5Zr1+rB3tc3LpT2POQ8wGr5oO8
aJ6CwLtA9AEi121iXTIAu1n2rWVPCU+vdkx+KhII1AL8fZ8YZ7zJJ43M5Dta2hlo4aTonn3of8YV
U6hdPAaGHeG+xvMuviWrnp5EQ22AKC7a1r0ttbEWOaeM2b0cFWA2eB2qbJ37T/NLwwRkTE7VLtTm
j/JAeaR2DgxNOPxScodYIqnyidLxwNHrrae/pAicNwC427+kRAxM/L7CsrRhgxj+GqSFKjipXEbP
JkXRcCetWeGNqGGdbyPrDuqseOlrqkYvSyZ295s6uZDBH3ok90aNGKYMQSRdrI51gWIDM5s/L/yA
I9VKbPKRaodYksNiX29z69OOR+IcjzFL7gzosvtfEpDXXE/21ULLgCvxemOo9yM7DdROQ+rMRpG/
pCNraADQhcMKyrChtUCAPwH37httFw6XmeLHVMRTymj2afMIBKKoX1Rh2ywVejfdXLJgITQ+eHML
Qj43o+yt6U6rCsuoQfW+FNMZ0b+OxFZrra1qtgBhrL089vhWHL9aJHQg0gUUXM8OUqPOsymhOyZn
Irn9TUgxQHxPPuC+3ur8K0sZKb/vYXuV+nOFtKq+v2ZiAZ+k1SZOwIp+HokXiD15w9zqymU+LDKm
jo9l3XES4/SC8+SZg/xQg1+N7AARvod3K/KcWxWbNXf+fn4Myu6UsR2fRcs70YmSoPRQWMFI/GLC
WwBsKrfSI2Yw1BKLfY02EFy80lIBG2nqzdSIvBNlAn+zsECMSMVLVN0kS6qOvNP1CC/KIyIUdPkE
tBBCL779UHaGFjnrsHQq2rzWfpO9qMa7FErKu4+e3aUQy4pQzfZNWY3xUqzWUnT5Q6JPqiP7g8lG
/eWqVr82f0Qm/hAP554VxCwV+c0pSvTK03hqs8Tu+mqyeOGeXDnFqE9jGBOZtZxRlqXhfOHKTjX+
YtX30Mdm3ImCvB/o0OWF8iuP10ReiUwhmRE1xWcOYDC58J6O4/ULSMEtY3NDZAlXhzF0b7xmxmpb
xDwyyGHySEBdQ1x/rxq4nkkw7Mym0ZLjV2jb7t5Qw5xKsZQ8Bx5UhVcLV8Vy+1lwa1q4dwNf1Al1
l5e+cm/o/jz4r7LqPhxhgQabbq/kVW+k6mnFh2vlh1eXya+5y86f7XVHvM0F8C7TnlsyZvdNiOUC
XIpQzjRM9bokzWmUs9LzxzHVgcHJ6X55Hu96TLoiaizE/ehBjRomqZoXjL9JvkUBaIgyuz3eleNP
/1ntozLxKiqXpkb8n6PcCWTq32w75SE+vcF0zAROFbI1Sp8sfcEKwB2xvmMqHmXC7LAZicFEOXbX
1qRVZ6Lp95swHKdn7kDFrDMhSY7g/lbaMxki5m0v5ImxIFPxFKMXOjBmm5ik+PUenSQBNFdglEd2
HLuonrfXjOZ8bwrKaGlCgc48lVb7CpldGyxqL4mAzE/6sQ0tG3/CVwLu9mSIkMmSpqdpX95NWBdl
VEJjSLIyx/RGrfHtZ7wV0Zv5ZnTRaIHVpcB0Z5cpglz8N9fGRgIERr6ZDkLgcrKZXCNpIBOLOJrp
qgnFUPK803VKMKhhbAMvZcgSxRaXt65hMn7TlEDIUY1CsBE2x89iThLdgT/tV5oo/kqjbI3foHLE
9L5TFx3gOt4kzSdc5plZfnKgICzuHN6TZNl/vsbcE1dAo7A+cE7GP2JxVK2eN4S0njpYdegskC6i
fnp9LLHTiEiLQjiFCIan+4ctObcfVl/GX0J8g01aEpCdZvc7OD8lrvP1JdnZ9vrUPVyea51Z8a9a
Os871vid7wlN5q7/pIiwbcCH96+SqppgeVASvp92+UqLz7nZFYCiUCDP47X31pH5QbIk9+lyz2Os
MglV+/hcQMqvq5O11D6kol0f45RY9i0BtzWuTQyD7dnjg68Uk31i56qgAe4iMuVe6F08YDYs2hTw
J365UjTbd8wcnTrFIQEZb0PEyQwouvFovhBJWQUycRsKizCVgo2WHneFHWifHO7bCCV37T1CB6lu
l3b9UscCFZa78/9RvjdX1FY2rFZzOahDcW5uddxAOV3anamKK0ryFC74XWV2mbwWf9/draRHzqoN
ICLuLaUZTBOHhlrq5XB2i0jMPrKBk/3mSHWQtiZIZxfYMtI/v59SCkmkxt7a4KEKao7fUPWRwfkH
mnnJYF8M87OnjVUVEnP+bsswVtiGv02ktdIFbUro2Uyk3hGLyEFfrKV51o6MTgmTzwYh5nN80iDj
HBpcYd3KhlAE4NeGVdaMc/p0oFPnAEb/dF8DXuIzeUscefHAyg5ZQGXIh5+xRwwY/2r9jJPCAqWX
rJb33PKkbf4ATxEeSNkDvnoLA626Vr9s+Jt2eXhk9aKH/d1zUiBOVJjS0HFL2iCenLP5YJ0nl9K9
xVo2rs8DqEF7BdllRhphBi/L9FUzcO8rK3+GJlD/pdcSeVrsV1OmSpw7kqc5NKIjMu3/0nxVMa76
ZmBWj7mz1Heu7geHQ7pwxCDQE4YNGo0dV5s4qhp1imiJvUG2VCgkNxTe0ZbcYYWuDji6mzqjx3I2
DJYAkEVLkWN6CWy9KpC4+pw1I1DmNfbxaWMTK7nNPq/wjFfaT0RFJUeNLJJnxepFbR87JjBmH1DV
m6+U/kO8WGtVLnOraE7U+BGSyN2v+CRcFCu7fhJO18ffqPln7my+HuPjwFAtnCTXus4e/Q9PVimh
JnCkD6jmvftrlrJ/mJGOcJV2TEFTgC9cM17/uCztVBaBS2UPk9yyfbsFi7FrRXZgSFj2VJ+vEyKM
aZvPze8lAoNz1oD6fIsbNE8K/jbwkrdVSqjx+XTZQv3UNrGKl+Bs/WEFzDDDSj50gavKqo+l+iwW
s+q0/bKPQHcZEHEA+VsmDidCy2XsJKqNRtdVFTQ/IwlPqaIZBufqwbFYkR2CCdFnuokUVPpUWAV2
Ln0DgHer/exPUWGwy3U3v/c8Qgp6fG5UHO10lqpUPh0XvAPerQoNBQStfV9S0WKg3op47RtEy8Bo
+4UrC0/NWwUQczdgbzesVVYUXctJRr5da19+JeD6gyQ8mAfgXHVr/VMMAjR4GmYmIPVxwwss+wu2
ZPkQfstTmlV9wICI2Gb+3CgekWpK9lOjlrFFiH2G01aEGGA7Gb8Y6zHcjlNXQvrI84m94jAC6zgV
7Yxq8am99R+rhqya0i2d/BYkmQnMhRQ2BQ6+MMLN+SRmEMjw5ZiXFdDIcqhAKwLeZPYEGlOH2r9f
YiD9ql5ntvdbg3qxQcs9xYCHA2h8ZEOJt1KzvaQy196pRdy00bgF75nE+rc9XfOfO54srAgFdsbG
HNZCzKZ/coG482E3SnV4Rz+8e7kBnke72iYP24+P7yCZF3ziej4CS6D7bqedTqeoBDSeuTx12EEM
AURkkzduIaBQg2UYyHwEs/Nu+dBaZuZFth7EeW4Qg/sWIEgwE1hMAYCRsOfrwzZ1W9XySg3Pydr2
gzklocpgES1q3Y2T5aqMj7avd4j5i2BY46oh3dcn3UNezTw40VaEUhIKjCIn/c/BLiQA9qKcGzgB
QhbRjxaPbMEckZIAs02/vNiBPM9kSrbY7OretDzvNzbnvUfGEkS5eOG/tuNUN8r8m5t2dQIi9QYI
ygC+Y5O3wPebD8DIC4WA3DuG/MvrhZtxHyEcoad932N2n5AtG/p+jNwNPtqi0iiDvGFF7h4zSEOw
lGgh8uudEf2+EBpX18aZsAdLyK1NfItEfZ4LM0JQeSFuUeDz4ZdcrWsw8D527bAGJURWbYcHiQJ5
c6hRTnOBMgnMhNfmBdaiSHEd0Eo+tUO3Tfij51epp/1Nlnlq1PHzxQFj0HNB/4Lzavi5X2u8Ea4e
wYjnMYJ/ajkYHWtl4gx0/YhIdxqBX+CDkderRAERZFslmioSpTkfozNW4VWv3zZV1Iq2HAW4Kg4W
yDNEzu1SJfgFKHKu4BmOUwaEejO3ti/gtXaeO/JTMgwgvLVhQizm/WnpNnIg6ayUZEbE4Ovwlcca
GRu6ALl1YtaiqIsCzyN/S+Ozs2qlE7wWrdiFaf2BhOnTkpuM84iFLBuSVAl0ywBCh3s2wD4p9tTj
MwJadDMHVEiFcQyegWLaHM8gE++ZAzEqkB25ltxYsZWww0abH750SlutEXAavBmGXbr3JXFRp9qD
YIhBu/lKvAaIAaEOk6y7zWa96wcBLeeapn+6RHpJ2F8+JBea41ipc7JgxsWEggDdvZ8cOJSAEsS+
t0A+3q0MPWe7oYr7EZP19buwKhUKSV8ZkRV6T9k+IZ3e1HHxugGptfIjU9x6d5kqVwMh/ZOWXsVz
iY36NwKVqP9nG6GnvD9tUT1Htr+sLkE3BA9WX5EmVBYD9uf4arUyGL3fw7bks79/pjm98cZO5SWQ
v37Y7ZIohQigs3bI0H3mCOsnfrhhflENBPD0PMDabrr9H+IgrKVbu2UlS0xOVp2Ok47H3kwyHkiY
mCKvgGwgD9vTwiyAfnUENDHzQozDtKMbdBYAeZSNn3DH5iie+0m7l29I7mGp2t5z6G30dQJlf5u7
75DKEpONnsQb4fC1lZrFkMANuou8awSAuQHqdiSUegzkobREHXf6XleulZf5uqqo5ewIxyQdXGGF
gg5+Vzc3jYcvYEkTW/OSrkDpU8994cBwgrzahqTcUBa/fZuUNFGiKuMTal+/+mavQHf/XLIcj39U
p79u7gCfFOtw7S/IoqEBNUx+obaEeQkh/IkCCFEnVhendLtsdqmo+MK/S7Bp2q95J8ZU3P/NJuyb
7Bu3H1u/EYDMIYv3ONoC6yTIxufndQN5RVr8cri7ZlwnxAXF/3Xuhyj3HrgO6uaZhPSeqqux24x1
91JMk85738t3NJirwg4pL1Ap1tdXHmLubh66rsd/8H9xZHwwpUMGXee7YhXB86cz2k6VO2RQ/uJ2
/F1vrBh2pgbNgOJOJasBDgp0blD2T49BmRhwceKj+YMGWy7X9odvocphJs9hBl9ZLsKI8trVUTVi
iVCV3qsCneNMqFxuByRsFl6fTo4fN+d/hlvnIXMw0LSq6OVtCj4x03LVgK62BrkIDGnLSCDoCQvT
4VOXtC7nwXlMgyUmcxj6EXpxIDK/Nly8oaAUORjU5E4wO+Me9vybCAdMQhSwWQ4JwwZ2QnoiPsgp
KdC30/eVguUs5ENQE7fUuMyICsdNNhAXtGKrF+TFia1C+FPcJVdfEXMLs389Mrn8UQDAnjFGgmBk
VV7Cyl6rX7jBA5a61p+Zw4ViN5yQSvevNfYXGK87ZypOJvXDT3ZGJ0ABldxK3L9FyCKXFCSnDFXE
NtRQMe1YA2Cc0xYYLcbhAC38FBT/Fpy2w+5lr4t2IgSfxqeDGP9b9qzCAZVApDyDNQbgIoUtL4bG
3IlX6humUBVamfigVHWgNqoW5nI31fFbSiZ6OwvIvkXRkXbEA102eokTrHkWpgCpebMalpIlq0aU
mUXMO9/Q1od166UyOxymFfwLrCDZoDM8jDBbAHod1B23w13HBZfY2pjEX3k6WqFpmb+QoaYc55xK
eDtsj0JoXE0qto+lJUP2MvN8mZ3K+DcjiD3KQJujujrbE4ErERQttQkal/HowpJlUznWDB0U2C8F
ifUI+yb/Qez1UmDm54LGI4aX6KW1bbQYxen6/e3vIEpSvVUDwqwH2SQV/NMn8N/r5T9fb/AoABH/
v51/kmT7zS27NLrORyxtVmpuewKxwLzdAGQHwW3tWbAB4oFt0rTtP5YD/9vt3Iw7/m+NfJF7dAiV
SNGCqyJxn2DnWqHMQ4kBwPhxkaIKykPHcXbiCcy2rbAlytRy4krLQg5P7mHFirhDywnuX/C7oPo2
gvapvvB9F3Xms4nR3se8rIDAPpwHdUhnruv3O3/D70rNmkyKOdS+rURYpuLw+WDzoWaCkX5J72uG
ZTY/0QEseClArtFrNXtlwCF/2sjdKbdOjZA4E7oUiiiOnOGw8GTbDEUVyG7zNEUVYvupvLWTSB4V
EEoej40/IVDcGCcCpV3jQoKpNesPDYU2aZiSpR9reMrhgyMYYSmEqDgfMDWov2yNvLKlqb5PyTUF
Q9T3XMKouZZzm3B7TTbM9ISg9zCm/8xP3vO2yrx4Eky96ToNwrjOUggza6XwzCFrn6/CKOQf4vGf
y+7naelnZsBbtnEKC1LYBF91XiNzF6CiuzNckWI7rr41gN4jVywFgBicPiZ48KTln0wK67HsuezW
3Y77/LzOXSv097a5y5opD3izvFOXTp/RLMMBnGXqPvBUYoy5u4YTQ1l7DtervVlUAIrWP3iFDF58
XuRrAar5/P8k/ujeGVYXqmQuJMe569PTwljtU7IqbBldq5fLVw3g9K0eY2l3FYULLNH8+bXh4CsA
aaEkZaPYtyVrvYCGVdi9KVoxYwC8iKHWED+mmu7EzdVtRtO08pDYu20ugrUN3LQQNq5knSfd+18A
ReFALwV9sbD2hEYNlA30huZhRx++jQlSV5VV0LtXczAFXtVfE13j+ONi/U0u+lWrlp5SPo2htRbc
AwSuYjfequfuGIKu9VW5IJCaT3LZvFVaCO2PHS+T4nYjgoL2HoyUyzZlFHHTGXCK72Bs7FkopiHT
tU5L1M8WEnxenJBmjfitVAIYBiMRqqWyvXnErbAqo4B8cOT1CfK7+xpTl9/JIHcTwyfmXRSnwHPV
jXeqRWUL4SeF+NmM6myStrrvMPqPNvXrhECMd8HRFKAQFwTo6TBgk5WujgHqhuq8nA2l26msmTb6
zW3AHt3F2ETGdSg1x4ATycA1H93OSRshADoKjB3oYoPBPGIqRywI4DhOOAigIgB1vjsdGqXauZOT
jOuUe5gnBpkTjk/2VHnB8D9UPyHAj5A/yHWAZgMVCAyLKob7EETLFmo9gwPvA3ciJY6xIFoWJC4O
zX+EzUy5WEo44SHAQ2yCqOXMQCbCJsJzd/4ORcwVLRPJHF0bn+woEUhD4DVahm7hIR3zp7rYqzyf
76rPi4h4DlUJU3WVxtrrPMsL1Y6gHV1oogmnV8rC3hsOpTB2H2PSZ5QXSA7D/k/x0sUS9YPw2S97
tSYsFbNTmRIcL9+pwNZXGUwsHdU/W0Q0jgUb+TPBQsHS5jnQs9RbQuu7wPECciHvv8fihfh+0cSP
e9ERfST2LLKCNzoy0bSPQ2gcXlpKE0T57TzskLLP/qb095+h3GSNb/f7FVJjbp2dnygSZHMiWbO9
TyL/otN8ui2tEieXICBTSXjaL8hAedUVRa9gGEA=
`protect end_protected

