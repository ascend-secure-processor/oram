

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jMx4Fl3l8KBQNYNqr/FVwCB814jrLPlSMTtdpxWTbrcWy6MoMrE6hMAPUlKO8okoavoipLMUngXC
XN17vI8fQg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aipMRgWa1rLI6xlddDe9OYjSp6k6BxsQ9ZtecDrpvJW6FKSe6DViUukadT90rsuE4SNGXiJUBaKP
ZNpkB2uzO4DU9Ele/ETZBjlMnJjQMxacvuPBMerAlJDeHKlFFlrtmgPwvIUtS1fpd7GSMUC8olc6
HJph/XkgXWDuELFZD1Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gXQo0gvMYVrU6gEXhtcf9+wfQLg0tJRl2ucI4C/MIVobuluaEcLuSXx3jN/jlkEelNCJP1EaMfV5
S+EUf4G2E3VepWY36OFSBE3A7S1m8/uonA0AVId7ZbO6eBEQMCNHKMONQnjfcIJfYzQwx5Y5GOCT
ImIxUVnACgXatld6wtAvms4gFBWGhJu3kXH0t/PurlgEDzOOlzFoMbrPIFgs8rNKT1u6Y7MRLNgt
VrOW3h1vZjzRFOQIuq5ULxGsjOeaz7q4JkVco1zCoaR+LRzbpcDH6fxnPctgmIpgz8aWvZ25BpYL
WY36x8VTMkSliEtgHMKZp2wuU9ZRTcZ6+XTrkA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C/uC+CRiT9H0O963L06rxOp1FJALrloHNqGcGGkg0UD9n7idNa5AHk/0b5QAmnFueUHxPeH6W5/1
aY+ZzTd3JoCk2LETUbDcrrauUjygugVcXBG+KcD/EMlAAZi35ROjH7xJc59PpkBieZGAgoNDRdSu
CvusBPKAGhyLhWrz6IM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cd92v5N9UnRL+aOxuo8bJe4fH1sy8VaoTalRHuRgDNBhDsfmtinD5ULXtFegBmFrl2n66yAgwqXd
PFZMACrcRbJO8LCnCYj3jwxlc8DZvnsiOGa6IDpNFtYYgGLxVJn+5gZbOad6QgpukBaF/07Q1LP3
l6iNefmd/rXLpCadRHoDZuKCZDbs115s+krqdgscnKVWVMSn/ck0kcUPf28JQbrizRPmKYzNFF0m
2d7ubkTOe6Zn1kr/dXE+1ybDR1r1u07X7jNiSCloPN6Bv93rdWWo5n3qrSCq8dAqj5Z3vi/K6tnd
96UsM7VMsuqbwqZ6u24WLLeF3RWgLlqUq+5QYQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61984)
`protect data_block
ePt+ClsLx/2y34VpDZ/tEU34k2lcR/4gE1639kFHkUiI2YhVd3shsJHEr3DcSs3UyoIpJvHobsuF
CPU09iatuyiRFgCfgaBAfNatxZNOGWhrcY8lNhLKZrfOFFJyGYbYTgCB8rizYLbPUlhAGpj9e+mc
Q7751A6oRGj02i8yh3orkiTCRkvREFc77U5EoMh+nK+AGQa92gatVkDzE9IM31qQbUGLbw8K9BdZ
++fCvvfJf/KuwvxaGkfPGMes90/539uN61Hmr+UZuaxDQRkDePOkbniaGWI8sQM/NKkT2cCFIORO
ccqAjMgxeYVFbT1KrmGGh0zfAzU1Fk+xy9wt6NFlHgG6hjF/ALJqzC5kkqeR5pe8N22Hd/9/katx
i7lXzql+KVLwjhGKa3d16fSu3clQm7bsA1p4sn27O6CENHf5R8Kp1z2Txa/FEoYOnXS8725ZHo5P
6Vt8v13QTWOmwEmRrIQGWEMns4KwrrSBhKCM+SSsaeN0+u83OiaBfn/eGQBCcy6AmaE2tGAuMKOA
goJs4gq3Ke6yrcty9O8manL1axl3/HeRIj7oxEDJFn1gBBq0/BXmJtGe28mXerEe5H5QrjEMWvm6
ZeEHg6n4s/XkTpe1E1zNqLdUXF617TVhEIbI8DdvgSUSuJrFqWWIt0qTeW5k4G/3/Zgf6jbEle37
NvihZfNmtzqCpdGs+nKQhZTJra469utdeS1fGgiucAzAfnjg0Cl6tu6PGw+vWs4qJRNya0VAUHUI
XhvJp8dqGBDyMDKam28FFyj0NM6DPNWe93jTFDyka8OA3pVYr5PQPDhxIWdS0kEeX3FzGgyQXL0p
R3dJ6iY0zsAZYcbW2BL+BIWVY8JrNdYlX27o1eG6uRcVgkXfQikk9p/uMyk8nPumwTKyjnNXGBpO
NRbwPXVLhdbv6nZmMvfcecTnFGd6bOVqOcenEmKZypDbQwScbjOTRACN3vYGmwGsTLm9YINrKJxG
UYsARIANUuk+Rz7ArHFFYin6PXUuaMGLfOdwJkDypqwOZLcWPQtE7MejfzTNptLJ2L4b3ULqZNNL
/3HHEsjFsZF/n9uc/8AlB5+kgI60vLEK/mFurBMzbSOjDgpFecRLozdU/gjHIsh7JtuafCAqMwh3
I6OZt0/HoUMwsqSBsr1qTD+0McHdtLZsVo+KQlyCP39VNj1RkhVQgOEDucJ63Lzusk6Ehwlpl2GU
rDUWCIrtRPuLdMAWmrs+x1ggn3SbyCPy33FLuQMAay5uphb4DVUlkDbos8vkRvXl4VFLwq2SEH3i
N3M1Uy0gp00zZdWlmQ/fc8gtLssjv6KJAPriHoaWLCNgv35W9hcrbbsTcROuU5M+0byjawtZB6IJ
9PAyaLsrpGHsx5pDCXLcuyETxYWH5NqSbaA3DFsbCY++h90a2tYoG3KxhlvZMmV3ryG3/Zkk4xjJ
EWE8rxgz+ikxBpgBtJah7ztZHokBkIuh2WZ2y4Ie9C5pwJjtzgtKxPYGvoCgwPa9T0Uyu08Pvn/t
5F3dWbF2L+8WH8BwJCkLjj7mI+PyyzyERGU/hvy1EsTTR4qGF2UdqKpaozdPtjwiTM6n/n76i1HX
+14ctRANIFHrZKVIxnVJpNnvr4eSYTtdK7MJLUq9w7seahqKQzI6Sjf1TeYVwJKo4HEfNx/sRV4j
b+U4oRNU1MtTlEv6TrIEjgztxzBhR4/xnbGsrVoNkErOzVLrnGVo2Lj9/XKiW7hEKRqMIhBtQ8M0
mOwNlfs3K4K20kd3020H7ADgDcopL3txgLLsZpRC/O92283RAODh62OkZ5SdjAQUUHgh5sAdrA/4
NKEgTZOHtZbzxo+c2PPo93Vgo7zgQ8Kd81KKK9DNl1khUZPFxxRomvC33830kkjCLruczatUXy9A
NH2NE94YNOCpRygAsHx3FX+Dk5KyWAszRK5/o16dgvHXhMPTessuCtw813exhkoQ2CIT2VaxVTXw
qVnes2PdLeKsgd9zASOow9whn0yT5dnr8tAsN2H0AC2xdApa/nHJRA4fuDU8xQJqV0m1ZS9gYCW4
bRXpSsruHaqr9ZhD83S+OXymyvBs3gvklen+ob+RdNgr18z60xwi1OMfdpzLIP++4ubZSep5WfiI
fT18r+tvWg2y+f2FurUSyZKGdDfTMrmXQGhjR7UnLYNmr45605HDqwGhmAo/XyyUebxP7/etvvkU
coFZpEzTM9/aFH9ldpQbEb4WY9jSMqxgEkZV1P5DWGFU1e72sZTDTZ/onAvu38JZTFQ8t4AnNNNK
JWH4Vb0Mq5g8KdRBylpD8zcJEYVu3fXTD8eVS6F6hv+Z03Gw8NZcfaG/znPZXFhTKxUmHYeMkOQe
vM6mdCDq7U8LT/Yf1PCjp+O0091AvicYHOWsPO4rPSq7ZqaJHKoxIIXTVLL7ZaSo451249QJ1cro
Q6qby/bMfBeYf6CjL+S7ydQms5BE6IEmRFjnpEqvM9GqWFuEd4QudSkuhI41EjPKy4vV51o/lhoI
d04Q4s7AwzY2NXw67esYFzoNyUDkk0eqcuPdr06M+SmDK561MTuIv5ExeqTAYAN104P0iS4ASukg
Ymkc2vB5UyLQSkaBF0is9CL8fo0VU43HROrNBRdRUvbo0vKgFp4ZsYIyTU1WF/89x7oa5PDzWUGm
9d9ADeW5alGZLH31hjZzJx1L8ojo6ZEvn+1THIY+JF8asVrRifsyEnwDp/+CT7KEVK5swsZmYneA
4UwIubNBtLGP7MSQ5iTibGiyOBdQjRL51/0CfqJj5bTRRfakqNK2w63i8iCUiCw8lGf9VhoSLsNx
i1uONT6dJ+gnQ0LTkJnEtzkn3v9x3v6KoEzW5MkTB9oASgOREt9k1SCxLEn4GdVCIa5NZTH6/UJC
OnSYcIVGYLdjGnIn2wVJ3ZCC4sTppImhLjDsxsg+kgOffvt6ra3PI9epvBTYJX92R27gTjyil0OU
8dDADyOiv0TA2Zdg1pYymjL7rYr37bBiSnU6UYG4AjMESxzPvMa2lprFyQxMQZYvQhxHAMy6fwAg
+gJGCXpcUwqNb2GJGAkPTF3GH8HtoZfi8p5kecbxq1UtTbqty6wMLbDHsHukE7TVTTrRPKe0ydKx
GqUEZxgbhuUMIcDmI3KbLvVMyC3qpHMExtc7a2kT5kwC9LYHVOUAWZ53dVnUfgFIs2G1a9prk85B
Mt5HrBpZxNkv41LfnuHqZxu6SrM2tfHZUMk06hCRTkGJppEwWsYRL4EprBhTqcPvdg1TCzU6mGQK
TZaXLWXzhMJHySG0KzniA3RQu7kQvZHIQhKMQTSXOJ5L/V3bVtA3dBLUNY1p0xGvsDGIR/ErPveB
vzqPATmDZT9nexDpx6BUG88Lc43Fi5w74FMk2/7peY+zkrugF3nLpgW9eEFTQF1J+OsH/9TPlisI
UTpVMCjJHoyqLVVSyJRwhsPR3zydSQkMRC94oen/L+IFdVloNXl+z0Szjkvfqh5+FIeYng/moGsP
/45DNDmY5n3tYAvP5NhpqGtToP0wTB5mWRaUTqr7e0EPjCZ/ZmNI/NloEKk+DTVmP3qiVEZWFALb
ZEAkE6KgIvVCFBPUFU1+P5Hh8gPHbPHRNdb+uiBG4QrwpMs0ZmchvUfVENRZ40WRy6whYrtrlF6I
69S20m+WYn6f45NvRasmFhyKV1JfxMQ0hXRbI85Y6XbvTf4Rs30Hd62hAy87OI+yGjaBOJg1hKCd
kiYVRYTnCH2DMJq4ilknH45qmYrulfxrloptuLADWOYzQcynFeMf/MtlSWrnMuO1gocMt3hv7/4b
plzCLEKu1xbHDK1ALN/xDjkOqnBQhsgvvF0tTScR8O1VrbjaTJomn2kkdfN7E/4gnl6OAO4YyD/l
xl8xmT63Cj7I1ooR5gkOWYquv0waEMsyT9PrUZHGdfLzhf2rpSCLfo+D25obRQkS15K0Nf7SzrJ1
OT05f7QoUk/hWrVTUq2GKGILcOyhPY73GYcwnodu29ygdgHbXOlgtHSTTyt+PGqg61rq1SC10Vxh
uGE3h/tfDkOptZ3mMB/Xd8HH7aQOWvg6EuqmUm6tlVFxCF4XetXDAcUmjk5k8/GSsbkvOAdg96mz
2fISHICfsvsfqg+zatRPKPkj099t+WRT/S3VC+o2jUJeeWQ3RLXCT85z6WD9cluQ+ow/PK4TDtUF
TuKPEox1SLJ912lFZK2Yhnfet6+MChBl9NvwGAfS71GWPbTz9OWqZQK9WzfmK20leUwCvFAkpW0c
aszeLqKmj3iWvvhafguLaesJpek9FZJhWIJ6qvBJSfKU5HGOk89CGgvDKwmqBNEbbDQLKehuJSY/
IvmNjS1zMd0KU5Xwlfh0HZ9Uz4iJG5TsvTYLi/XfmhUJE4Aku5jLxzPzXTeIE2C8gPW+HtS4T7ON
xOSXJRwZnHo6Hva/i65SObYvmeAFIy4ASSIGVgyVL7+06MbUe61adypkCucxY39Dco8L6O419rK6
Ewk9Vws+o3KDQRCi1IGROBdZEM1b85rfxO+779lRcH8I9aR4bvxCggNOa5/XR+nVdRfIrpw2V18G
8RmIn1ZCmm0qTS6VhkDWiBdng6m5MTI7s2UdaxyylkbBJOWxuo+2GeqT8DCz8197sEO9SuOIx0ye
uH5H+0e+NxPcb+QB0LkyeBnSg2A6sO0zM5wXNHWLchTzUCede4P1NNGzxdCR5rbL+L9GLeEIaMkw
2VgdxWDwPXK6hSQGobk1AdZf3H7Hpv6l1FzHLDBCXZGUzzaCoR/LggCgqogO5h9puiWJKHSmYqjT
1RAVKwmIhv8f+zbAV6Wi7s7AtDLcZEhpOImdL7jWXpJL7np62GEvK1Efr7MwvzFmp5ENYxD3v+bR
nkH17l+QN1viDK5IhLhJH65gZUaroXAKCKKUilul5uKO38sfy6vkmsmO/34+dqP798lRLcQjuYGn
VS2hnsrhwMDZBD7tsUujjyX7+J5KyPeaAtPXK5/pAkx8kYIVxLNzVw5u2ZqiUSWENRY3UCJTYcHv
XQlFJq2ot2RAJAJa0LIeY/8+thgct/+UR8Xps71czJxB/BBW4rpiOq5mVopsJLF5IVkhJjXbIl48
k7bPZuaT2ACBVsOY919qnSk6aTRLDHVc/Un72wo1HtsXYXygnoP/xH5P+0xjuLsgK5jwVWUB2fZb
9WojIIyqTCnwTDAhvaVtiEqljftncNBWsu0bCFeYB8X2MLygra8mdc02EJI2Kzqqmxr1U33T8gDd
qLv/esVIv671pUl1j1W6EuSJ3nyg/Dm0Nin6bc2OAqKHwZemnZsuHhuMQ/LWdqsP3hD3eFRPaQL/
Q4R2vtdJI1xWraji25i6qAyQWbpr1P6cyLiXLctbvezrIEeMuqHDE71Yk6s/Ha4BWanPaunQwuT0
L4+c724qp2C9IgBpeWY/VEKe815mU3zp3Y2vxsGPF+rtCJupESk6149B3vCO7NSafGiyVSAD8P/D
1iwXs5rceGCn81z/xUmSZggqEjbQomUkmugUP8dN5Os771NCao/veGPoGVKVhPvdgAUmylAt8lY/
gs5CXED+JnKRiIfnMTUkr3D8qkA6oDzFrVQVJ0ZS9BQD+ddpQQ1wINASPr9On3QFDQ4QwChw57CV
5IbkhC4nR2PBfzKB5y3hwV7xwf3UXxPlaJzMazhEZPJLBkXk/jKDfg3AxJ4tjXK1WTTMIJzLeSjh
02NtHBMQEwLT/mDgbAIBwtpo9ebsAvzbYaiRk/Wuv4x/bQLEid3HCKtHgB46zsEAoiIcG1ThY+cl
2WwceJ/firwWWIw4jET6SqRGHuZidFImC3YN8ERj23U7hflCOMD2Zq4HjEi9xV2wt02JusUn+DzD
cib13b3I5kWKW6DLKEcPQluOaTgiwdFBwLdsIqXcG94Nq49zH16INWVNpWa4w+xkT2dNRyzW/HSr
0uTqWTuDoIeLJTyBLTxWP1AM6+mAJLmwED5JbeGeFuh9mChqDNMbdDH0W6xJGIz68hBjKybfYrfe
Cbbwe0w+Gvi3M0+6nVq+2+kUZO17AlagEP+LvHbWGo9RvCphYFq9TINO/K2gd7DAt4P9H+Ocl5vo
5wCKTV1pU7iM+B9PTA8w5cDcoJuZByKdlSy/kGH76EP8Oss6przhR4d73o8EyLS9B+S24D2drZB3
7ZpBMOO4W4oj2XpUgHt4nUeFyiUMriHbvdcRPOfiPeVcDWosAWDkUB8VsF44oOhLTiyWQsv6PAqk
/cjIxF1eqSfrMoy9NNSvPSKvS6cONjye4bArZsAnYBWTI9C5xEB+sd+sHVJqUNKWBEcSm87+iCOo
YuyGcA1oA0cnrbgoipkrLKT4D+iuVHddyaeqOlWrrsliVQJQSfGmmCV12yCtNLfP/LVDVYRQ92NK
/kw1lUqrYUJcOGVgYaqSECwsrUDgWFu4DY8N3M3aI3aj7udUsKqIy3mLmCTP1n0DTRyhXAPpGtO3
JicEoqan6Aem2Ys+UL56ulyjXPrc9FAYsv6rCHBeKHZ0Cq6irYGn5l1cvctDijajf9M48psw/FXb
0du631qgeH7/wIxDqSKEdzgvMMmPN5o6JKi2gvA6M/vYfmrkLFyatOuhdJhWa5x7+aPme9zxjl2C
jVStencA8GayAJ6liZw8mEBVt4lKOVi1pIvZKhaHchh5ythuL1yHQSWnaS/vOemcHFQZZPBnI7Ab
F9nSLAfepdh9v5pCNkU7XZ54Oj1PS9EHGJjfV97iuk2u3KlASZZ3+OjBtqagn3KbRh27X1xOulue
0sK+2Gtg5bahzZK/p9Qhu2mAonTtyl09m7Y7S9PaCRi2+Ru5AezqyO6Pm3tIulF8dQJR61DBj1Wx
2dHWHzijuprW+gHfquvWDG8sKFkWlq+qqIkCAx1Cu32p/2hjAQIRIT4vDs4h8tVf7Gli+yBVBAOy
nrx8hbe+nQsSA+tr4JgVi7aP/TVeyaheExJDvCTyRRwrXj6q8ebgZ4Xy904EJquCvmaAJSY2uT6e
1ioQ6dCow6Eg2DDwkg7JUWSVxYTS/IXdiAfCEUNUJoEJdQGpGhuYmtNHJQWJGS30B7/AznpZSspD
xslj98kDSFpHsBSFWPhVetzS4qzu9wMD5Xa4588YlZkGlQapPLWnyzmkYhXHFpwTTLZpIyO61kMl
ExmvvKOnWhH11N6wiDzUJlq/YOgsGSIS0Ad8UQkQAN4XuytugYO/9QpoZGpHSBdFfKGuFmwxjLYH
E8bJIAFn7dcAmCdhY3bSr7W83liW1hNycGEELTHvkv9V6JLxZBUGtxA/eeWKZe00jbHodZie8/Fs
2k2xQ1CbTjgeaoTrcNwo5KFo18jFTvtpT2SF/sP9oQ7bQpyUv0PkIMARjs4vPHyC6ve5WkTzs9cU
F2f7fuu+4/EH0ds76oSevJuWfkqusz4PIwDOxb93vpJB6+ghwWvPrmu043GRxMnuJFUkUvakU3Rl
m2dFf3LnO1JH/9o9OueyufqKChyYWhy3FeaP3o9OT88iQPl5Jjdlay/x9F5iJsxwyU3AitZN83vM
5ZHf6NLgr/xAV2kUjHz5PfQGHhJvSDdTVIo0OgdHAe0idx1badLJuXTEQQORRds8dwNY0dQUCKrN
RGkzGxyqanxNQTTMLQ8P4fLFirEJfdAOS+tzyk0PpAlbtKtgh0639pyVf8IFPx6LOuE/lHEGC7Ur
T/Hn5Wvu69Tc2XbwFQvE5QgaAfw4jzwlRd1Mj8nmWPYkM1QYW9chDLqDBtSmCkrLSo+9RMX/DM73
OFAFSPe5TE31VXP6z0+0flDa+dTkfE7d9lpc7Oiwr0gusqaquHH8iccQal5GblBjKrI9zHeo7cCH
iF2ub91D92LFrlfM/plT43zM4ZR8NaILr8jQSsKoG+3fdX+r7066y+xCbGJ5jVysLzHSrbbYHK3f
wAFvbUS/R4CJYY+14hViBlOUiRj/UnujhCCguwBb7ZKA03JFqQiQni+aRBtVDfdiOp1Xl2Aaguo0
Au6d/b1C/l9A9W4iXYCtvt0ok0nlEKG9X+aplU5WAQRnETYAdMFz4Fydt8vb7UWqcgEbdbyQwCsC
4AWhyKO6VSnEX4jU4yWZgMBUcTwkPKMadgS10rAZ4zGfUCIgZTWhKaSO4f/0NcaJgqqDpwwVcXtb
evr01Vz9/bhM8XFPKIKzRWwdsoYO+mthog2XVgtJCagHTn4r6KyHwI1eZAIZBl+9hTxJxPanH4Qz
Ww4cVDw0yq8+CN/m1m3r1yiiul3In3qLlGt0je5fBKso0enCcUpMC8H+QIbRY4l8lTq8K1xQwXMQ
tftQVZapfeUYsf6jz/XJMeUOX6sLxpH1GGkgRpOURbZlrSUqnP9i4J43OJbQI/j5XfWDf68RHGRQ
vcabGIInHpU4KdzfEdKKf1wTfT+Ido62+rsYOiNGXjmL5r60vjoACUn+KRRQyRqLJ2K8h6V5Hwm0
b2lOG00qv69Ymreq4AouaGNH4GZOet+yX+xJhV8Us+dcwjxJL7Zsc+6d2lBuarPYn9O+/hbuSaVn
SaLG0svodN5Wdc+4qOXh0gKTmPL2fh4wrjEGvq7QmVvD6iiJ9Qd5eeyxAk2n0FElG1K88ePhZEow
QbvOTQ/uOSrKVgcbnrmhDm6GEgm7lSJRuZVdnMcUpOK1lDuO2PbTyB89K81NSZ109WaHFkELX1CD
IA3g32+HwPrgGU8jsPs0UKedLzxpfc8/YDwixHpr3YgXzYRCH1ovkeMpP/upP4rv4seIs6wr7TfY
5cfoL1fMg8s9ylkEd+AjlBS1MO4ix3HaomPzDHt4sAQaaKtBJIOZvzWaL7eYQErBTD7ZIhVSkC5X
CeMZmE9aXiYiY8IpVxKSiLRTWKLXHvaxBgqj3crZaFMuyukoT7rlxY5ElfeITVeJrOhK23sm5MUw
QIQU7NDR9GdD4W+FBwrcJC5UcFqwV5lMSQMNky31UqzG0CaDAw7Fn3B40Yo0a1ecWCDwHi7cClea
+kj2EPc/YOiFOce0a8IxR/M/BObtzO88dPY8A70RxKTU9f4HhhPPD4CouCl2G3PRUK4PQkl1euSw
AczFMMRwj3N0JoEVRrmzDLoPFFlSA0ixuEjki2n/lyohvA4BC8I07L8qKdWwWsm4CGDHG/lkVPtH
AYYQBAVQVtbldJ3bGdQOodDGsjG9PgsYq6mCkpqtTXV7TKRb2/F3Ituda2iBn20h9F5KTX6AF3mO
zZDgsrC0kyBa0dqDSTbztXFgec6+gC5Ak+zzMTIeweP9lu8QhGdYwvNXNjevj+PT3r0QTCIG54O6
BlIv23qSaWcHRA5Cqeev8i/j794UKSJ9Xw041vOowDQadoMHGcbYzpnuSbf4JOkO9uHBC/47b/aO
wl2+WWkUlC1WdQyWI/bITZg1nyIu5q1ggpAjJan6d0xt4JKqNqkhfC26IhA7jJPqU1M3y2GQZg50
QqGUuqjAlb2iqDQtFRHLtRsjPu6KO3goBN9e6bCc5Y4fKFa+JsABzD0UytiB6EWsM9oI84BPpGU1
oDhSyeXTkz3migraav7EKP3kGErQlKlD8QdTUZievm5DWJCBBB+ES7C5hXygMbkFfQ3E604wcF/y
6MirOYJlKhxlTCU7kjv54Fz8sIDnTZtcWnsgrrFWGevj40A6xUnDrtZHx4szI5wROOIQEEJohGrg
8Q3x5EQCwJOkzBwOAmM9aQxVb5ykkt4/Dycd7tuMF3517l6q8gywh8uTw5/3DQKPNS9rsSBdGKaz
YHYVcDEXsUsHCMYKVchMLr+0NscE7cJeUuLFPW0mWm6Imv8d2mKgvzYxAWCIeOd/CsBPQGuagS2K
wsrS3HSt3YEx9YQTdnLeChuhAAF5dTH/ah7IJu5cKfIuZYBOXYaPbUhZxVHQ9YF1XiIQgcAHeVT/
Y9bUCc+kLheSVc4iZbS2U7kYg6maCjDUmkJXwhaxaBkxYEGq3hh7lG9OvwRRVTpSPBLeWe5Itk1I
QRhUZhybgPGCVjLzBMLQ8Ll8Pc6UUpgrojDRy/4ngsP12rslthMJjcozoM4SzwqrinbZ+V7BjQku
/lt7lRFuXHFeIOKGX5P7/UAk9TGAiNXyDayCqY3uhvBSARgLvMlLLAtEijAgss8BSvTPdOSgMr1B
hzUpAmJud+OtnOjNeBDrZeVjrfwryY2gWajFG9cjH4lYoPcTO55uDX/yn2DukBHeQ6ArSCqUxm5y
5mB7CHR87vjeWh+j0l2i0fP2mJh6xOf6th4S5OLtw6schw5yFuI4YZB7LeKdkfFYeww5OqYD6nqA
bu+pz2JtxV4W8FRksaZU9BwZPdt+mhhzTDFVY+JN8muPBctejTveFYtAOZHmZJwJ+MjqZmT4MeT9
aj3iAegl3fd62yba6haDOWxienVW/WTZqETYOe7WPXFWoVQpAMoidMAxPjN7fLST+kAj4M3doDwk
h+jy9Yp5w6wTa/YkdW9GvSIzK+JfuQ5+eogVrH9Y22M/9fJSHDASaShoeAE99iSEk07vvbYH/78g
G7lqFQ0EvogWtZ4spwLxB0NiykQLcNMuQFmJuFVk06V+mHN+/yvm65rtZO9OsZ9s7GzoI9yjlIMa
B+K5ScD/kzhY66W0fPZ7TLGVsUZB5q4u5oGXVryM4aVXI9q9AwZrZvqxw+r7KhOBDbqc9GNEAgYk
cKhyDNd1J1ME+XuzI/KP8RFRzENJnPawM4kYzqlWTm5HtAojCnIocK1RK/qkKSPhkrFH7yAJPqLa
0xa2eyFRIoAzpTFrxgmSKFsKOQM8SlJXLRCh/1vqM+QVwaSSOpFyrUckvsogcwU2sIl5gC6QBY2r
Co+LICoKu5vye5U+2tAZ4j9Xw2OBNNFMKSQ4iWLbl97+jFjA972PMwdbx2SUI3TMovm/hVajamFc
WlUiR+UKpNBVG0Tcnu+5gBs+zsybUckybdAyRDf1yQmhfRoo/mGIcs7d1NRwKH/MtYUc4w9QGZoV
/lvMzw1NFhNEJS/zORY0xYv9vI05jaqaHn/F67BR+fdjJinmhvDhn5ib2DbV4avSPOR6IDPaWiJL
8lcIGiL7rktRzfVMJZefySnn7HPAp3FXG1NW5v+HWp6PonZ+Dcm5JgoQgkW2KEsHcK21s2eBuSAB
bvrfo3hCQOvEp+1sqU26PgyvauC+skD02QrmCk1UjK7sKTpeHVUEzryhrdIOBX73/Hdy0njhZGc5
r4K3kf4qR1TNTtyj1V7IOIfzJ7IN92F8dIKewov54gtAfTu+lRIqlK7ch4CzK5d8b7g6P6+z1j8l
5fZBtw8ZIXS1OloC16yYMAPiOUXwjrBggommmpA5bqVu1eZWFURdlcjqmWrub0oH71zMH18FTc+W
e4YqiQNZWgIg+imODwQyv6qyDQsKLTjXfWToGKuQqU84/YKQooV3ORBhLIGOqZ4v/ddRuD46Dlys
trAjAgJTTRj+HM1W+bUUIZjj8uL7+6SheuPhlRqeN35YWdy+KixDsCI0+MIEBUxAVDNH6N4OWx5/
5HwKcgVrn4aTEICRA61BNyWDMu4cYXxvBqr3QODVNWKCIZbnXha76zfQ+xRv/1xTPgwYvVHclBqy
CxOv0uI6IfJ+sOx6g41L+PzNUpO67Cpz+avKFNXVo8k49plSje1ToTYqZAEciqmfE+zMaQwMVd5V
U/1J8dfvhmWWia6P6MlZf+uROfko64oJbvqa0UEUGWnfke6awoVkRrDBrUsBfdcJQ2mLBrJLxh6m
WMINYv7BfhNpZcHxnpkAcd0kNO0xfCbDxbZJH6HW4mGLNSP81nvy1FNFc9rPnK6MbCM/beqL+G0Y
piO0qvBgtA8r1GKQzyefXeTgzUKMikLnuEzjO6pmKyfbjYfQerJGEr8shakOxM6qs9f/B6vfJX1u
I3ydgR78on/tmYsH+8NoHsRaHrjaLKhPGAt+788XUIfaTSmNSQcKT6iULVzNlWLjx7RSW17Xz60v
Apv5p8LvxxO5wXH1GsmLg2rvlGORP4w32dh8kirTfP3Wb2HvearSn6MFVhR4WJD7fmD8Z6VwV61o
yHdDEmlChe85SHI71HX8fpxIDi7sOa01aGUQD8n7uyCpuZwFIxgraQRjLAXYd8JOCqgHSkKW0aiF
illepauiKxMq1PZjMZiBe2LZ5aIEvTmX6Aw8hMUBU1nQ6S6ua23+lcEo3ITkOF0WSI/qhlxvrHpP
CSDz9G/Py/NrfqfoKsIJlEuxieuOtm1qisZasLy8gwaH33hdrnnVN6VCleD2ehfkS3YujUxmKMnZ
5wDTlSMUUfMbJCLR/EBjsJwmlsY3YuqUsdkh99yAYYUprJDHdg+8Djq1DDmt8uFpnIwcd1wTd877
J34YCfxVCfAWK6SheE1/hbGLVBGYCWtV0nXgpUhsoHzKi58g27MuQQ5OixaWwa6dI8D/PJY6vPKe
MJTYP3P0H39Khv3bDWLT+7CWwWDJQcvyoSUm8DUgg9Qyuq2wOq05YgIDY4xWB2hkmJcGgbyJHpqr
580BHYXrcCKVCojhG/4hKItYfbji+ohZIEXxyQuapAHIAEVJd1W5AwEyjMrSfxuRIjwKen3TY90Y
RBiH7RFeDdVTKQ+B7B441SrUXQ6hZj4NCwlRO/77FmnPdszGDcjiGxS0rsJTKF2WCAUMPNQQx1k0
h+PdA4DJ88zlYc0Hy1PB1KNLp8eGN9knmK9splGPdQ4NVvU5wMTTNuRCNw/E0o2UXk9WbsL+0ljx
T4CBhkzBMDZTKMnILT75QIpkgyyqmJq6l010THsGlanD7ZyrhR+RQ2w/MyF6CpfffdUxtwkJIePo
CGatXgmv3pa9bFB5uA6brEPB2EUlxGQP1eaKOEm+FDAdlj6GXuX5GV4uVa7YDMnUsq/olIxdfOJI
+WteFfdECCK1z3Id04eKcRbEDDUsi0zBL7haJ6fexDEgRxmtJZgX8NCAskCzWdtXG1B8dbzl1t0O
Akt1xAVZL+I1RuIYANQ8eMT58LTn9SAoZgNupAB5M1kGDMwpMzySFQt21z3aBi4g1SX2EW5Pq7Yb
aX46GAAcCbAaJitnsq6SXVff5E0wJrfE8/IUgeLLy6Xbt2jcOw2pnv2ARQM89Yt8AovVqlBi9JRc
kCNgd5IZ8abN1f58i9wSNBnqXJBENzIETnzuUZT18an+yO+OQb6bqST1j3zUm1iiCHil8VZRKsnX
548cDMhTmHOLjMyA/f+xRQTRyl6oEG6QdLmetJoaKUpEDnW8w91rcN1/FT1es+2TC34xCa1c98MQ
JeriNUMWhTllsDHV8qdDtTIzh1CUpoYIuhfdYqG+qKmZ3lqIPrKERVLKas5neDGv3Q8DEu5WmGxv
GF2yi/bn/sgTwjLS9Y1k7rVMe479pSUD+kyEUfxTRySgM7+FrrIsJ5pmQ7mnUdeFI/5jsfmWwa/j
yz7wbXAPeBMfFC6breS3SlAszjTQe6LbFG40iq2bTTXkHDNOY5xEHh2juNhoN3dPiZ/O37M2DvJq
RwRE1DbO8L1ntECM9iig2ou8zEOaEfsNTQsj0zwucHsmcmIQvxprEIJVDjpRE+Khq/Z/0x7AGuhB
t/LJ7VlomK2GwCasVAzIvNVDrHyT2zwIrCQclQ82toJ4hW6AIJmNtjxJEAQgTRWAOrnm5WIG2U9S
CB8UkEO1hMr3B9y3+qLDjAkn55C/ThLaPS9pYgIDUn7HUGD3kJpr2gmKyPC5h5usUkWyRZgm/6At
WJpv+/anglUXnRFkdI3pMU8N8Z934rtr8Dp4ovEwnaOKOYcmBSsB8+fBumW6AipgbeFILy7i2yra
QqU2kiNDZf58/WtU/JtmDfiKxbrG8HlU+QWgoqUPU0XgXr5CyW05+6lDah+BqyuIEy7YGJs6FwGk
wsZzE0hWBcizKONP2L84rZtOL3GSVO72u7Qcm8B8mY28GF6qKFtk7+qgr0ySxCKF2gc+LBYVS0sq
DjUTbSL6nnOFs9IvF1BmzpXHZ87nlzWIcQE8Di00T1EJVXeYZG/pJ3GO5uV1fBgH/yiObFoOngy/
h/NvM10yBrUO+dXKJhotnTsXwiN0MwR4NprnW5mEZ7QQzFR6+IESXUTY9D+o6Kn0mAJU3hZVEA1V
BO9pCJzTKmvXSIySGLxl0WKKEnhfagdMQTGuGYqkmiEFvSio2ukO/EyJnbZg16kDbF+R/WjlB3Lt
zQfwiM5h/gX8MlCRELClTLQoxkx7XYrUkSumVAXE511+NvOJw2E0L3eMFyg1iWldizHDyifOYsWJ
/7HxFr3k9KshX6e+tL24qbbk7Pf8wMTPvqTVtkbpZNejzYHhnSoaLYWRJAgGzmFtPhpV4VqUb2K9
LIWUflQ8T2xJAPle+ZNjRYSvjsx/FFLcPCgrfQBu5xmU0P0I+vbvvp66xNNlw2AHB3OVn9PKVqoi
zzvwh/licYIy6yXTSyysDtCPswZT+N3b238ovOJNak5VpYG7WzMmX4EA7XV0gGB1p0hOtrmmI8Zp
6McuiB4ucSrxAb9ox/+w+hRvtKH7hFJ7n0lJHu70jCQJ3u0xVGIIu5heJ05/FSycDeULVbB3Qddb
v1K9vvKzyj7DlwUIM3JCv0p2B/NHvPZe7n5w/OEFrFbJXvP4cd+CDKXVATf2gB+IFDjd/5NAhCW/
g6fgVc3Sq/b+Kyx35KQ4/oF8ObhLepdUU24525P7+PGq/AachgEu+wSjsArNyQP4cuG7HmLUzmSo
GbiTPsk4ng7hX1rotIRqhOsb45KerRdNhFm+axEy10MqVxBJRMPg4dAU8Y7c7cW5/p1MYV/xSUEt
DfU6yqWYf4xxssE/RZDubDQnScurkyzVPh3e+EavD9ajIeog3NjqdB/t+ky+vw/Fqwf0y228a36j
XXwkxbvweDpAtogWrOv1Do74HK56WSALXlPKC9D8TmuUmo5ZgH2zC4GilYM37gFPxl8fkKgpidsQ
D82qWEXhjwhng4EneADENMNzUs57T0ZyoRMJwJXiZbYEq3Ns/1HIx9B8THVNUcnA3554MwPG589D
70K/gtIPhgVOGjkU2xiE9P9uzNMz+4b8XVdkwTNzQXE+NU6PepnYqkILi90uJRt4aIVIWzQzh3YD
F3l0kGwOYBXbSyKEeiW1kEQAhcVtaVcnMXgUSla6LkEXnrHEvWMyTK8OBBoNagf16+eGRK0VZJIh
u3Iho8lOC19CE9Y2dBa19i/rahkeE6kw7XXu1XJyI1YLWK1MyLwpxSLWdCMVT4itC9Bd5DEzpXr8
jXBHV5uaOReEtdnmQqIcOKw9hhF+XFtntFrI6IhhKd8sSYKZZI4GMzHY60vcqyg7PZQik1z8adKK
WTwXLxuchoGqIYmHUFEVUvgvFFdO8EPmvWnsQWYNJ988ARZ1kZeVe4gncny/1FcZvSRopWGTJmj7
Hm3hs5HpRmIgRWAEFvbTIl9LDGPln3nO0AaRF9wwMRmtWXrmabSbpM06ssgrg4HhEF5DRb1jhahm
H6LOSP4cF0ecGGDPmROxE9+VBPp7j9sVjD0Y6UQTvS6cLTW9O4LehtPiS9kUQKLpXpaNvszhtM4M
sSBnAt+jYSSRWjFrIfwGyj1EjQ5+r4BCWBU8WJ9BxXk/WmRhygmvkxiOb8Xo4A0Nsk0SDd4zggGV
vbCVzyeXGoC6RPy1K8p/sLljAS0UEQjP2Eo5fJEZ7QUPGCddsntlDlt+vJfbPsOQsyM5wIAWI1O5
MpR9nx/Ra/r+KUEVHcrmfWcj2kxtNh9NnkBS1bhFRtLxdoUXLrntA4sm/v96ZfbbHZwVkplzLte0
YrPc7KXc0CBH0q2Ri4beGMDDR4+knzbcHF9sOB/g693qqKQA6IMTTckv6AVVP6+ehQmfJ4RG/Q0N
gGr2wwLmbPb2B4/kmOZy0XiWzecOEXIHe++iIIOidskmaQJrdvcnOTARsKlU+X+VAt6GDqdY4pkP
8WJnxJYwCtlIzSXngXNqGmZK/8V40xs/rHU2Do6y3HSDP7NWogbdsNyo+4y3KeGTQksOzUTllGWm
riMAT6WgZAxLS5ojYRbnDUtYag7h4Ig2Zt0RCH975CoHF/lIRoE1kqTJ0j2MefbcoEfSoZT/0H2R
9evBSsJt6ZVBo4xoY/DbYAB8qaHbrIHSc+3d0/oUOx1uu9Y5LnExmakfa4YVZMYf7/vp6lwF0hL+
gbO9wM17OG8D57cXHfnOYjPnD3rEkUj0rcdvIFy/zMwNms3N5fO5rcGPw9gcgO0ChfoY4H1tN7yP
2/Ffug8pYbGe1UdTwSpgaz0F+bGDO6wIbiAIHGf0otjrspoTsAlE5h8F1AaYVyzVaO7h0+sLWUqa
zIIikyqgEHJLJIsOqlj5qxx7TAnaOg1k6v8U/Hpqb3CPAl6uS02H90MDGeajohRaGCYTMtZJDExi
VOvqmkTtV5Nf+M0v6E+h699u8D5m99Sx2CqKjtTSEX0MIC/VTJEBIa6uKM3QUb3ZNj09v/K3MFHB
gDFmPF/Xl+xNq8Xw/DK6Zs56JeZBFG3c396wGtfM5laeZ6VnaNlFVO3js+kluG6OgMVvzQ0mHC0X
/WSPV0etl6aCN28xolEhKg6AIiWpubEQk21KA8KbKtu8PGUMSV32+ekw9D+x+FmBmDjpp5LIZe9C
6k5ynCbAXiP/O/bpxDGblQX0XtYkiw03dlscgvi7HhgIK1tnX1N22zNTS0vv8TLUhwYtJhwadb/c
+A/Y9zGFlSN2cv77Vw10B0W5igjiG+eKDEORH3Orz9sW/68pginh8Dx64Var4pb39NzHHlTa1Ai9
2KyNOaBdayaOZPy9Vbhtm11MPKhZ6o2gpYCFa6lkg5DpTmNLwAH4vECt3EzgTwpdU3M+g6YSXS27
0jdJZumm0kBytmn/0raU0hQ4E95/FLFn8FQAUS/1T3b7goYLbxHO0ja57JDq9X/c4kCJT8VZWk/I
YUMZrcitwWGSKcugR+qYV4MPqK0UGA6ha/Gg8mjsJ0mbe6og4MGCDkrFzmDJ/8rmYrsKbcXiOD3g
SE+4eYNQ3ULNe1/ODvHgjqlp+FCdOsg05Kc6MXvHF9Rynyt3kZIg2445tUfOKnDVknbeXlVyIJn7
c7NE+MVekIzF9NCkoKUohmQ+KtnNYhR1ve2PGUQ6cI7Blre3iKjH2Ft+6UVWKtimtSxGfP2Wkhze
Cpue5bDNDYj+gx1N6Dql7RGR3QZKFiPOD/Gsw/BiYXX7IZk7n65u0HuMsiamM/LOocz2l9k0qGpj
6QQHZfGSN+OjNMN9u3L1IvhFrXsaIEKKjUN0L7zyGjOCDu6ocYv+B8rZn8A4DwiZBNTG4d0Gr26/
nmLP5FTBxZ5EpoXPdgxiF5ISVIhUH+2CVMUj3h3WMSWRdtYE6+kr/NyA20JQ1l8AwwYahSdGMt4j
H3c485egnp6AsTRTqo+5M0A/ETKuDv5Ko+kBbbcEPLwbPfoEqmoFpPcr6IOFbwbGXj5WlesyVEMA
nm7pyQwlAHOwziIeBNsl5DEBxWT2o+I+GFmFrTjnmMLTmxwTok5HPyBmTPq+U2Y5aeKeB0ZUquM5
fAuDyfWuhlfBsPp+dptwYdvDjIuZtUXwqDeCzgIOcoA9hp3UDRjh+UAIyLUTDUs6+bMuih3kAy4B
aPl1CywvCMhnHj0us6g+XFLMq04Z2E/HrwFzdZiFMFdNkbcMOEyqx65hZf2HKQEOnMpj/2WfWGoS
Dpqi4QfenKHKXubbLk3zeOvWx2kugT12QRX8zJ6Vta7F7am/8cTl+5Fit8WZo2lsVS5/pGJcX2yk
5kX/oXgYvoFvS3Uno6Fmo8VSYrRPQUD4eI5OomVbZNaFccqcRIy1VDsjp7c2ahyVA4LPihvR2TYQ
NRu8ikNqSMCrM2U7+KlJFOjl0Td+RzTGQ6NfpwZYxCQhVSsyprv9tDIUguiAW/s4XCZpEHO3pu/3
j2F7t/WpsWg5wIt7SuvpRCKKafbAxOVVoyvL6ToYnu7Fl3QTx77wVppx/HBOdsbARiaeeH34YOv9
4OzX/mnAPiuOsaGTbtJVAV83axXB2DQHiqfSL5o57T7JyyZ8Ka1qk7zFyZ4LigkT5JuqZYdByGYM
T5CcVKobW3SlI4OVFfDZ5q7Mr0CqAIx4WDoT+sPpQjMqWqA1ul5FmQ5/pmXJoA1/Q2F2Uz4yjLCD
FEeomYIgZkSjJ6zjbjkcEWXvHB2PC7ZPUFuKImfh1vSxYgUd1UbPySD557p5UJPlzHJUbvVlodVk
EKQurx47qRr+lhXvXDrRLfmN/zb01PAA1KG4hrTBjzlE9MgmYPQ38g+/wIggfdUTsM7PFIKojweB
0cGIN6wsC0mYxbndJyvmMExhw0hdqsSt/pjU+/hLroELtWlAUaFDGldTSSMGog5a7FiorvyG4A6Q
CfUmGKOEj6DXwc2wFLz8MAcX03gWPu6QFtSPnYPCFOYCMfCaj9qCeeuKr+PmHU2JWItBRzPyAbek
B5umXXMZj4mgYElkpFjxUtUO94JmzQVVSWrKnVqeAEC1zs+OxiRCwepEQKZLEAJ+hUBjKl2KsiEO
1YXwW0UUSnsU7PPTP2rEJNdK7HIetoNlaQlkZIFIBsAcTejBamqUbrZ/dO5+xCParQbXc9wJ4aBK
y2lP8GNDz8Fce8DceQ2K2UEgVA3LyJNI0TRjrWKGmEELTeGH8t1o36dyyTV+V5CKqTm8dTeKE88L
Gcjsl8j0EqY+9y3AAh2c9qMqOBmcPwl2osxQzV2PAUYXACBynFunjcbm2xflXvDzueAnbHxxo4Zo
yW7QkuZiTcQqqXdZLaNAgSrqxrQjLPT24GTVhcPpbKI3jMcbmrU/bsX1KC1vtb88HIDstsKBaN3Q
5Ql2l79mtU0+fDhGXEynmBFNe4bKn/WZUGzLp3GpYMVraZuvNf8MKdP/9P+fhNKkx2BdBuxt8Lt0
jifKYEDxxMzib0bgLFM6K1XOfXQK9woi2babO/J49TUAwAzC91pffWEG8rx8/i1skhYIEyBDoNsg
YnbvOaw7pnkOK/IHJZEDQViau4+SpTapso6u7QdMPEZFC5FWdqicX9t1Ixlzbl9RzfEPHhS/ol6b
fq2DdT9io3zmiBZBhwVjcCmtmZXdrA0i6rKL593MSQqP/MtOuGdQLLTw96oqZffzqAVBiSLF4bEL
NFZ9aQfuGSQ+4KdJAw213F7Ys4lAHysX94Zx/a2S98rlLjkz6IE70gCKMoN2QAWf7kcZsoKfaDk9
nB2chsrcyldXpIYQhuaGcr5OO6/FCWmoSwvgJPO2AlO8i7lQBszoCwplP5NO0RUUeV0qeI2yKBlK
7wIEkPyhcaONhQB1IAVEE7MOWcIY1p6BY233l+J2Q/YYgBnN77Fhnc6EQxz4rAxlg5VPpNp5PuF8
u/LXP/hg3cfHq5GIFyF5IXl4vR0kpmq8mzTN5JxeS3IWRvQyTbsc7Jwpnga7NdfUnOWgOKe5wvQu
QJ2Bl3pi17ksCIDkAQKg52i95uBB1wOGhhOVNCykkgv+vbPpqu4mXsmj0loT3L/Tog1lJ/YDLq+3
aiKyQWEfz0t9ZhD3DkkYN8j4Z2Zd0UWbqtvQdLbm2lTD5KrXsQSMDGSybeGsGKTSOKBoi7Stx073
ZYPnc2NirrJJ81E5pBj++v/QoGtIPn5HuLfCkfLPeuU4chzq0tQt8jH7JiPsdLI3s0UJ2AiWQR9U
9XOKX9n52rbiX/MYd9he5hXe07/PtV/eHi4nLWm+NsAdktjU8qO8JCNiTec2RC881p+cXET/3YoJ
DDa+H0Yk4PtVvHycodwooGX3dUlsuLJ1G4U0YqqRp3860cMsleX8JHeVUfpaR27E437+y7rzlCv0
PY72wJ3XUoJGDD8Sv5LzaNdMWahuRcO4sPW/e8CRS+hcdn8yrW7QINKpmdGKLnLnxIu//ZQ3UIgc
PHPlHMoRAuMteITSaxCdsLFLMEN9+VKoUp3Z/7d0blUxBjlupsXSZHxd6L/1paai5fr+rUsHDau7
7V61/h5kngS5AzMulE624K67pPaUPwKFdJNXiZvF8NXE/LvnNVzKc/G4ZPwI/w5tGwbp+6ieAumW
irOARwd9u+uDmce/5VLwqxq1LqhauyGxBB1sZdhzFuLMS8sQOByCtrOtGUsWvdg30ckTS/LMH/Gr
kZ+TGa8hfjKYA+4oZvFDXJ+rv9/1UFJ0RRSaqLlq2ul821iAczsuSx6Hl3riAhzzrF+dLfWaLJe+
HY/vZhtoUPZlDMO4mYibhIwA95BS9t38/9hlYdXcNiRZT27zPKA5v2lJajy+sqklBMV19dQListN
xJcCqqJvlY6JvoETw+SijH475JpfwrIwz28EuI7ylk8+xwTEMpWYmvNp/8aD0zZBaU5pBr9m0okE
HsN+Fxzk/I3RKeSWCFvMgdnKEjreNtLEPeKayNJoRFsQelidjRttFLgEI1qhMw2V/Z3rcnv3rKiB
/sSsuREpcpC9sf4vRQJaXo4iMAs2Vkiz6RFYvcNfiGdKjIBUEByUMCzX5n8D5r2IHLcqhqEmFXm2
5cr9Idch4dkS8kTBRK5zGlRRR6HAgccRUE9YvMDSGGxUtl5WIsFsKj624SFtsUgEgyyBHTpZxcUJ
38sf0Ej/ca8Y5RBrbqh9fm17wi6QJe1Knr7xtLSfJF3dngsAIVtPtG1eGkuaoZlezWXEyq9FPHza
Udo9QDCr6frw2a3HcydV8bRDSa4ma0DmOJv437jKcq+Z0NXMj6ie8LR/cjMs6oNsznlhacjX2zVh
6uAzTbSVrP1EAnZgmFQjdK4CbX9DHQnmmxvmJebgIsB1vvhOW/DjEWdgbt/9YbSWjZ7wbkG+jmIp
GPqhGNXJ2Gv0tiVzQH1Vw+bJpWNNEnzecaaLJYfEDL+QowYiJu5bqmxxu/V/IbiZPhME2irIoM78
A8vNYugCunlxWNtX3boo3tL5gbN1kn50GB5S22F2XT4HkToflWO2c4kHw+RlhWEwFsrBXo+o+lH0
gFFsgbS6Dg3aWdnXMhvUj8BtX8LnOXpk1uC0ZUq22EBjPtBt9TzsXe27RzLXmTOdZKiNO2r5COHQ
lHylNW5itwmpvgODhFjGTVr4eSX8aV0wYZlgd0rh59NvXVpxDSfazWASXi46VGekbxiEppv7Tj/L
6eELWAh4dmMMNODacOGERRUJs3aIiOXbWnZrmqmReb/PLf5mcEfu7D5fdhbawRu1pg2LPGQaT5cG
EdObpqshgNxOYPvvPro9caLTN8fHLuF4gTY1q8M6qnMIZ6NKWS7SEZsM7n9XfbZnbAU9WP2bvYX0
ZYvsICElnAh+qaU33Fd3Gt2CY7avT342nzeAUN5flDR6oL3mR1v8dzH4noln4J5AAuMa4rEziVUo
N3sE6EKEVfKuvl/66pXYodQD7ygUGMDwK9ahv2Nvvgf7eMqJcG1BLddloQmz+MFE6uG8GwPvH14p
lGmnsSd/A+AY3HOVNcXMbhQ2xQSOIzjm2bK2ogQmeY/J2gfgi7Leh6djvV3FrpBkiTSp/WoJwddq
rm/+fZOLcqFQyU/Iu2mfJSpmvrAi0uF3FgtoCncGFbmd4VGazMyYg7pWxI3msjumnY4NMRCt/eYX
rgykYPsGTPmiWZPqoPUOShXFrZyeOh6WljPY86qQ8gk3PKDkrbTokrP7Eg29Cqc6xIAG/O5avN0b
JmETBIKVFr9++QffeULtk38Dl5sJeX6/zeNY7xJ8bFephpc6O+XPZFdc5mTIty1dRiYN0ULIRtEy
oBYSrwxAzKKicr/DSITzgdwet4KiC7MbGI5iT7K5AratpMF4jJTTe3G7ip6kKrIfzgM9vqxwz1xu
jXbF/x1Ay9h9Sc5jdBNa3FAh5IFP74iEVF+4DyFnBUzePObKO0CSvw80QE12o5C0KuZzDuEhx76x
XLnmLIW2bsC0RVd775jP9e9T3Rr1Q5iSf8aZL5qeIgp5ZWUGzOkwF1iw2FN7atFTHcnc/9nXIDRL
PdYJD58S0Yauka+2c00kYWO9hx+aN6vZqfi3v1MDfXen9l9nD5H2OQJYwVtOVkTa06Pn4B5fr/fT
/GpqbAZYDBGWwbVkKphH6A1jfwcgY6hMvlCxSZLhC7OgM2yR8jSlzra64Y2qsEu6Bbsl3NaPg0QM
DTActpH2+G6urKLmpTiWGyc2/Ot1nNtVtLion3BMzTJ4xIjdRPy9UzaPn/es/ZhBLUTABD0Wrsw6
rHQ5cEz6qVX/qGif+TbYbcCXE7jnF8xTDG5N0jyQRcp0zGqHkGsAR5iQRfui6fqTqa/DXoHsbzcx
4NO9pf1ulw3kk6PFzFB5As6Epjg7brFAfnR6NejXqGpstx/cpll7hFPLsvWaov/vZAtLgJpj3322
WPGuskkBpTxEpKfYgzIr6sFWsy2kRJF0ZkFuooaPmYhdrqNZxfsXtW3ybMsyTp2x14f5DwTFkrQ7
gmIRN7kuLre5J0YBnzB9K1S71ZnTj1NoInSUwhYAaYLMQ0oKB+KqZP0PVYmTYEcV6XIMeUhk54k/
FQ9O2jNHelGQzk/vIc/dEOFLZLjFNWdLj6Y/f9pX38LAxpYM2gVo+S5RB6WGq/GlTzu9Auecmh1J
yOGhDVGf+5FZqfSmj0KMaaxe2MevR/xXOpZKojLzC22k+1OPvIwdg8d8NBo8t8yoDbMl9HtAVy1W
6Jbr2DTHg5O+rPYOJZ4179Jh34z1xyeSeRd/zVmh8yol63/3XCP21lREpFs7hUyi0Om2JNgZerDg
sMyxIV+drpYboquHOcDTht5xQxU/xPvD6Xh/VSEig3A3xt8fIojI0Ilhdfy42IkJG/tEvcHDbRvc
Cn4H+pWF2PB9ipN6qTPgqBAcnhZasQV4cjiaY3/21oAf8tZ393krxRZaXPiTxCmsIxg15OEpMM30
FntqUNVgeBU+H1yjAd2BLFRMvI0scIrOO1WmlmgvWC/15tRWgGYh28fWteKVVW/2cbWgyN+ovdNA
5oRudfaN3bbV6PTdTdNZcYqVLK4DmjpN9XV5Yd04QgabTYQM3ZgldU6XeVrizP4TZhEsMD4auvsw
xwlkMhk6pX1G+6fGXoV2es+TkcoUFEJE3sUsPxBQjI4j5XbV4cd0hgxA/siUJMebuWioZa2ibzzg
/InN3H9VfFnNvPTa6jbW95zOOJ7EipaE0/Le8SWe8pFnlgHVk7iyZzqPThh3wTd/MJpYYEWlqISF
Y4/s8q/RMwhWmc4zpjgqW9jkD/Dgwr1r6gGoU3ZUsNQ2M94bWN+Q3pOue1CtrTu59pEt8OtOUVL/
5ymbS8Jc4d5GSKMeQt5G2rnJRVtabMMFvooInbzGrojUU+DB7mcOlvKg59XHKJ+AbLcz/wVzyOQc
QC0GDYTuEZ5d9mAOH8GysGw5v8Iz9TihzBQymuum6h6p8wHwPC28pdxmH7Rwo2UAtclaR+F15NSu
O1usdv5RlU3XEwm1YgWWYg/KUEED+W09HpbHlfmqX2PMEOblOTLOlTy8wc4PLq86HNVU6jQ9kIqu
Mx6CjNYw9/XzurwUSt5AxE4LbjlzUTAueWjNFzOCy9X7WGICBLwH/6FlFiEMjzCgcMEI660od5+x
mgg7sMSXhcO+lsmKGDqs+TrcqSMryt7UVxISql6p83ToVDTjjmw+YLjzjWC3twfPzlGCj0jZepmY
nccrPL53zmLqObANjD8uNYrHZpiOYVbfGZiK16CxJVnJvUystGVuB8iF0ibK8X5N+vnE9xA5YHg1
CUk+i6Y437WjU5dS8CI1uBUuEVtysxBTnbgQlYN0wRTreXssK900njsgD26nzEG3vydddwofIzAB
tTsXNzib3GTfhVilfj5M5rsLDbrKVr8ChwksNcJSP8M91svjm+BIAfJyMUBQNepoPZYQ1zL3YlEf
ZHaIZELUBeBaobIDA+00CLpa4Ov3kzl2IYaoVLDg6YXhXalJom8Jyhz1LN5A54D2lBxcrbgwGejR
gY+Ui1pJYSqL+lpPhSsd7gXe9x58mn5FD3a0dsKM3qRq9Wga3xLWIwIhde718hbAgF9XB0B0SKEs
BvW0xWgqUJ+Cjbec+XMnncdlD4+rm0bL2oTRAE/UW2VzNS5rH5BKawltwMSra6N+CHhksabrE0u0
utRTp1VFaicPX9oNiIJF4M3d7+3JsGjo+EP5swUoz3VshUsFeo4jG5UQ3iw1/6IjVCA/mBJ/ayOJ
WNmEvE/+hCQHxW0lKds8eMIgP26oH5L9ZrLDsCVJO+UaCC6V6JRzhE+mdVvEw3ulrlw0EA12J53Z
LSXByZ9oFpj3NHFj0PGSJo/T/3IjQCsejo5V7Zbp2yJ9P7pSrESV+KNH7HlRL/Ebriyh51IrvztF
ZVDTMKX5gG8moCvRC+zQHVVR1sEfVUzm1QO2JIdAsMQKJMd5mFuo7awlZXwI8dLJ77PH7ms8hBn9
SRg3sac4EWYLlhP1VYoebKeSa9cNyc7DBWfQvtx+q+0KeSIB7WEt1ArfLEnbxwk6t11F8UOmwZ9f
wl/VUD9dSONg1If0ehwLw2LQ7XrXxJcoOxg9vxJktSbNWjLd5hSjuDfMuQrMctMcNSH2lN9FBtFx
iP0I8EO+y38YDres11wpBlMcVQ15qUZJZOBWYdYASW6C+mnIrdGYxSEimpQdHCX8k8ighumUxgK2
I+8bPcz/hAgSwZovLdpOUHsLLRtlGXp0TK6W9JGauLY+WsEnifuWZBeN23DJcbObOUCnVK4IxDcL
iwFPakO7eZbVlAZd4cikwovt4zSVHasM/rBiuOwhpRW0hqkP9G3/EQLFZmbYyI1Mq2BM+u7E6FHM
TQf26nKa4qKpw2dLKsTPxetWxe17owlT+3+oNaTurGP5cvBUSDCNY1ygTcr4B5lIzCcpNgotPbWk
e6IlRcppGeOTqkTDLMBuByPisIsP7cEaoIU3pnZAz0fmfu+Dz7pqERJJRs8BAqZHXsXWcNrUPFiB
FWlLxiU1arGzNImFLsaAK24oYqtNyAVQ+uvWHG/PobO3G8FV4gN0vaOYMVwEbCU18BZe1Wgz4sdC
7UJQq4dWWBuksGz+YS2rE4wAn2WaDdaL/H5heWudE0angPylKWcQMG0QQNAFriBp9fu8Y5c6EWP9
v+pnUuTKl0/BoSsk01ShHkAT0AtO2YJTg73pbrQF9aE3rGGYJYgzQqKKto2ImgCXoR4Be3izfyqE
8NEBiEY+0eMaxMF6ZxFIaXZxomoIDY8fy+/SeXNiTtrUqFtIgnc/pCFblv38HT9JzioIa2gUjkY1
b8hLJ0+R90/WAqyZFNW0gCdzauJ7ekBbnVW0zQpamtPQyMSZZi68W/TtVMee53Ep6VM/lRX3t6pU
XGTVUGL6crBjU2RRq8jaOJ0+1ibs8+5E4ofIIsuhwWGqKx7uFZMis0wPB/OeC1DhjVbyrWK5UIv9
hJq/pseoGT8kE+cIdC3gxOZtU2siuMU2s/4e/LiJ4QgcpgSBSnGEBGVaJz15Gal1W2I18AwJ1IHE
n2hREQtoWttk8/whuVbAkkxgH9pCcLUi3FNDvq2/ql1qBfVtUCLxopKzllMWan+Q+objkHDTM5cc
/aOMwOW3uaMH8GVQBwR9R9FLZdGEUX9Qg/XQ+FGPqt8oKwsh7PC3avz0FJTMPn+L7BONT0fIziYA
0Rw52t41c6I1mAAzad+VbOJq3Krg6ofWvIr/P04mCRlCXcEydeTWUa+dkpbzhljW9vkdV4lyVZdB
IC3yXbhDRJ7heAduT3XFcrDUzQeaJcp7WZkzt5wL4mRLqYD3fuKse1GcgMZLLLY4Qq56gWCsZ0Sj
bbQNxk7i6xSNQjWTbS+ep8Ls4HAToB7hBN/mbg/zkgOcYKhfYGuk4rzvbZl2WUhblrHmX5+FSugU
A5SKPs4+rleXv150efX/va/qof76yK/Tqr0thWbzrSYRb7gnhU6HoYsHvgLK7pAcWIqg1A/G4DqJ
j9YOYaqAxqp6h23x1rttj537SJXGhIoGqRWwCMpbGCSOpeD9/Sy6FZT79GapNpIBikEA1iik84Ip
FGMgJ2inilXEv0F0HEbFWKLOo+U8su+PBYeh6Fspg/q9DUEHkxkAfbrhanwl5k6myOHaBOsguS/2
xBDgSE5xM4VPf3MX461tvo9eZ6zeZJFD9YiQKq59rBd1tJ4/PSaXNj67fOPK/8CMcNh+ZPvYQS3v
aIAqNCQA45mV/botb92Y33qrv2Nsu2jcyo3wWZy9iXg7CyLw+5oKSQp93Sl29fSLPKQspiNEEESS
fQVGXrMlCqw+FKAHMIobpugpPkgI5yy51JW8jdwplhofixKj4meZAYwRBawI2hJ3ULyn9mN9hfv5
8RdLQExyKgBISqk1diQqvvlj9IXnXI1xIbPzrMyvNJgH8yB50VYPFuLKLFUtBm0aF0kGq8pbvBai
l5hrgu0FofALKXHYjwlht36UlKRYKPOJabQaZPCXvVsCatwwB6ioovnj2m8t2t24Jc/PF6RKUKNG
f1qDxMSM90VvI5W3lMZuz7P4Bf4eimmxljkFKeZT184Nldr/qw0lvn8KxZWYRJGNbZdUWdQea5mz
gt//ofPr3tcD9q8p3AuCgP+VTJ9S5B5nORJQ5s6AIwrDL9OX8o6n4KRShnRhA4jyBZHNnsoak2a4
+BFy2bTAv7XaCEbVpi13xv/C0nm/TBiMLUHcJXGo9gJzIllfC4tDBgzuHTCviv16DBlfzGbbcRUz
xgytu8kSqOhj9YAxLiy2jmX77pOft+qGdic/3TeDtX7G0TW4vlWMx/UynH3iLaZ4MCk1/s9ZYYH8
X13Hd+ueO4v/eg7kxIBaM3v8RZTDnTiCZMpIajuyZaEWlMNnW+K75k68Pq6oQcDeYEroYjaMuCmA
oyxOUM44if6mMh7hCbhcfhWC/a8UyKsKN1LaKpGdceFI3H5FaxR7hKKHp0YgRhkzVRewM97SY7RD
jGTsMlR+QvBiFryerG1PLHiRZMN5/2gYRhWGPtCltOAhbHvZDG/gLh4ZceD19f40SmoNuxv1cnRR
wuPA6YBI1ePX69TRguMdgdsgeuVg6PqSQlb/b9rlbDqZ64ie592f7W7HbSQZL8IE3yXHKG3zBOfS
OZ0lMiGoaxp96WnWgWQjxSQHMhN9WRsCZ9r9EeK6KwAQt3jvRXQ+lFw2CS+DuPqOur00+/nQpM8J
6eBSNNMr6LGVIA50VIA3WU6+UFntPT3oEvgKv/MLRGKrLB8GryOhA2la8t+sx9eqrWB4n8l27GAJ
yYVMmwRmBQdzx7M/q003CrbC16TxWngAB/6Wm9Xm/m6lGATQIkTTKy9JqMHrkfsa7pJJpZiqJEEK
IfAnIe7rwBvKRuhP0B4A+dLTvj0JVTJi5xS2JPNH3uPj2P4hyOgtNuedamsct9oIUghFugo0kMsV
v/RAQm6PN5tkSaSY4fi6lijuLlccTuixM3lo4LtMC9YBE+uMMOgyC1oCsapSQCa3Oa1s79+znOSG
pqRHQiwNrL07a1Zgmtx69OInp/pd7ps2fvjPTqeLDzD6JemeyZFM8ItyLbjbYCwjzsUlA4DMrAX+
lnbYDiZCeEsWJs7nL6j4Nx0P7xOStBdj2o/QWeYBYyjbSCYUsmEN1S/Zk4gBZqXL9r9z0SfgWtdz
cbl4ieUfYx7+joDBZH3saAwMFNs+pq431fDVmW4lja+/EyqE9vBGM/FTM6mTOn4f24Na/0hXg3eH
i2Mn3PIWjKsNoHysV26fTEk0K7vGeFCwcXOsjRxXKD+L5J9YW+XEZ/zdNIHwCnhQ5QXC/PmaunNR
rMzSD+c6hrY0qSGRs0c4/CN/CS2Ay/fRtP46GcAQlNO9ZFAq22uY0hx+D51eALtLX4+dbx5Ju9uz
I0pzCXCMhT1y8cQYKmeduoZEGNND3l1IE4IJzdFwWIHf49i7kN/e4AzI5ZPlP4fFAkFPKxmlktkS
5jqIqZa99pi7JW6kOLSptGbgxs5+ssqFtepWSrFkyck/OU/kk4UAIWYMQkWjlUjsHwS2sx2RHexS
RwDrvbiKvC8XLjPkVNndI5fYdoct4XSllv2s10MhI7sFPEEn2dU2q2jacs5++oX/bWwAlLGUXpZg
1duDMRBDkvdoE4ctZUN0nx2v5hNwy9ujqZDJIikLpVIt4Le7w5oyKItg+tRAHaSDrUGeLqK3nMch
PR+QF7il9l75Kills2rDCtaNBxL/Wxi3e5zEt/04/GNHaqYC5Pc+ZcmZOvJykPhcLyY8OBXjeUs5
2Z5RNx59WUyZjucJdRmo3kIxseFAOQPgeNJ696NBy3ruwrH5ZAT0++kjOh5L+wiBJi6uGdEUc3ux
uqHb1UF8F+B5GLWN7flgciRbH4wTZXEukxBKq/XgFrdpDgOJJEKlXCktrhO4J72PdaMhaH1Kwm76
bJ0oDIa+WWIs6xPAZA4bdIaNh8V/hbvOIebTWL0ZqQDOS1iSqvXjyeCY68dBE1W5wsVniPDyu0O+
GVsbNYv61TkWOBBxYhJHOfY4z7TD+sGt+xoqKQE5udRCVFnB8XnYuugvIse1NjDKyeJRFiBhsaWo
9W+sZphiF0HkywEhIsZwdbpHOOtauY5Tu5rCRVA0eZw7vGlSun9Msl7F2dB8kezjX1MN4vOUDoZi
CDGCY8sMiOAmNonp+frCS9mgiKBNL3PkZNqEV8TtS4g5LJEDPXSgEJd02em6r5HTB+VmhAM5P1OS
AaVauX8tI36gCX52SGl465YxXvTRBpQcnOodXs/8+rOdjI6tTNBBANdx9lIgsJVtUaDzy9U88VW8
kLlcm32NtGR67g+zhFCEwhFavHep3oyyHMbe/cfpxTcwhS9IH6PO62tGNlhdDd5fkeuZTvBprWKv
kkrwM0REfaXuAFrDTPtsD0cVXBpNq7i6gPtZr1ce5VBvMm6kXaDFGTb/E410uwVhTLmnhRSEZ65A
iim3jlOyCeiN7ZTzbUPvOsL/xIxR8b0w1pkcTy8PMoLu9/cL4U4/dvfrBytCaZDfRXsICVJg7tH2
w+KErk3Q88xVIc9tyKVy50F7gCEhcn+hIm9sjqqMylu4DT2kNacqLhh6QiYrW0PjU7okrXEs6eDQ
2dFVV5m+6JiKdeCGMexy973a31jyThi72eJBFs/avesryVnFXadUPy1zNyvOW3WT2EwZZuWRqlOZ
UsQC+2DmQi/kOzGwtnxFsGj8xohknTqx+yMvcMCc/ocx/YieSoP/HEntQEWcsrv0KTOUHMBuzl7F
9ZturtTYP+5EgNmsHQ6t8kJBjnpVDL599NFvpeqHQGz3vPLtqJLI3LpYNhRh7wZy3EXLc7yJPTCW
5NwidRqcp9/5OOLq+hBoTrCdeFirrQrbRi14wThLwYOfOBZFF3ih/1f/dP+2gGYtq8HqLcYJb4h4
pXm0c/FgTr34y4hDBNeJ0yBUFERZk+ACNWjqSfqcUmM3ov9KjNXydqcIpfQz5EQX6DuxeRzlJzw7
sZjmiMdBZ0KDZsVrMs3oLB2hvgDUKcun1d7uO3UURoGrIkBmv+3V8O8X0tpdG1wRcSTCbRyiVywH
EChBz1f+cAMdYcGoaNtuptH+NZMYjjSeUBCBbIn75A0/blSbGB4tyYwKNIIbOSP2zuHCgu94cW9v
5WbEAmD2ABW+p8sBqIHkCDYybAOkW2pP5DfTcvQlCWy8YfEeF8UiyEcKI6Uwuz4dDOIWGcZdwPAL
tsqrhsfCeQT9HIi0TpZP0q57XjXLWU5txVq4wKFmTbD10IZCl7Ivvwe7FDP2jCOBxqQv7vAoCbhw
Im1cUh87DNbxP/2xekmrF2BwBjirIbTYNmuuSY6utuqX2fVMRKLxMCoTGk5PIlbzCwceM6Gm+F0s
/TL5GQd5QE8MTQI9m2Ec9gzFmBnA7Pj/IfYhTY2qDjg7485ebzNl1MhXm5a2GQ+fvYVKyHrMfLS7
91eFskFGPFz5bQnDCDrY2xZ1IZz0qstpuXi2cA5LOoXLJlJ5vgMXqCn/P8ZpCyVI/ItVNjUpQLJJ
mGVquSTjLKm7yswqePcmQCBu4cNy3VbFftrAcX63esYAq++fwGxSG0m6TeVybzVGsG74plyKuHOc
aAvHDGMWv6GZnbLubcrmqTAkmt63uoW06xrbVbNSTY8Q8rgEgoBAsmLln36xm4q3iKVp65Xzstwr
8GvxzG1dIbRqQNJRYyMtQec2XdlZRvzezRH3vlo3UmXEXOJNh+785e2oc/pBjSs/KiuH3a2MeAI7
aQcTPTcB872bFYol68Y/cO05lMZJkLZdAxVoGthtSfosqlSxyX2B8K9uoGemh1VE4Oi75kyDoBC2
gqqpWT0fpVqD3t0XQ2DNQGHDnCA2i5VDl8xPyJVnKUJ76tWDly3XXz+zG7EcJ3VzorXXQQfsjKrl
Ajb6wpDfI9wFcuYmpbob4YadWLJ+LVZEGPJBUfeWJBHo+ebglHrcXbAX8NaxA+mUE/9GxH3anWYu
0VtA3q+75YKLnmEDkX5qQeb5qiV9ogJ0XcIwtRxNb83Vh4Ns6O/hiz0jSM2EoHh0LmI2zguzC9RR
zjzpVFe4RWwx4rifMau1C1o7MNHrRlX5PFh3BYxdsbBThiCZ1JBeRwJPuoHAVlbZZN5te7QBvyeM
1bYb/RessbtaXIZKT0B6vqZJWtB28BYuqeCAl+4m9wfZatAuWjCVvfiINd/HuQZxm3yEgTK2e/0m
xU1yWJDnWpsN7D/q+kTHx32Ifg8k2LQu3Uuntlo6qLKfgb39pA0LrA/vwdyHaJKd76kK0vdXKhaT
z8fn6s5Rls0gTt11GaiwI1/mSMgG33gQ7ivvSXvzFNWgKI1TFwlj2PPdIRknOt3ebBm3dDdzsyf7
ta7wtWifc9eq0j9drveOeSDIz+u1bEAxT+iV6s6XNsJ8D57GvbkTiszO4/uk+FWn6NY0I2v5+tYJ
WcJufSbLkJH1Ma048clbK++MdrhMR+D1BejXXMYt6ldCif0j40VsGxiofTPSD/O4cL+a3bkXEDpR
caGMYqfs1nRD3AW7MEg6Jbqo9ma9k6MPteW1sMYXQMBaFyjqFbiso9N0T/oxKpWgYJPeK9PUx5bx
8b6VUs/z9im2iEhoCbDYkYIGAvBSjSW3gYSdMQ8OhXudc3EOJ9lc/72H1yq09Fj3XlSOV/qzi4Sp
9faIy7D0Y3PMMyFcYIuFCzCq67w9j9+FDccr+5mOwQQyj1qeCwE29O8qNkl45lWXfCgFn82BSTRc
LshEHX/VL2D4Rhnx2jRDUrBOnqoUyfLqsT0KCpntY1SPs/GX2Gnf9W4Dktm/lDTAo4o+4IrBmrjd
l5Eg3DV+AVUhVOavbS66ycST0M0YA626u9+MOsbYwAbOKC9R6UYlR7gfra9pPq8E36mczz5c8CX0
5YUn6VBy4BkIwCTZEfwvvPZ2NIAM09223UO8QCS39tDzE1LouY0WZMtFMV4UYWa/xNi1z5PIINRh
y/FnIQ587E56F761LtcA/7NMp5BC1tE1fcYarE13Qk6jPx+eSbcIpXciednyzlLqgVxQDZT4+sMv
BMkLpD1XCV/16Uo/wInEaAQVuNX2eL0HaVgKxKr3Mvxo1WAthXi4wTgU/zQ58f21rlEFpBtZmu5D
1T9yrDl9QHcFTrAv6yn+mafPUbY5h6lbBol8e/v9x3aLK4XJfdF3ImTPiB2ibu7A4StdoM0oY6dk
PU2iEERngLbg7QCDBj6dxSVtzh7rcW/X/R5JtCqAu5NU+ImTyKndoxsbqWqE3PcgsQiFpAYp+N24
OYpEWe93HjnhgjKU1edMjkFcLsjY8ogKcvTt/p/CtjivoZG6NpqpYQIsT/b7NfIAf5foaViDzUyI
mM3DdV6mvewJLEJ3gVteE7oWkICFpp52srYvMb5oG052hPSqjzBSAm3IR7fvV0FeXx1EXc8yp6kb
5rK0sR75Jk9SjlSKxrHMKG6UKrlQCk1B+FDijyoAmMpy419xP/Xs22JYyapdQZemrax+xAEDBx9c
iPEZPpan+OOMpkxTJKajOD5fur8Y89t577ZRYBye1RwTfwNdJ0eRJdQFtw6GaGYfw7FzLfV+HmsY
29bDW4OdkgL0Thg/0SLNjLKfsqy55H0odHcor9euzzAEp9ddlnIbLd3EKF96Rth8bLy6UM4v8+9H
iIHxoCq7+oxA1uEXc2J5XCepHup6+q8NWgqupgOrElc2Bgl1UCzSKzJ3k/b2LkmIP0GoPOxcVmcG
V1EMvq61xdRKDANP4LGoD2eGKHSCHGyAYRSowT3/7ezKpopLe6vz5vW3R3n4UZP59uPElpPmIaUe
xYmwE8VLgjA4ctUi475oHN+somr9AZ4SC1GClF8ubn1lb7L6G+ypAGf6o9+2Y05zCylxNqlrUD3U
2dHdeE+cZ0qSDDl9E91JdpPrtl7H/C7pTLFnel0H36E8LB3GDo19mbmdY+vAwSMV7/GCXZf/2OsD
RkqiYoJX2e0WqDECblStJGAr1B3keDYTk9NOz5TyqYjRvAkmft82UiGPK+ZXS8GTn5XSGaDYizlZ
htCfBUQ99q/qKCDjqg96LX8wJV3IcplwdOSeFtPGt+sqadeM0Pa+s7EiQdbKsyAZMzlvFc7dJCKf
UF9re9hXGqpCuu8y1JtNNzTp7VYq1QLZqh6zBXoYElRbXq8UXJ8v0WKbnfoUclQzaIIM1AtfM2VX
ilVrVtY7ntZxnvuNjq2jUFs2Th4Vestb5nbzGMgRy98+vYgJXvOskkRx1UR+MakCCIHD3pLfOZ1j
p7IlmlWQOxOqXgnTIoIkpUFTauKGva6gz7jFxgTlTocdiA45/+gjNnGjE5ti7OIRqFWXhOaqjylZ
c1nAf2AKnqsHrh2D2AOHxaLWSW9IYBzfgC/aIcBqqHi6HXei3sU65wKb13+Yn9zMsgFk+CtqCiA4
jSNiXc/Kz5EkPaLBBMcMqOvWCSsjd0huldlZsV+qhZvPdmaE1Hk1zWy2pZZvE7YAMLU1aUcUDk07
1wecG9xbCyIBNrpwou32RU6cERZHdutsVs0JYzRpevLsRyV/PUVnDJfrUJ97zboO0HjDPEd4GKSg
1Yfw4rm7ujX/Kqt8hvhn9QhR+WHc3xy4Z8s/cG4Wn64VkNMpaG/d0q6+36meExeQOWEEesb5+XlA
HCicZV0+M12CkkKVEogNUXZr/20eCQvSCHHTDtggET8JUOjyYGf+R8akny1k2Zsa6NzuyaUIQwlP
urFPeOVqcF+2l6YGtDBruxIXGJdn6BMLdtKw60Vls7Z9w8cRLZ54sXtwFfaiXNMPn36dk4MX3Lx6
R/RbiswkrNLbfXGDgJsHuVNuhfjHwga86UyYciTOTAHQnRpU6aQrnws31VO3hB9gjktPBtU8iBRx
IG2YL7cCjf+ebE1jeu5vXzLznAdFPwiNx9D5TQo+zAMtEAc2YPrA/ef0Yi69jPzHJLzIUxuiAlFK
ND7U6PEDzeck5t+1uxCqL5F1AlIhxHSoa/apGL9nGIm7DzbTTzwFwrT5tSPEJ6+fpDE/raBmz9cm
5DdZ9mTKr+CFRIF+nHm9i13EvplVIGCvGFSukyzWkTAIQNxBiMuZKe6UUfEU178HlVoD9fN1oMhe
JI7BAaZbnF3Pv4xGLi0Yd2JzjH04ca755VN76sSw9jRlWoJug7DrAspWIsai4JT3gAI+nE+Mktud
BwsrAK3qn2rpMyDb50zrsIaGr0YIwRUg3S+82UzxjrWsQDgfJS8l1V7htDnjRF5DmU4Z6ksqpfTs
UYchZDCDKNM01s1onTNo0Yy+LxjhJrHlBlHeaMT31CYr8YH+CBrH1AZN4eOL58z9hjiYdpHlPjR4
RabDz0niDEz6qeegWw/6ROhJKgEhmT9LJyeKSEWzIS6jSeaCtSyaM+GrL4LF29TnJnpBubN6zjsW
ep/hVPDDA7fqvuC9c3y74JHyrxnEEguT1VNDFELRpbTRPQncJeUwNANIDbl22eRVcu3aYXUj08CW
M0HB85RTC/uv6HGeBc+VnpNY3mWE3V2L37YSWg36me+ep4tZVEnklWcxd/yMaCeR42525ijDLifU
cmdfhdn+6CyuVSKomiR7vGGUvmkn73ppDLlsXEp8fa3lk2JhmKjP/4oI2XSfpPOZQmILrJqco6on
2+AB+fpqVN2Eehb4U4mxopNqw5ygC6RIefAOuyh7Zg6fbWCT4yDoRc69uSIma3Rpl0Av+ZzwyOLa
6rlJmiIN6GQgRyWuHWQ8ajyxRpIu5bYQYMgO8HqD+l0vhjVG2ymCN1t/CxoXmJAjLalk8TPTjCwX
p9txeGtCWYUWJYko1RNhwaTgJY3YfwjCv7d+xtdHkBne4EmkY2aWnDmT+mzl81Dof5U/sUUBarbx
jDjiKMGR6jyHmq+s292Mtwqndq1DZiRojXnRY9zcTuv+gx4ASDyCSRPYUaUiEaPiqesqxaW1oOZF
y0D7aBRb64fcqpfVSfB05IFMnkzj25N/DufiJlCmelg5OWY1AUkpJGYaqT8zrPUxw5njot8XXxQT
k6YtyH7TKac6toqKiivS0AqeMldlcKZKCjMToBR7/iUtTqWkN+Qv5wXzN2lhMEHLqa7btpcxAHpP
RZu2pHNDlVwi1sKjpAV5XaF8InvHdx79Szu3WPapYYj0zuGae2YI/yl+P2qMcbCjy9SqYCKHRH3C
e8LudCpxz2Fgd2zuBGrIc4jNUkUu+VWCWgcVCvgtx/XjM4ZkJjd+J4BsveUVJoY0ONnr1+F6Mw9C
XmYuG/evdVo60XKzajgK1kAuc7mNQtkRx6SoKj5Bkax1HLY7kssvS8hN6v6H1v7JSEG6KRdpox4y
mz2vCs3R4Cl7EjyTHpgI67r213Cg4HXh7TkJuB4l+s1PNcO5VwiU+wsPaqpBz1eeEZZlkzg0IaQe
y49W9+oTNmNc1QNDVD6aMWpQpmtgMC+UZdfutEzwo0TTIN+BMXmJdtRmXm6753sKRghYcN2hkXn6
BKdhqCCG2vEgvSx4MbaYspLmoUsEfTQMFuh6S8OSxmsZUFBFseNkLqhm+dx4Os3KPaS4w10xqARx
RyYLwmkr6D/NWiA+sd7/WeLSMudi1NiYAbg9su9NFV2pRpUpSmgtIJvH20hkS7Ig7aOma9X83VRp
s8xbiwcwJQ4Y/FUVB8vGKramqq/Wpm5iJnyxm4Rhs9niJONL1TH+mKimCUZ0RH2XwLRPBoQGckzY
PjK/GzcCR/gkAXRh+A3m5wLMtYQrKvbLQNr1X5PsMVQSOAtOAXJ7CWSEohH65JzzPk6T0kWNmn0e
Eb9CxwBnOjUHJ/JBwGTddN7eLuXvyBHYvKT1fjSIKVfu811X2r9lM9/3X4NvYN3ouOY1lIBWn23S
68ny7mRQ2sx28/TW7GKnCdQKJt3D09IRNKjLQ/wyMBDioJkN7gGJot3YIE2BEtuYh44SicoODPg7
XOhNR+XIH49O/Wb6q4ZpKb7whBzpK5zr9NaF18Q6kH4pZT8pn8FXEcmbIz76jNK7L2Bxyfci3bix
NRgNLmPopxC4c50R9TePQS0i0gyDnyfVH9kvooXInmbLnkwytQ9jDSzL1IGuqFLeMXFWqVRf2E34
jlV4RSuZ9R/cKoJ3UhD8t+GTgn93FGV0R00BFIxJAf4EBoH4SwvnWM6tSVCIpKARzOyNR5yPf7dY
uSxWBF8bodIlpbGNiOe/NFHgznJtnpHCCtOnTNmwCL3RmO9j8f06IkwBunzsBpB477GvMprlLcIi
TtKZJkt18BRir1WPofSKvnNjyyEwlCoMpSp+iLut1ipvuRWYqOTvk85mc7efgBg04zKaxuWrS0t5
n/xw3+Kvdsslk8e+bUzw5OxPdwcSYULF4tcq+KJpmolcF+85FaJoAeKdl61rJZ89nsiwGnccfbcM
07FyViM4sRrBPqiSCgXdABVpjGYfR1QKE0mQhVhNqVrusu2kCK2ZDQAfJQ0IX4HZLNt6Vy7mAcO9
7+MrpbTEquxLzxCrVOBauKkxHhndkjr2gYjG8aO2xji0EZkZYqDfjOGXhv1LDFf5oUvgKDx/W5sT
n73GsK3yj009ALh9iwL9catHRUPa+gmSpWO5K9IV4oZCGk7a91IL+QAMZaqzzvtRaTrp8BrNjB7l
5WIMpsAI7xCZc/q79Dgmp4sTO9ZugnfmPJIIbKJkL5G7vahDIxXY6WEtm2wxx4C4Tww/Wu+XFNZD
1p8IgwPpOPty8OWP1kp+C2Proh5uZT/jKLuXY3Q3VFGU0hT19qiU+Nj9azwZMLulD3U7IjdBwtAG
tb+6R6DVu7fBRKQMVQndlScQJUFwhS44ZjOalITH0fjjwgwfBF2fI0t/7D4gDa2nnK4r0aeHVxv9
N1OTQnUuDlRi6v2+58OcVIdrCFDOv09tdNX1O/iwNVc+aabikfQvPPovPoRF9WOHcJgqbtALR9Mj
bOygYN6m2uDkETP7vvUQwuK53trnQ/MEA2Amryv6razaJgvFSA2EFeROp1J1SSIHLkz0X9dwkz8g
VcLWJ908u3dvwRi3C87S8E1ByET2+iv01aAToTM2kReoYjwsAjqcLasJkck/g2lIeXB34P1Rb2Ic
aYMwY8G2raf8vftV3bM/r2f1Wji4R1A/7EdCADgQGeqD3vLR9EXXv4t5WB4qD6c1z91yFwUJUEu9
ORtIQNpv2vHd2+5S+EnEmXLJa11ykeM6YpSondMm4a+/wUZ7mwTVkQTM/301/8pqqz6E6KT0a7dv
qjwebJmw1YQSOmTePFmn0TTA0jOEIUS6YaG8D7clXg3QijVf/LkYxG6J9pD3rzr2PsO3EnVdrReF
UolScwqSV4CCHVHUcR4iY5pIhiI1aVDS7pG/J+d2BnpWs59E4iyggxGbwg5ao58iZo/5RjFfz4K3
a8tCQcwch3bZFnNewBlp82gviUGsZnd2exrgW7BYdfWcD3iH4tTItWLUh4phMM6WQrXNkUvgjRh3
1RtxATheW6c/j78pIra7iRAfosf6JpRTo1lJg6gSFU1vEYZpanKq8xrB/+U+Ys+/sn2Bg9+oXbU8
6qRWxOSSSSdo6kSZH7A/wi+ST6Csk6lQhIJDfzyK1G90kpXMjqUL7fSsFVDjps/gTo5WaeFwGo2C
OuK0XCM6ROw1gc/ZZR/AAreoLXiThH9/qAtjr0Dnujn4h5xXmzx2WYoguHxe9XXKbPWl+9x1dR1i
456OgsCYGSCh+V0UZc5sYCVwo94b06HF/eqhamkF9sm6G1AdO4tSD7a7KyRKII6xsBZcYtnE8CVc
2bHxbKjDRe5iqmAe/wvLwnbkz50px97EaowzQRA3upZ9EyklKUxE7BafiRqztAjTOX3HQY1nXLug
vaSz6bJfZSUUBCWBp4dR0bp1YTPkT6RofCeawkwRAMz84wBrkKIaI1f4SSevgNH2wbQA1JTh3sjI
hLrHZs+tversTCj2SoIiQR1KHapR8P7EzKDwpcC8DUyjLaV36c4XLAYuufEFa1P89ABl/a3FpRaq
PiF+8BGmSRJf4I/1e3nE7IfC2dXdGKWosSTloOpYnLAR9ONRNo+pI9O2Le4n86ZfVg8TFAEzRuS9
/VCmnJZMvj+VebkrDCjPPxIpsDGS/zJ1QMlg3t854AVWf4Smo3eQqGHUdUEGNVfv1Y0Ntvy2fPhH
VTkely2Flg2g/da0ow/eqjS6HFBD7synrS/JKCg42TbqwiJjRPOcM1JuTdyxHJ2MGBnPv5Fprcgq
A4hXK3ylDy1F77mLazX1K3wKbOdG9m4ouv77QPwL/LLqieVQkZpcFFnY3DINPF1+rOl81KeeqPNQ
I9j9YdAdzy4VC6wti8OadIt5xeg4Dzf5JRyShRl7GM8y8VUR774ehsNjPOfKI9pNGL7VNzFhGEjv
ceidsFj1WwOL6JnpdBDw1UKiQAL5C+aApLd+GPTcoyanZ/hPG03k1QxRzhLvrmdcp6hje5wc1Ry3
dZAcuYxLzF66WbkS7eosCmX10tsGlGAz7oKmG7SWGKEYAb8+JjHu2vchzuQ/m0Mj0kcE0cywcXz9
zjs04cYKFDvY1bNhtOtIWaPnPF6O9qYpV61LSZB/kWpr9D1Xd4EDBtGdwVT6dnyRedIhIV0jUIiB
1+ir3Or5Hgl0muOdyoqV4yIj7EKyCMC8dIV/TYoEEpWllj9HGLfZRQuvcc1W1rAMtv1QaZm5sbH9
TZKs1S6gSD2PYGZhl91EdsYz0y6TXwTcwj2jM3aW43BzN3EHMBGJbQ9q1kagM84lruBVrFUyKorJ
IfCD8WqcjC295DF5pU3qzSCBp95qPDDBw9G2XthI3tBZki1kaUVynmfcqPXuu7NQ9OqQEyWdN0lm
1MHlXG0TuMA/Z4EB509DGbqWfqIVhSrMeKHYQn4BxHnsqcp/lL1Ftwcy9AGN3K64e4wGUp6yufDU
+i2epR6IjnAmtW0a3QR8behOarAe5fXCwtgkeYlUMqYrP+QdlltXkTNLzQ/Nk9z3RkUDg3L7vUFt
cIDJ+WgdXJwnNQRIS47FBICJ1aSKPQpioFD7QOMkXvDbi8Mn3w57HhH3w6bu4SSDpHc6a4wGPenN
r54LzoGGO07bHTJxbetEIKXM9ZN5M970BXKlc1ZU8e0Gjh8rSAMsc0HqadCs4/PrTTRliCPB9rLV
WozoNybzxfqfA7PzC6GGfLSBaG7mTrRCq3quoeOYdu+217GPyMGclbefuqUJyzlv35uAk7ogndHw
OQ4ykJA5vqYYKnKpqEZz2x6DEEPYzqgaQDGPW1Rn+zx5DBnseArq5lOM3SfcIuOGqeWza5vLG4WB
HhNem/WbrPusfWcR7P+rGxtisMK+7kYM30qnJNZZQ93voI9WSRVnN8WRlE/czTvVxP7DxG4AEnbi
P0byYxg1Aqzzk4ulQZRVo8j5ISxMwP2SxAHn7hE7IuJrvRWK+P6oD7JIR7eqIRv9+oyW/m/OWX+6
wS7rdPzFtCH/CdQioRaEIiiUtWoDSBdGPrV69kZ+ttWrKegXc3/fbOxLatYNUSPAzrgn6tSsV7Uk
dec50/5dYR49zElA1/PntSW13zBjj7yX9k+iZnfhL+cpn6nXLAV03Ue90skTXB1qjIJOC6oTxd2r
nanQFwoGZi/UQfLMh9dRN7gSXfXM9J3WpD2sCuqAq0LrfE565QbQFzKHahhtYb/ltykvTefB1hI/
Sj2pZYGYWWQuWUe3/+xeRMlBh+Dqe01jy15QG78GR+euzjGBjd9qClW5SInPM8wY8vL9quTPtv5y
P/XGx8so4BeonR7YXG1gC9drpghds5MbT1HzVORkzyWkTBMXzTJNKujLuHeE9foSdyg/367/8ch5
nFsUiMIcQLVW/OTCcikrjHc5izOj0q3MYKmKftCYZ7Qz8i5LHp9rXl8+1z0Nf51TQ27EgFWA0CL5
a+fDPyudvTmqjrI3QO0r9zbhjAlZvsAgzR49GvXjdRMnyTiPALEDh7NypSo8VdLI87ydoedKIwsE
1MgpocMmo615ctmTGYyblW6kq98XQ4HBx8V+B3Eo64hIm/ekG/NB/WQ/mczFEZpvIDubAjXEVUAZ
FYYJfqgmZH1lXKg8ck/QtRFSO7cRoogKDC3oglo3iegzMt8ZYKTYdIYrnMvpB/4BWZHC2p3cwiRT
swpsvZq0u/5hblCK1AsQPOENidD1QVvwPK0tKRc6vFrJNTbASkFy2WF9AyiVICML3DIPBFmPtlgO
+dAD7Zhxdj4yvda7fron6LYTcWWcaM8Tg2MVH4ffQx9BgI6IPatbTYsEY8tU3A4wHY5vzTniXUs+
6JVirsI/TUYa+YYvTaJk9zqyHzi6+ocA9cBMOiosU0uT3ethvLZgy0o6DFTkESw14gaQkuqGyDcW
oX3+1db5HNhulkZM7tk9fDGJCld/quaI7md0qYRViqnrwvvedoKMOuQ/JFGc9Fc0D2DKtHNtzkBc
yWdH+HAuYemOVxndu0257dLCDj3uQsph11dYwmYONPa5b4j71vwAPSWKOR9fbui3gpT8o3QJtb8X
xPWue+MvXgw/5vPKrraiu2OkoRFT0GuJUkg9Bwi3I54id5ts0iXDYbN97/Taw45Ys+42WC3JtCPQ
75tMoAKVVoXKM4fYu8hiV8PkqAYr4lKU9RZggILaXfsV8bgzVZysHZZ+I6okENz4FqadY5F3zzA8
U540K+9tfz6yZQE2GZxUQzOXUDIxs26QsDH3yOoEDfVqJDR19b174VJTaS+VgH/5OM/ZITRdJLEy
/Ax+LpSAWb8Z07yXU1VzDW5pdhdODrGTRqvt5+xYg5/m5S+8MoiC0MfgKCWytQjLo1mmu5uCv0P0
8M5wMZvRL744+yLHANuBFxOOu+lEeeWjWSllPv4wsLHLzbKf9/kGPZ2SzW4QEE0YOCrmVKkWXxeF
TPLWaAO9c6M7qKcMDG4OZAPh0ktq1xV/lwKhoPDTTtCpfYO7Iv5EZMHtXIInzQf2L0aZvKoNMiA6
Q7Ym5qP7N1oMY8XDwuvTEt5h/kAn4Q7o4VjuA/euVERI2lSBZrnqnpEpwbXDk0FPLMBo+95voGYM
2IYXT74mf2+mZZ6v9eMm8r3HGDKf4j6FOsLIsiQGJGn5lnIFxOp33TgUIfgEhBGju/yaNVjC+4Ew
foNR/jumwtUb7LxrEsTAsFnLbYmnZT7oloqUXGF2jUa0JkAQ9aRTgTJ/VopSgdlasqKFV6L6r0jQ
BcigMoZxtuWpabbLDTMjQ3G6c3eqUQjc+3lryBMBSdmAQVCOZjn7+ruNGs/6FUVRcFEBU7Gqu9ou
uHTcAn20NFJKU7GrqXPbiJjgITrI5RPyeMbLOA0eVL6aaITr+AEeWOfjOkrnYh+6/QwTra+gIZlz
YID3L+/KG4WY+2YbD/wzqFfw574s58k+cw/6tzbjBhOx7YKzjoHesUFX07DNlq0TqEiMbhjEwyA0
epbgZ319/S+O6gS6uKRBVu2UL0oqorVSD8A6KTSOoeOHMxn+WXaZ3xcH2envbawSWDa/iSXn5hzu
6/39FRbV+f2p1DmgzzeCxWepX88aPFWBED3gseGdP/kfdzXzbjmYQHFdXkd0eZxzf2TsZB5HlHSX
F7WnlOQYSUgnsgvY6TTdJFQim29jJwwmun/GhPpkymdr5SrGo5uJrbdxKfETnutB3D3kwmAjOlid
B47uQ4XurfxllQQgeD+i1Bk4WCopZlJsqFCutu8zkDJY4HnEampEx8kNWtbjhGFn3sOzusEvm6lF
OTYB49LFPWtVRFO7IqaKUd2vTf3/0yC2RZ1bkG0cl+StIoTQ/Qs37YfYMq94usREW6Byv3SStw9p
VLvz8657qcdmAqPJC3h6r1zMsTTPLD8WQj/0/8vpMP8skfxX+lTyA673EXXx2u8hbEd7CBEOdHz6
aJLxvgVGVeV/1Nfw/fZ+IniJhDH6V1z60GMzslzBxMJn6ZIaeiWHPVIo5LCa+ZdzfO9zEWH0w4k3
r1jq4CrrZKsqVSw6v8DLGsU2p/6rFmMKWD+bipbhO2M6K3MfsZ8lUS/uJkpp2CMTkXPQ0UDqRCok
j6NiDqxkmwa+jgjLClKp1Jea7V2RhXlpxOsCeqed45rMfCqfTFqZ/PRdMzanuMuPMcLEWt/JuoRj
/QORaMle4z/zz4Ic54lIZVei7cfRHXD00F2MiwaJYYfZHAYabMtGpLLWHhnZBUHsTj9bBGA0NDm/
utk0UPM+2+O3wU35juZDDSIhW5lh9xbCEjEnoFzj9pAtcPc7CHhPk9jVU+q9gecrZH1FVjcXfk+w
MeYhM+S/fxeQP2JHsocd3dKKN0SXg9/QVg35ZghnMBqIqvwXfoIm1K57Z2ykpI4ZlKf0W8tBVOTL
Rz/zuUsIx/FyRr+y5WJcVrmh+dKiYZ2TjxniLsR5bW6h7SxS2iJi3IzLhx0HXN7qVAPpOfBcb7d0
Q7TowjYArdkF9N/v33aV3/SftAigJRyokTgyc8a77JoXjgYXrCfR7m1WtmRECa4rF5FEaOVh+g07
V/y+WB5Ie3ysen+woeu4STD4ftzO/zg4r3tlhcMA1OH8N3Rt/JavIQ+So66+KvYY+ZyRO/lZKK72
uOmSJzndioy/cT8bdDXtYQoupF3spCVT7wuYzZEfI88GPyOEiF+T7YwhJyG4qRo6z3TZEk7GOv5F
eBo5nTHtB/2gH5ycT7QTucV6y0aQbZ/ZM+ATz0h2NTr0qwwRRxY1FQsYJi12H1m90MS0YPdl/4dn
SWVG8DP9dJH2fkSchiCUQ2+ZaQzmQGKjDDCleZ7nqDPhhhABPlQp2rxfGacsGegpnwX6oVLDfzTV
AYtUZ2NgUCQnZGXstBRDqK2NATn4oB8nnI9RvHTQ338OdfXSy5OhU448nAmugEOUyXI0AYkGO3YY
cvEMTJEIkPFqtwN6KTotNSbhlByD9wD7A8EO4tSoImUgLlSaj60skdDokCQsG/QP9FZ5l3eiV3Vh
f2LDSV60dytbE/KjqV0c2Sx8gpWew07Jh7gj3ezo9tMHKTE2AR69gU7q/4FL9I0vlEqnYDUO5Ubc
QokHS1hKGzYYjMkL291JD6COSPpK1TtABUgbVYqRpgAP9xTLcoN9ZU1nAUoN6CyCeOX6uKp+Ae49
KCsuZnRW5ck8N5HUQ72uWAA8Pyf2yvybd86pppEAdOsV8Nwn39sWSpdKQQw4aLoWoUucVZGtz/BU
wcINIH03o0FvsSkZ1BObo4gGmHl6uJsDFUMn/r+EeULddkTdszoIbN/dsxl/TuIGPcfZhQMFpmtL
1F209v5ldh944BGSE6A4tm68G9O6qNh6RkVydAtna5F5vJ1735+7dYEBmaTSGboGwTDG0S1a8sdj
4BUrVV/Sbtq6CBe3JQEatPrsGcswADtv1t5DvuAEYYez3kcCQfUuznPunlylpg53aG30wwKcBuRL
qf5XEZtUW0FRbBjQO/igvRHwImwM7aeaqQ7IocrYSxkVqDZrEGkoNgCETHh2MaHb6LqsOpL+Cdz8
qHA5kB5d6c+DkfWsCWpWsqiJ+tgNTJVAss8FrOzi4H4nvGiGlGn/3e2LOIii3iZPP2tqp6sCfyJD
npqXdcx9UUzojb42zMzK5qytjaQegpkagKYOulnqd5rSHjQoJATpeiKHPFSSQsu3N3bcol2xr+wd
MaNCV59gIL+OmhgXJFPp3L12ryv1iENkQT/Enx/qmR0vlpWG5Be83i2SX6NBhQi15enxthnhP0H1
xSEu8p7K8jf6XLjQOWgEkaU1KZUEc37uvtrHssvmPLC+jj9xmliDwhkS67x+RC+RDpwX7NQLg6oS
NmOEaNcpA7qrR8Imk122/+899G208KLdbnFk8+FkMSWe9PYp6lb/5ofngzgT7B2ZDbTu36LiSf0X
cG/HovWJFFWcIMcgYOXsvcnoaCKQ9waaNcxtJjuNTupqrXDom7jy411GIkPrfEkksYJA27f/HWeq
44b5hh3PiEyYKAwHL8OpXUJovQlNTFkseStTuNGQBgOqD45BQAXC5jRWNen+pVU2D7NezW4zkxWW
yDjPX7avVGO0r8IJHuYYyroPnUuTi8uo/jxxEGpvALG6EptUtnRzeChzpGFgGmdVMrr+QlR9Ul9i
FXritoUcV0+3heEMVGbeXhZnMet+SBSiBlg1GMh7j7l+COVcYkuBfI6fsV+x2jS5m2Lo8lc6jUzR
oTtAKl+r8W/+H/leKJCQkmzVItUOafoRZi8/gXWG9bm/eZTI/ZVxgJAS43gyUA5H6A8P53uNGtvX
pzSgXkaZ6Pn+7+DpGmR08R/J5FAB0vqE9U5JRVokekcRNJ6sdaqIMAdgmmg144vXadbSAlDzgiAD
KVmX21CYcaxVfRBtop9gv9tTKbS7u2eeY2R87Uw0q1hYSgC4xkrea9WaCz9nJA9Q2ydxHgldKvyE
BPqfVidFjvZiU1wjk30dXgi1OzZ46/E5Kso9hI6ga4Mpy6XaCLWNHRwN12X0YZKMaks+LsGj3DD+
k+/Oz1UVRe0pppAeyF7A/0y6ZSZY2CxTnjTNZSWnipidikFLDvP6/0OMKNkbopHqb98MjPgLlhKM
bbR0LIsyVLoNmXZ60DPYwzOeI+bvmQEblbTP/O5kRKtua/zZS+bkXLjBXXikcxSQYXDnjC+Fdjza
n5P3/x8cCqRZKXND2Ur6ynmu003TfPNxWQcKcOFwejat2keZzjgvVSly6M2YaU0dIPHJSI1tqldm
V7v3fEKAeSml3U9+wSC8QDcO/idmFCadNunrAOarnxcoLjmZT7i1DE7H82nLg8BwVrneJbNhyEim
cRABea4q24w6+SB9RONubnO35EKyN0QZf3lcjgLkiLnCrjbjpbmYkPBoh1K2Xgd+404XQ8uCr0dk
g3A2ywcP17rLP/Hn3EZpO61Pr0fzwBxUnhbldDjiK7g5q8kteSL8MmkNjF+G+zmfQ8pG/BQZA59z
1eIi1madyuvMOevKIHktCkTfpkt0Bd4EwB0zu9u8FqO/5GmII0ueU6U+T5ofWFLwK7gBGtu2Uncf
T9Nohyc4/Z0DlAMaMoRb5Byx61dOeMlzrt9xk36hNiY2nnNt8/DP/M4lg2yEnr3Utz5FS796Uc//
5zEsTST1SiIYq/doeAMLhqNEuLs568hTUQocX4l5JOULB78txhIZ2gkC++2E8XuNHVPTmuvD80xh
D9+TJhpkosuXZ1NDUIkmA42fK/R5xvmBbG2qneOaOW646IYHiB0u40gKS8HKJvn/iQqDLcZxryZz
PYunf8SXwODDiOfJwYXuRMOTgxInD5TJSPoGI56wo5+e2zwmPQSKRDa4d1o35CJA9BOOaYrxWT3o
9+9bINY8UsnJwW/n4rnKZnvz46dfnZVQoUdjSv6vCZOJPIJZMEu5BCQKH8ANHf5bURMjoLne3IWz
LZIsLCldFbhIzbHkhp4a+aV6Ln235MX1UEKA8ssvB6uQJ5c95fZBt9mOtypur3pIwt0BAhTtWGRa
K0QWHWz2avpmaEdogV40B6cbB2qTXQkCfLaZo/9CkRrWLNV0cXimYAJY+z4z6iuiOw6heMu7P49Q
7wfAeQO2G0cCSvee3NOiVxZxxkjWyUN8f8+2QcIYY3jdYx5peQO5MjgfOydqlBi0i77oZRntY8Jm
lQU5mESrMARvGNNPJ0Q2X5SYjgZF7tHMsVsGlKX7+LROu4l3GrbTnI63bRYIOEYTMA99ktdSwtb6
qJaMQZNoEIrBkJQhWyMP6qOo9noHLumR/VSBwPbfMeoZC1N42cQRLHRAT7OZ6YOJzPO9U+gQze8E
Hh0RubCg4TMr5VQTxksjubSkY/cuIIW1n2brSDXMp/MKAzTGJr1aUDClluhOYR7DELnWK+V7RUdH
3ArLIFJFlKI7RJl5voel2kxMGn3Yb3dl/Ve4Dr7w104lj75j1li87PQ7+x0WbgRgvjvijjP7drs2
jqwyX4ZXlPTmnsDevHg2GS4Tl85ROLqBAlKcdrSd4rDVZAWEI8edtOXceVY13Ag7KWpbbHqtTX/t
JAFqk7nNwtV8TgJ4aUkN72n6CMYNKf3gux8ckhIQvzpExF7It1JA5r+TdxpT5WVzo9CI90GjamS+
CdRyVtdS/p1buCT5bPjL59WajC5lz/1eiLtogzsF4tpX49GJaurCiw3K2d517ZqsqmU8lSx2jKyY
YAlED+ab76u35z2Qte29mCgXWVabhoKJGOdF0vE+Cv3UXnnCXmgVJNke86z3Z5r+FdGCXRi4/oOz
2wfsFvfXGf/YQUKyG6fUZXRDPXEH/kItAlOT/eK9qikDB7A3wntSRWWQ2sJHbDWacK4WGmIjJLbP
ec0ZQ9xPqQSi7Rt88DNIf6fcweJs+Mlm168/lm6Aoei3grRGx/SCJe53RADOLH015q1n9wPFwNpP
ybWgU0xuoDXwSJ1k2swEpufQAmOPDCm79+tbWHBYBIQWvG3z2dwZK1dD/7L2onFbFxHlwSWKyXT/
TRW9KU9oAzb3h4Q4dpak+xAcDVBU0OwPjI51DJysmzEpSt4Rf6vaSnxnUfSsoavfDnU6cgabwDe4
/7P4IYrDL+HPM2qhhg1qnIvAyXWn5ArMxB1R6HT6JDZ4SzIhFuB+DJLOaD7aVVU6vluQUkbpv0gv
uFnTFaY7BKEKxnVWL6/Ha4ipXPT7FZy0Np7xGp0fkpxbYl56OfiZn7TicXt31qjYIJxsi8DQ1R2K
z/mqkaOyOLfzFIifT2gyyN+kUC+KxWGMLqS5JtxQRwBQxOK6gM040RBg8Dt761fI62Rj7M6CqZ2N
ZHLK/yDXOAyPKe0V6gfumkWg/X9Nda4NkhWdKb+2mZ3fBTQOuGx22V2UUAvfxjU5g4Zcn+bpHjJA
2qzFFuAz7mAeqgjZe/t5lemAIeu2NVSLGJcedOpv+FsORBZL9r/8IhXqezZNt9hu5WMjHKk+MCwT
G0oVdcMeePZfnbNDtGedyyWj5ZgdM893+gX7kP9VQPeAooyGXDBfcG8iJ/68MIzp5u6BrgN0vDVB
mPYtQz7vQowBTih0rm7sKHN0bRO7X8FR8Mb+TJPuBbKjrk6asIASqV2QcljGBD5Vr2dy+y3T6oLW
grZo/SIkMi/6yfb0EK3MU1W4XwvC94/cEaWpZVtytZKjGnWwDkSe8KU5+cpNWW4F2R2cUqZWoCot
nNU1xwzEyebBbUQj2/eCYFWPU2yiWH8dpdkK3UvSsQzyT8SGSlNfX1BXxcKQ0NLDkE5mRrEDidXl
Wx7P5IflUgtVsDAa83IR9VFdSiWQO9ExVDffX+Vvk1Gbegrq7EcY95eQ91nsrAK+EdPknCbiwfHZ
mUMRl/44A6442INGby3BPelSZuTat8ORuPfpj7n3Yf6x9Mi0HrSNQfDivf2rjHRDBbXRrvrnwkrr
cj5Rs5w30/Mt+F8oWgvx2ci8Lcj/oNCvXnrUwDtdOjXnAoU4acPdtYln7hrqjRUIuCGJQOG0Y1Xi
9RGiJQeg1P19j+PSkS0ETkK0NISG/HZ72jUKacDMNByANSRhzOM7VZJ5Y7SR9tYHqoolSPohprtN
6OWycAGQbWBeHUAO8Izmg4D1NOz15Sv0YY+BHBKpqvGXsWqvOgzvVQdACUwfTcYAHD13c8J6/PPT
gHch76yUBxYh0N/8kwL3j3oJ2Eu63sOpd6un1f7cIyTDty2cMkBVQTpeBZcYWdpvu7RzuozhN4KS
zZumekUVTeiAtr+1r5VBJMH29+P5CchEZyC/Qf4a3Faf8RQeYvR/ejdvSOYfAYnqcxo0XP47qP1v
kqS/nTv2SR6xiSVU1tcnsvKQNGkEUc9oJHCqWj4Lr1+4CiWA8q5WdNnNnylul+dWmmx1iAk0mwIA
8JfS5TF0iN/I19nyVse/ztl5BXZlGgyJrEBARnZWcTOjEM/SxhsCvZ+p3dF5gyI1SHKDlOZ0HZyL
J+OMhSdt3NUwgFcd144tXvjgzLII1MHcfTG6i55xzVFzJdK3EnsaDstgEM+VT3yU/NjTURgVLH1c
HWaEG/VbRlbGz/eQvBpW6yrHWSScXef7CnXVHKTS8V1l0fIJdjdTNHpOObtMh6iIbPMbCSgjbVdR
BkJKVyu2qBQxrxItyHXVbQxy3ItFG+rmG4kp1539EPr9OYBopC3/YOLtHyKYxSWMfIsNrFoO86Fd
XoMy3gj7uzAscwTEtA3/I45jB14wbvxMmGqp6SBlxJcPfSAYQ2j2XSl3uc8fcFqy5GWWCsaPBUNY
fZVqDv1ktyFKYXImimEdolnQhlF2Kpz4lC/bOluUJy03t60+oBJYZExP0Dng1evlq/x+ieqJVn2L
5Q6tglmr1i+hkSwzgo1TN1W14dGLg+pfWG6awzVKnYyGogZAl/0i5UFoFfC91ueS3s17k49WHI3r
thqzhMWlZGzRro7OUXNf/OFtPEjB0ujkNToGBhZyIfGcNEbXe5OxGIfpxvI/bptlh7eKomqc2ASN
eroSNoUdcIcxo1/GlPahflA2hiHm6+oXWAujLXC6QSymut2pGUJCMNEvNZNNZmjxOkc0D01vx5Fs
D15WUd1fXthXZimpz7EddG2RUmvHYZ7UotvsX+Z6l4rsINhVn7+Ufufi6zWXrWMIAlWcwQZKuBUB
Zx6YBsS+9hRRibpHJTaj6XRcJxQ3ULeNVxxAnrtc7hSBJ4cYlziJmW6WDbQW5ZMBDKwaYBRgZ/ZY
q1G3LhbQvvKSDFsGnivqzTM27wRK741UhmL6MQv34wYV/4V5CWlb5tBAM41SVgMwdtefKr7bsPVm
6QCwJPn1nAJnc2gkrfO9O/kvhSkn/uSs/HV2Ert8m/sxKc+NgsR5OovySjeGUatDKYTorXt9bMlw
9McdQZVlyzztrvPUg59DGw1379yE9TL7hB5GuYKRZO3lu4jo0a7SgkGsliRNir8g3SvfI078OuIP
jKgdtRjnKOHYfLFWWdzgngOVwa+RDczbaP8pi46LDFrebSBGepCSQRu9c9sgQS7M0vuZCYFjwjzE
92eyQxdbdivg668Qgc8Z0tbEFYx66KIvVtTl6OJslY1X7mTFKsgO1mcIIyEB7N7AxRlStwXZAHIb
3LqQ/rxYmSJXlmara75Aq4Oc9910FU/kKNjphurPZ+AlleQC4O2wfnElAbPcbqVgSkg3mCNjgvrD
JJ6yC9/YCZFMpXOX7GgyBKEpMRC5iDOZxFPLPvPuAjqGLTnJI48/ZOPjH3CepjRj5Yce0To4S+fZ
krcQVRcCugY/tEQwSi9m4xcuMoB03brdhoi2G64VNPdQG3jYsnG2x2QPMRnKonnZS3SfGR6LahAf
fXo9R61GvK2vF6vZaTLcWDU6qyu+0ECNjJcurrURtbL2CEsH/5yG1bDfSE+25bPaxIw4tD/XDRJF
9QX1I2FpDSSdpFYtOG0Ok6MuRJAyT8t5p3LA2kOCFbTW6cxJBKwzinxrzFBOoo4OnOPkcZmFhn25
/wJvvUzUIjSL102uh6owZxbbpVV+b7h8/xisYkpNpqLO5R1zz0mZSuiRZUGLXItku08GUab9pw9x
fW0tIUHxH2Pv6C8T39Fep5ZO5Xn7LnPAw0GnbmpA09s5j70TPA0kv4awsR07yIKZ1LwO8XjeWZbj
Ojrl2yh8dVDM54StdoSEquZr4Gft8N+78ZizaNUfG0bqJ314Xa4ncKK7hfycmlUTFFt+ZD/O9PRN
4/qfBzO9t8lE3EWLQs9gXKJtqVBW2Lc+ppMj+HqyYY/Mb+B2RTXyFHTkRjX1Kp5mB7m66HEpg9E4
MgQ27oU4q9uvzmr2OYCFwDIANNHox7t3Da5b7yg3WTplENZ4Z7igJYgrHNNswnI51BBTL6VIlill
JgXAdqDA8qdD/qBu+bZWlDhkgDfffDg14ILU5k/OFUx5nrfdjyNU7hvTxats2NHU4khLPU4gWZKw
skAOq2K9oDubmkQcY8KZffSR+T71suC/sOHFAvIyO1EadDG89l8ddwMKLy3QwfYrWKvMFAfql25f
5zTdcpjRHzfpVWV+6V1HqfSrCApcZPdfvfbbEJJCcjxnxhZf3h+fIBJOkHDy0CF/vkbDne004Wn9
1u6xmKWNcFCNiPj8tr9ZahR2Ut642qfrYGVK/CWU+xN1cIZ/rn7/z88P3/1Jujbn8yN4Hi25eRDL
lxUq3/4Me+LhlYPFfLbZRvMaiScYWyGuXufOkBbCvndFRnjBUN91uviov+4ChPbxzFRkVGti1vcJ
1o5G3o2BtwufGPYXzTyxF577YN439q+oz0dASeLCiWOe8Yq2Jw261mekXnbY0S2lJygxYQsW7+PC
QMpiYjbWOkP535N3bcJ7y6mvjXPiYWi1AeY7i7kTW1WkK7Lr58U/5umhW3lPBBCOnXy58U0kHXR6
bR7WXfa9JbasR8JqskSnPJaV2XJyUtzPVjD3oLMVQYfz6zYCOtRDg64Z6UVO65X5MbFvVby3kWSt
Yc5ViUkhDUeBEQgE5luB9oOOYyy12rmOUPX2P/fS1UZeE8egGQJraBfHH4gIFJRcAIkZEKuXCAS/
EySQjcTNzRnk08LjCXPx8kQPfOVnI3Cd5E2pAdAM2tWLv6NRTAhuqCXLddzAHe85qffZa+N7gH7x
18kqTwukuyAezszqx4SljLtV5/IUKlSq/1u5k5hazj+GfYhb2dRa9QDfyAwItTXLIfCTB9JM869H
xHMKiDwguM9FO+wTUpNAAegIWsO2VjEE/jEuf1B81vbEW/A1fxomgeMGVjlVvYX1bfE/FcMuKEcf
XVcLrVHm2Q7CNg9n+86ckLt/KVBJH/fpjUJgLtbYy03NCFwl+bKVKKNXWntQC8Uy/t1HauJjo+qJ
BeaFvCfHYUYTTPXhbXqd+9I58Y0MgAXR8WnH97T5dr4VVjkoOMkR+2rcLpS112b7O3LoTF2XZoPL
nC3zqKj++N3psT8fWFYt/5qq/xmCn0M4kEL1BKwprv2B8LxtJm5/6koP2lg5K00RAUYiD2Qb/avc
gG0KBQNtT9Y7U1394sSo27KThLhewY+1czT9ig8ZKEm++9sgALWbklh6vMvPVEhjSS/ChcdBRtxN
K0U/2fs22Wyb4Ue6Ml8B5NsyYFz8BGQEI+UjzZsFrlsYSSVhheI4CarhBkzuU3x9WkjuMepiCQjn
vb1aGDem8w9UbBspPRwyT52noxEs+w/utpihLp6jjlORZkkz3kAnWlOmhSfYHRAOxUQ4fp/7s7wx
DCx96S97o71qsh/MgfCrVdfBpyzIRXWaDO5eUWSFROrwKUZyYbP8iKZcNhZhaIOQcxYg6AW4pUJU
tJvVMeivGXwGa5mkjvM0iGx52g8M3ffLsTkmSrby3MnPnn5SsZiWk0uKj2VK6JqqG0KiTij/bCJA
mf1kDvbABMhuktBq35u+jtcLTP/iWD4CdgJoRiWh3nNKiI4PpxIikhFo8daDo1N5d0Ahg55EBxtm
f4scJFlfYV2QR1SRPIpJWyBjZ43vhPLSUDCmi15D5nBK2BDT39oj6rZ/KyZ1L8cNY1HnD46xauds
IX9FmUvqROwMBAFBuDp+QrtuqC1kUxYmV+stzc/vBQcQ5gtmwZpNu4Wxh2RdbkRQcU+Jf6GYgk4r
kH0QPOiJne/iHkoi5FLGPX/7CwNN8LEnmIgdK5453xrVmTra+SbImcPgT9yiU0WEFMqe42j8pJe/
s+VdMKxINU9orlDT2RSuazFoIi+XvwT7R8KhOnJAB2uQMZbWiodm+3bDy0TzJq9tP6KL3/l/IjxE
b7YPKaOyx0y7FX5uabuBOXqqy1MCLflXtZxDfyTaGlfKNOjf1esSgIijYjG2DxuSOo5HznERj4cr
LqfPn7LtbsqZwe53OEys8QMMna8kRJOXERVt+xKztJXj+TgU2+ivLlX7XQ0pwCS9y6t9r+Y4GSlf
/G05fRRbzWdTJ6NkPXhrReT69yUGmpsH3q3X1KtMhSZ/EBvC8A41lXVcxQbEiqyHZmEOWGZkBOs1
dY1IDiAi5jM7MfbGS0ULBhv/txJ+CC9nMzralmwx5QGxPbPpPRUMVA1lpCj7z/nac7F7cPXC4RPY
iBH6aRqfbtpBlmMMU0GeU2kNoREIXJRXKcdr/O5sO9fOS3T5SsXWcww1f/PaJ3fLPlYVi45cJJhR
SAUaiRGkehdKDblIVIcb8trdPrbAjKQF6dEQ0GDpQn5xU3SUCgO/TW9KJ9uW0dfg/j1imciU2Szj
K/PM28JVYEI/0DTg24y7QTXsjbs7z1KhNqLPkixZ2utFhtRwPMvLVDKWoIro07mQPdlW1S0atXrj
BXdFDZ2Ah+wUwk7QZ53DLQRTUh018TuTnEoboO6OpnRm0SEVZGTNOzxXAcE7XytYoUfyQMBYjwQ4
QTf+b2sczE+/MgKzD9x0YucYahyIydGM4CAcJ4n/50r4U/tCYc398erNqfZmCNjSBWvatXxnLbwd
9rjNEEsZrJq25yEmhEkDeSp46ci1mehDPDxOlQM0bO/N1rqfSBGpFqQ6DobosNRXCEX6nFz4yvZV
dfgTC1YO7zv/wIH6A1vqPODd1ID7OBZRg6YN3g/hbG17tOsP0UDtJqPMRneeiZBk0B3oTlFGV2ku
4pCxe9CCa5qC0TORQcvbPE4+nKSO7HNq8lexQSNN6OUWvxjOXRN8uIYGYzdCwmvScx4FLH+nP/z8
Ef2fGynXf3V7RyHodepD0ifeVUmrrX6JDUdvXP0R1GeD4rwzG/Q21kDtx+yJi/X0IEEqDfF9vUex
/Eg/H80ED00Num7ArWvppuZPMHvjjIEhsn5xZtOJfs6x3W9issRVreVGJfuUlzmaLlt15hdCJpmn
7tJrNT+YVpV1GT9G41OHaNGtaeNy0C1OEZ7YCuNf6pK7AgjKmuJjJpLE1/5+Dh7HMJsiIsok69DE
lLjCDudtkL3YdznFgan9TG/F1l/c3vvD7lAAHK+XgOE35B+cvLbR4/nh7/8wp+C6pSq1Gdk4cBNe
eMLgEBucEWAGwMu3kjB3n7v9ls56yyrKvE+qAqCfaSEk1Svler3NtiQ/LFi0P5FlS/taCpXCZtnA
A3E2PqdXfOx7kAMAcoP+GiRtGHCp9TtCPj57V9jKQObDiAxZMhoTs8y9XYwqb5NgfSXubLiBymHW
mS7OxpQGobYZp8Y96oAENQHCYsaF8WyocOxU1u+4T99pHWeFo99oOLT6BCBMsbkz8JGl11TuupQh
MdYYyx7pPQv3Wqopc8AwEUB1fGhzsYbpq7tZ50JBiQHiYDJxXWYRQ16p0seNSZASqWAAYIxo1wUJ
hXV/+HowH3MbI67JWZAWGq6sDP4iODgEaXoJpQJEORKtGEPk3FxoxC+1DWtKTesWBrHlHMc/ko9a
dzpuPxAYbwcFgOrit75kBL1I6FqmFV1Hv6tWk8BZ9pS4Xbj9+djXEqa+t6aTmSCMAhkYSWme6wT0
Xle2NSiyswTtKe+xU1oL5XOw4czU6MYP0ZWq9nBi396qWjrBzkyEfMvDZcYqoPqzZemjA3m6DETi
d9t0B+cASnJ4DyXT0ZzJmbiwVmXEkZLIpHNsndQ719IPEHFT9W3y/I/ADUnu3JHESqZmpzyTK/Xq
r8gAx36NeOMhJvWydBfCPVwdqLNSExObNZiEqyW8IV1Ro/fmeltLt5LVvp3EB7zJY4jGj2tJudX4
YVbQ4vJGJzwf/kNa6j7ViO/SPKNglQH4n0W5rYCi2Glq8fkQ4hAeuv08/3iBzEbHKH429ifHX6MM
/qua/1XKECzFAUh3xQCT2ThoyMaDW5++XCj6fR1uO6KsryixWIDRqWEBsqgM9Z48nIvxCJytppOa
SjAgkj0c3DxOhIhVWl/UeUmNRVXtr/7e+j5Bcx3Jbbw9OQ0gfr+15eoazW3Act2JrpfQMaC8ljM/
D4WB7cWY7Kk4dB9qE2gusJ1RUgFg7XH61xWy174+wPXZkzmMfqmhij7TjppHcKBBUxKfd8mxUFVZ
LeeGj2m8X4h7umG2VdkHJMQr0bvxxltNveip6WoQARK2KRjp6s86wGd49aZd3Dc+EjqltwfE8tsX
3YEURNlb/2E1yVLN4rt+nQ5i+Y6PiyCsazzxYOjZnxfeN/u2rPvhXzaUMrJI9pWCh5KXmar2TgVx
VHyuLgJ/9Zwjq57F/8F6DRlAa7EEUy/r90zT0cYKt92q9gefMWHQlEdNftFupwYV8caiymsszMSY
SwcPyOnid23QT1Q85tqfWJN0B7fvpjfXyF572Qr/utGW5fwm2fEBnqTdhkUnZ/NrAbdxAQS6ec8R
utVVa1p7v3X7Ki3VnAwFWKSHTWB+1PsY1DV5ZGDLxlV11TlAcEjDuAZ4QZ52+QnCFWC4G3JCgSdU
ACXIiNQkx0LR+cikYQp7ZaTPx5q610d88kR6D6P8ImFHHS75sHPGCljYLHshWl2HPp5pWtQQ4DF7
jogu8BTt4Gtx5Mde/uB6t6q5+gzC1EB3OhMIzMV+yEDnWio8RZmWceERYz20AnuLe1HqxBZd9KtZ
oc8Hjfx9Jcnsd4EfK/Ae7Swnz5FH6pVyUCaTZFuUCknCZRAplsPZGnJNyz6MiK++qmivLVLLvK1+
GudvAIjETwqsrvr6CI3cKujpbRRbgtDKoY8sszkUXuZ4Ci+UMivyhuNC1oqBXut66X5rw6PRFIJU
Tneu0DU2QYWFquAnlApJG8hJM8yMAVrbp55X7CEeQOktHzH0eFVaw3bzvY0oPxmACHYfS6Bed6xB
dA7z9MKDM0V7qzBGEjjZbXI8ZFlJrtRWxk8Xr5hoCyEYWY5WvwUdMxQbN11CRF/z40tGJo6f45wG
CIMiVCMK/Lg9XIgB7nLypTcw3umBn/crs4rP6t2XPGBC0RYPwuhshFGW34vO4Kipphg4ZjY1piWd
MIVfSKpDdBzCBP6BIhQ5OGt1OeAlu96kgqz7UwIMsOVq+a76mv6fGPFzhyp4EBBV+Ohfp+SCNOl5
jpD7uusQkUJQ56K76JCTGU0eF/gyD4aWqTq7Js538pKemrRwBNuY1+jDqF8aAZ6OtgTbXzdJqRZN
EKGRNFlU0atgowUU+q77C+VbszyVXJ6K1pM2hLFzVm9kbbIGCunV0shuKT+/3tjmExg4+xuT4xjb
lJybHlp27dNPxUHOcVWnM2v61pyRtg7nRF7zcJRCX7a4JltUms+QcM8mYwr/4JuEOHpS98dKHN4a
QaFEDSZQfKh9tgHyrr6Eok9EvFmyJHDQVddZOW5Qgb0FNuxPO8VwWYiDYG5NrASPp1y3wcKhEzho
cXLdCT02AU6OfIGyUQcEqOcb0BS9dbV4HqicMPRZkn1mdWLiUxwk/K4CVQgbwdbxchcI4RTZApMV
WAIftdM/lRSdLh9rVzN9rZKKInuhJF1yVFfLg0UihozvpWqXgPJVo3/dyf1cKfEPCE21OjRdUMCj
N1lJID0oRjSH086BGBAR2pU9XUD67K1CQLTNE0frT/cIBcE3iQwsgPoRBXyZMsf+wa6Gh4NhqHFH
0sNrXUHdOmwJjJSoOnMU6+w2L1ZTWwW2SmWvMmT3H9vFl7teJAipfJR2nnyyiJiBrsbGHEYNvvQy
AjStu4RqTuxtLz7LaA4sww7Zp7VakZWq1FP7kmukZPXluO7ioXjd6SqkbUPMF28X4LecR7YJbR9O
vI7bmn7FGpoK4evvO9vZrNhyENj+39BOZJbL+uJtvsXepNbAEe18ln10TQFSNCKjb1BYy+IG1ml2
JW9z3TSgPZvcVCDuwWdvocrpmH9Dc1SiPwtzoDU8QEhpMsX4wkHlf7U75LTmbbWKcX39MLaao29i
NAgXJeVbsZCPQ/csSu9C/hZl9H/8A8Ev5sWS5QNUW3ilV8mTCjaMVumxUH/xhzztE6vPil32sGGh
L/1t4khJZRHfRrLHkhc0oTjb8L3dn0bxfXCgu8eXcF4BERVOSjVbgL1aowqJmZKIgBugdi9lBEm9
4e5loPJbNtPl8VtsjPUZKfyqPDqrfZIVu/vNv9BrRdVYaZ9mHKeEEzdXKx5vV9HHu3TIdZbnKmD9
RkzE8abVh1rxd6gOW72U6jjST92HnukgYFlt49WhRfd7Zlug9g85+6IsXdfVA2FqnMXUFLKI/1cg
1iPQewkC9RGN+ontC5A7tuPn8VJ6ICQknC4eGgCM7pER6Ow/i7YPeGOrxSdhWqiKubeulw3qONhA
gkw0OYpxEz6gzAMiQtWMEgQ7Mm7nNLVwdETgw7boWlgIjeO+Ogn5o7ODTP+l8cK5737GQITmHuq8
Pr9cCQnsbc5Um5SCuU9IR0VbumCTjJmyyNTzLPjstzpT3hQWKzhs3BCIONOiUb8vaDoEcEZt+uDw
080TR/Z2fvEmfM8slYnNkx2XnBUtTxjmoU6L52kVc4Z9d/vHzVVoI9RsdQ8xWTfBOTPfQIk+lGk+
1ewDgaZvT/oWWGcBMotcWhkOCWZKvEuWx4whd5eeP/8tnYQjwh8GMoNt30p6mFklarOzR8ejJCIx
AN4p0fIyHEmM1hGcMrKivrchLSxdOo4VS7SEusZt24/lyy0lWr/d/XHq3JU9ywe1xqVh+6SI1mEz
45OC8n39PERjC7qs8HjZUtXBghEYPOJAHlIlg/FkcszzHLCIxm6fZxT19b9T0PT6RdL5XfX4yUld
e6WC7dxub0UDoqFWyD/HDR2MgmEeDmfm461Ijf54rKwZaUrzfeefartTswM/M//zhZHkbtXrsu/X
TpW9CFd1U4LNyNdi5BQGL4Us7U/+4OZkabWv8AKYdBWqrgyh4Hm2k0MbeFD5aNnw8a+g+eeaqy8m
/0qsBrKepaGl0J+Q0xlv052cHLRC3k7KYsc9tSMqq9TcDNlPSTUTD1rd619IRanizBmA3HFat8c1
3GoLYgrULN/qbJMm1PaDk4d4HzcdUu+sd5oj0ad2ozPzAGwKBBQ0JdBxFJIPZfQWogiZ16rcc0sI
UEouQ6svoApYGAqV8S+uhzQkh040QYSxCpXFGoHaB4Zykt+gKn8NTwx4Jhtnsz2iaY6eWRydJSEa
it8AjEJTEXzHERJRoz/ew540/kcOVWeMvr4Vu/A5Yg5JUUJA9NSWB3bj1LQ8FvPVFFL5K7cQPAU1
tp6SWp8ASVSB4mGPEN84U8roXkvAa9HSZgTbhi1kyzq4Q06lnpV02DvzBYV5q+7UvA5IyDPEPd9I
yZSHVTGndVOeVRkfxMlwt8eE/lTitjV9cxbiGjoecwrkl7qAWcadhHf7C/WrVnJvyY3sCHf/Z3pN
OEkUHwF84aekoStJ9m3vI7/yCl9MFeJu0aDdlRbIrWbp2y/dF+iOq9yn1+tCZ+ZnaSU6BNvLwVGW
/9nylonA9jtDSBj1Kytv/nmaVs7WnGuS2Vcgyi+w/8cHcJUgI4/8VeZlyE1yeQcjIdzZo2dVhkTF
aOohoWchxRsQ9DVuC1Xo7y2hydeGvl0/xN/rioq9036KDCnOhdoV85MmY1bAQ0jafIAH4SvJiPtv
Omsyrnt355t/cLWR/9AloJKacjBHpopp9hFATyVmPggvPnM4I5oeJnejvpeR/EEAFOSzxyYvsINs
bpDHgSONzZ/IJSU7RDY4lE0H7bSYAhAeWudw0nZFRQNreqAgyj2R3wLkzI/k8WtOloBfvlhlYTAG
IYsGg+cX16Bl4cg7mK+eXw4N350ELUxhuO4GrZ/aeG4gcXECoKknK935io6SEdbwvuWOMZsfp0I6
g4NuGywF49Dw5CILF0SWZZAEB1wZKi362A+8KyaEo6maz8icoxdLeO5xYQtKHjgyrjXc/0RHW4Mp
cczQa80iFtPsyP3XzrafUTJzcailkIGKKDUa+GJnPmiEleUkezPresgu6V8CDfUx4vO7nspdaDA2
uzn3wtTBEBjVLyEZtpj70jQon4eZ3q02rTQP195GEkLqdOhuP33ExwZsaKeGYWz6Yp8cyZDF7qOC
q4A5oPIHPHcfOQCyvlphp9zLYsEt8E585du5p6qTm97HIzINszCDVVqECS89FmrAqI39fXXUTMKY
tZu+R9K1xBz0fuKo9UwsVJfe4tzkliqJIuI5KB8TQoj5bNNf0zaT96cgcVRGf8gds3hTfbieEkhx
9RnI1GeyYJzxX6ag+6NClRfUs/7NDUmcL6go/i63d5uaXgq4B9YTGQ59yEgdLu6IPOIxn+V/qVEy
7N/DPCXzC7k5YR7MrjBIMT6nOQsOdo9KLvbcMl961qQYueEi0ejhyhE7FeI+rT4b5gjM7AtPwtn3
OkETLP5IIxNwUdclop1j2ZBm2/aWLZQf30fIHfIc4FPAhOqYHCYxGVYUiNP7RgOQsOjuOfP9Uji7
04Hg+JqonN5W1jQFedbTDBqwGSAlllwN0NnB69wEPtJbuMrEXY88eCGm8u+Iv5VA/Xc+RcbxkI2B
UOfV2K+G9MmbQpq+PFRZF1WqSywGfsd9yi0DGrfcs67KMvgKHV91FSIxICqUQs+zmanDL+66OFd5
jxfrppb5zlRjwYnYJvGYO+pfKFs8WxGXeeLULG7D8cVmC3N/hc5Rvc+YxpB9EMByQRCz+u9dP7eq
0oaOPKvS8cyUODfepaHY1OGVRdqkqxh85onsgd9yBOxiZvyW04fR7bFf4OY/ExHybI6s1cKEX0MO
VFC06VBtfSM0G6flZYkIhkYkJKfCTGqvTIUjog/XUvG2d15Vbby/0PhLxL4LvyzPBF3VFSsbg5rz
vsKMjjdQeWW0Uxxj1+X5sImFugRxJTaEfCYlxdZzeKmN3GFhhwK3+FGZUXnIZCfghPEspSZ7e0um
sFNZrPEDrpMkkx/emirNtjzn4nez9o7wBMQ3yyUbVXAx3juagqUQ9cIxpNbWo/s+gKw6NpKJeLuD
WWSBRhtiDVrCkD1X2IcnPzV/ux/G79YY95Bm+iLRyLRLjGh+QApH7Q/yzsEIAN7by6TfBeKvE4q5
Pds1iWARntBNVnJUgRXxynJ6tpKwN67to/1Z43IH32JykbmDCYNlNrKuZrCf6XxxYwBpiiC542aQ
I+hdSt58fu2bARIsnsHlC79oSLCgiZnHWojDHInK6Ru9IHWEUCqT/YHBRsyhmzXGaSc8HjTcf62L
dTMuCkI6DjKLZVU5XdDEGBv3wu/ghAO2vgfKEF/UrM6kgf3V2w5z3hLCFzrgA0NftbP8V2PN9976
wYLgTiL4SJL9CwW1hr0QzrxHSngMWSnvk56bVIE6ZQYTcG+FtH13MAM98rLu0H8joYtQnlB5Jtzh
i4+10a9+To+QptR0ZsYwnGbvhmVwbEvZsF9PlLbKoMFwL2cAvf5pu41jWg5WR2ch4SlHnynhU1ua
gZK8kHHm3gEb8Au4kCBIXZv7BI+90akBsQiOJ+Y8f+m/TBaOwISI7gvNtq8qgGts9EMupc5oRByO
zy0sqERDvQX/9dgu+dknqg3JTaYDIZ4T9K/E5Mgbs0uNJPc0cyg70DADWiPeHuFlOYGoxKtFBK71
mZHocH7SZtX8pTz9Tk31UcWzSV3T3aJTDiPxs9SLr/353wS84l22G1CBYURBjk/7kg1nR854R8Pa
xQ0D1GKXY9RT46YUM9s4UF2et+aaNVDn34FMU+cZrWGQWtEHyx1Js9membdrKwOvwxzvV03+CUHr
E+/VpFmzq/sesFXKFD5uIP6Ca4ym2UKA96YOHUp07uJrXlIDmL/rMahWxB/ucIX27MGcFsIFPy0o
M6DUTheFR+cJTWOgXqEMgxxVYpi7o2uMuYuAIWmwQiVyw7YVGkjVf0GoDOAsxDP8M95WaJzmLlqm
fiyMZ0dCg9XyDv/JtH9rjSGht4Bzi/OIJ7ZhSSm5+DLtD2OWsTYzFVNTe73zAlVYnryMDCWJgXcs
zeEPgEh7UMlM7uv3MyOR0p5UGLsJu7JK+PLSa7colwT2nvJvQrhnWPTtqjiObmELvwbXr/V5JLLL
TgEdD9MK3nVFvNmcSrES/bNRude/9UX4FPCa2kYhpQZ9BfyXsP23IkTj2jtsOxxQSdsnpv6hFVmi
oDQr1Dk4Jsud/Mw/vwyzOpBJf+lIoEruSD5QAM46l1bIirU5olfWC1C56tAj3d/muajCS6WdoY+/
vNIrf5tamCSMVQylRXUWob8+VZcfdIIncFdpOoQqafcmNmBtGJnB5QrZE3pBKd53fLT4o97a094h
5z62+aa5x97H6BWYMftYqkvWruoPincHK+UShkBl+PD1r+h4m2vewnvY7o9c2v/IAHT0Bp0YxSq6
MzUHP8q0OQT0cvufUq48gpYyHXECCtrODjrEQ2KtxHcuEBp6iT1MaIPRx6xxybgTAK3W/8lG2U7F
r/5elqXpy/hpZ5vRflSq0X+G0xyo8bUYKDK/D8g7kil7x+td+Xf0mv7zoAyes0LZMDE965sdW4FU
sVGWBMJPlnH5KIE8cnDXbeMGHNXxVvlstI1B3GxgPPFBevirfXrr3yYyHwNlmBihgSCj8KweJ0lJ
qmfM3dYXwHd9P09G5sbunn7zyMWPKjC5QRREX1S4VXM8TOvZIzlup+N6s5f1Wtbmm0ja1YTkM/yO
Ixdb1g2lR+rv8Neh/U/HbbGyaiMNMwBSkfSWItJCdM3j4QbvZITKUUUGNBtjJvHvenSGaLphTbVG
sioqSAKYoSbXsxsi/LxWaQZjd+29oiMmJlvpdvxprMiCSTiNbmXCRcnnJNpRYb/SJvqqDYgNkMeW
k8dfrSKhvNUrmz4vZbBhKMCc/q4FsMEtv9ASXVCLIfnH99Maq0GTtxVQjCoyzfg4s7Xz34cgg3BY
coYEpUoeEb8tORPNwyD+j+/L5NBqBBltjkQSfZPmU1CrH361R0wDV2cn4b95LfqGWnL4XnU9nReF
pZWMJdC4Z58GIDDfbouTZ0Xb5HSXqQX0eQTrPrg5VW06Wnfzg+yJkygOVDJbd/wJK26P/3CMLEJA
J4pz652bEnMxkCVJA06n7fmyqKaFVD7HlwIc8zO2vW4dqscxiQAEsZUru1mC/cwSi4HXtU4l/b1q
a/RSIDKV3PYou+p5+DNY3JCINCYb6B7iIPKDfiE5FQAXHpE21EJJdafnXw8C6VchOniwLmVnPUJH
l0FiUbWAsAZSl+L9Sxi3RcJH9CF7Axt+siCDWjzP28B9FQ1kl7g2iJiVapI/8DLKOjfMmu1Q62B3
4vg+Wh4TjwRxSOyIOqFLVsHn51VHlai2Dr5giqhFj4kqb6DrzQf46Jiyi4EFAok9NTBS+Lbf5yF/
Hc36Q/lDnVgTqa1Ar9JTII1vj3Rf09wRpCLIljNmNa65a4nKdpaovTNrnDFCf+Q4EXikrSBQpx2X
YsrKqx7cuxmjJaNSfYvafbz6F9yMqrAx0qPSsEN8+20ucVR0rOcYIHZYneQdM2fMohUdgDEqyIhi
+WFWKP+bTI2v+e8IpXPGEOvzdoOHdPGhQDXMw6b4mc/b1O/aOjocixTN8zb7D+Bvo/ZW2DMei9j9
b4oC8E8C/gUudx0L29GWtjjblMU5ojr1imO47rSDyIpEesb2MYsosr7fuENO+9IUkTKSNT/mK5xU
+byA66AlMgUYYEwsOGCOu16IDxwOYPyyUCqLjF29sKG/xYdvc7aVTJwVXb8d065d9NY6wu7TpPZ7
5kMFT0ALUQKz1boDyR2a6oM60KyzjTfhl/T8tSOJ4N/S6lJ4SmvhX3zbzpEKINL9CtJKucxOvL8M
6kczh35m0rWYc4XljiAv1AsdMRs2/6DYnsu9IBFxvyf79OLG9x7j/uu3ADYcIH5L9TAAU5OnXJem
6v2ktD4TRA3314GxEEOy/n3y7Z9c/tl6pEwWoyR1FfFsVtccBGj+UZultC27hKflC2ZpR8nXFrSQ
0asnrL7A2hrgHAHtgM5szCnw1Tp9PbjsLf85PBGYHsBBBgLEgZtNutxhTANU1UFZ2PWZt/7NKJgp
R09n1Azclkty6kDQU5uZbfSGMYJnOO3ycVqeIAACR2hNVXwo7o2xBfQmYdAgHWjDGUX/uDMjhCzH
aMnVCu7q0vA3M2EiNxUCXKXuBcOUgwcaJNiEhrVzH0AtWukZh0RehM8Q0+d+AsbTquedqtZsk/Zl
DFcXg9y3qYorz88u1Nn0qUbM+qKQ+tKsxWCcIesYplqQ8MgnNjhBok/VpqOb31p9CSoqfSIrY0ts
P+dUG9vrtFfDQw+tGrXx9VGqVO76oc6p3o7ZrUPkxrZU6GAxvYel0mRxGxslw1G6p58Qpo3Hp/1C
MkD28Ou0+tkFnp8GwQwSIUcRuRCmfOjYTBDLef41H+lswvGwDQ3q7wSfNegPlW5sRbd8Bt1Sd7pe
wzUYwHv9+9jBmAPyDSn6OrSzWe6QgKcWP7PqQ6nsCjViBWx9GFWFNtAP7NysvKu/xZ/yaFk7qoDo
DakAEOwX2QP1gAIeSc2Z6RbtFhIk+wd9wn9b9GI6bXE1IRP+JH6Cg/C8CgSTYnaso4XlcDeRW8c9
5rTp6HiocWYns0ECFewg4b2q2mY+pckeu+OOc29L80X0wW3cLqbEuZ4sSdY8hTx/bMZIIFDZPufO
4Mdqi8RTR+ZqGGIW0nJJ2SxRXOe418ttpopCjGpvvrbPoVQWL4cEldT0QWZO6gSibyPLL+pf4r6v
J8eAS7DkeLBR7UOlr59W4EIoyFcLTcXpzWb2jCbqzECRQ4NqsACdhto7ypoKGfFrm8rkRK+IxwEG
3BPORJsjLov0zlO2XcF5rSyROMLBG115c3WEy5Cw55GS2N83h7ZzltjThFv7xymsT/IEkn8J3yce
KgGANfTUFFBxfVcqtH5yVH2LzgaVax9jyEurHOC1sHDCqHqzBwlFpH359NFcRqt8l8TyUeT/rUgy
t0ZZFrLMch6Xr3Hg7YvrhqM0i2pAuLPLQ0vqMqdYgs8XkO+lV35T3Nrsj1gsVcbo+U2zZ8O25Ot1
Bc3NypEjv/51z9DTKr7jV8Aodg4gyPqj64ZzKEi619JWiBur/AbEQmDg1PSbx6T8ZO5/2IxlnNG1
YqTXbxad6hp5zuxNRVq2anqq5tyGnPdHV4bhlU4VfpFSSTkrA5gtI3iowdhxJ5FTVdNWyX5yCX8V
iG++m7II7H+P453n7TbwqX3KM01DGT78ev6z/HIRyN/1Y9Z5FzoaXewqcyIKSYDkmmcIwSCA+N3R
ldEZYAwq1g3DmBdiq+CyYCUbD6W4S1SIUy3xmbwFnhude0v/yhsCAAT4VtzKRGwSt4jU7zTaaLzk
k/jDTMeZgWY17goRT2cNoFhzj+Xz1tcDB0xHy85L0Ib2zNR5sM9xM9hvdJ/lRKDSRL1IjsrmeA9L
/11k00r/a6DATdT4mrZcpKy1TqCeK76RWKPGNCTG2Vk1JB5QkQaFQYNtiJxMELAz1YIo0v2Yx824
4FsciRK2z4NnvmV6tWbBDbzsurlKyZ1crO5UUKArxtCXHuiJi1AtHDDE6fjgyW87p1hbCFryhRNT
7dBRJGSkXH3K9f9hTqM3CNqSlGLgfIbbGtpRR71FHo+oqyzNM0M3kPAfnc3O/zTIkw6/FnrsVgSs
5SkhIFBozC//RsEYnA8kT4di8wu3qdxYjpzRQJ49Bk4X4imwQrWLh1+cZ+PzDauoOqZ043votAKV
rDlQ+FQlY4IPsAe5MBKeezi9K7hFbqfkG4mYWHhCcV4ebER7Jk/9u07j/oOPzM94gT5BE0MmHW48
NGKdqxcnWcu8lFPE8khyyS6ACPN28qRUPR8MNq8l6gGVCj0nddkWD8I8q8nwzBTqaMHcP9mDzQmP
iBk9lu8g8aIwHZg5CgyIQ1eAzs567rQYVXLjNMki5yqC6UA5Uzl+7nTybBEUV6+tiR61wxW+vF7J
zVJ2GlFhzTqKpP7h3IqLVnyjjH0OsPXLCrQ2EhKUGTvtu8G3IhqTdrnFQjt+U8IQ8cpvyAJGHV+b
cF3mNDGwMTrHPbVMV5gCpqHy9wtiVoSA1mwTtJgUXaMxZDNGuB5nSDprfnhPoSN0NIopRH6gKXcV
YQmF+/0cOHkz4Cv7ME5s5D5ezaILriF9uXCTBcGmJhke7rj2Cipc7trsPZB+LfQK+j0xw14Ouk46
JfkQ85oYDlm0It8Mtm4PP92lVj5mDdYXRDjXdriF+T1yAt5u2/N2wU3M+dpzV5PfNEIyx6rPV1K8
QRxjkOKnZ04xE7ImjVULSpfWaHaHXqRLnMBa8V/HosZR2R5xkHIAdVkW27MWVlhcUaqTaeuFv9DZ
V+SELj7wyjrXMOkOxhNLMCJAOSggZYaq+5heRRLyOnYVMK2IclTg1GquDABDLp7trY5DKgJRyRuN
cNi3ZBGFEVEL9R0vQOHaQD/epQOIuwiRRz0B16LmrwG81ILsgQ+evZtLjMMQLYTpqOZgAJTbU6E3
lCkQY0SBoamW17mD3/EI3uxgx8/H0fGc0r5Xz9pT+A6DN1yqqr9dYD7NTJu1SOC+dM5JryR/pnXG
RXp8/3KbsnqJSX6RaKra8SeKfaxe4aCeZP5+jFaBZxVyrkmXnQSClnlO8f3qH4yptx7nvs8K+Rsv
W0GGAzYZ1T9IS8DaaoUAriWXJ61/t7PvN6hGq90kTu1p+qwG0rBpdwixx5eWGOt/DU1RS6vwxfj2
KjmK2/3DaXIdVThUsb9zGr66Fp1CxsNAOROGY3v3wBab/SAd8/mcmkewhcQ/I9x+q8ygu/ot+Rje
Ahf3W11yNdI72fnJQOx92H7OR8vbcFzZbjA4AlhkDmOktB3uyBWqaxa5m8t9a6znr8DyitsbRp0f
p/P5+Qq79kZC1U/qr14uew0Rc7sT+jSQbZSXft4IHMH9C9hm+/9nsU+ekYuJxjMPlefsh737pdmA
GUR9FlzVxeCdfTTwOvpiFMO5v8S072Yebb+FEDzTc4ajiCM8lDvL507JQrYSwYvCMaaTftWmSgg5
OpXUBXW7i1e97yuhtfapB1LnXR/OpZLfdn6+0ugtk3TAnx2aCM4MU6aX7IUwUx/58BoN7417rKlf
FqMZLUN302xKc54RzX2FU/yMLtfbVeFkJt90Fjd4pHzR86hZdS4fHlkZk0RDiv3hGT87FQjclgUY
PV2OsIF5UZCBXG1r8OuVl+IHwZJ1nFSxi4t1By2YIZq4sd+OXhqlAapODeyJWh61hAn8M2r3IUNF
uCFnia4w9cqwqQXJJ5upiSm+MEsSG/F3IZPDtU8ocCFvrp37B6Hk0U0olxbCnsYeHZolI+E7qvB9
l7I1zgp3369Jf20ZlJ91UMrc4K2WhL0PKhluMjhIYUFl8Vr82adHPVhpcHSmTB3w0KFK8IqflDVY
7nAcvjqibH0HIbk904+7tE0d14XC0+oCRloF5GGSmPprZy0OTQkSwQYS1X36ncY029af+OyjIWS3
+vsiIsnpQo3Pgkq1Ltnz5Fysf4jMQL71KYzRFg82ufvvHy67c5mG7WJXh6DUYocHym82Bkjn0BBT
sVhoPrmX0Mi41Mmg6sRlIH5emV64T/D16/5WoOrJNSokWkwaKu2wkEnvQ55SNjVEwOYvNgNISOel
qSITujaqC8pZAdjXv0cdQaDOs2wvaKfThwDqza3Td0LVb+UV2mZDOcRrdGsxQv8fYk0kEYKWH+iu
sxFjFfzUgOHxqXGPl34y5Jq9LbZl3jXBMU1JkmrAXkIkZmYO4aXXwvQTdxXpDVm0SvjpL7qly5kM
lFGZ+XjhWR7wAZt7i158fHkSrLgNrvCHk7PWPqjGZIAr53WPx6/7w42zs86cbN89s3WCBxdL8szG
oGjEIUSSr50Vr1Kv0pbRSPz+kc/mKTkwvsPPBVjO4gvwm7j2qxGnYL2g9voOgZmg338YaHQDtL54
6rdN9/t+5LPxQMQSRUxgLkzQGMLajKQjYTgUhBt/wb/h1l6ydC1ijmRx7ks3yqU/3O2UhAWAoGz1
D8BGDRbnTC0S55GbbDkys3CLOBNz9y0PkuOmBTAw58QGeDd/8HloNUyGbe3MWbt5scsSSP4f/0AG
4PgiwHpbmA5mRz12YMH8hW+BHy3x/d7qHW93Yw+vCwfBqEzuG6xzS/3YgNP5kS2tFHVPcbH4iVp3
2gOiXlAjd836/iv7fp7kO7EidxTGmPmJfEPYiI7ly36LORpdy2OT1I9iiTKrzmAwjrqWIC9r/IYu
Z1RwV3KYEM8GiO1JNLGmjP5mbUJNCXuwmVs+nDCQ99k34mhsFD3Th7JtuDx3FTOrID/g90+9MtE8
LHKhT2DylZ6j8rbClXVG35JrQ62gJ4eNtMjyQTLan8n/uFXRAi2SO30/4r5JoNGsXEL6Q8DSAWS6
JH9+YmsLRKfiDHNhehP51qqJlUvF+AMyfFIvyRLyvI0nsmNKfR4fYYsQ6uZE/8x1tWhyf/DEVxy2
42qVWjx8DU8EflBmCfFc+M+0KemtYEHS5e2MKOaJQ58xiFpC9mybKtM32aqHl6Cll9zuR7MQ74DI
4XnNihnZowKpXoWRQgqAeK6ACB6ig5GCZhI2QcDCcBjB8ztE20HAQmsDBpEytMg9J5Nvs8f6Bf/c
rEJWfdck6f6l6zifDZD2/Bc1kaPuJwhP/oMIWN673I7t0zfJGilh3jFNH3xHVOFSltJVJw+bjAGm
DQIwmsyn5yRD3Pb4NK8ZWeQmv7Un79fr981E+f5wVhP61qJDLhqY+FlCxFUiHsBUxj1Ce4Yi7yDm
aPwXwovc3d+Vs9GtcvARH5EajInyoaKvVc2HDdX6pPFnaZXZPYpaXybpeqeSDQLN7Xzorc6MTLiA
QyTVigCzuxz/O+zl0AMA1u7dD5UAm6bWia//3Tmi22qyLs/vWLl6pInyNMKQ8S+yKKXgvHo9+B7S
+xfqgN0fjFHrb2/pCZ+idyJ9l+CghzLIHazVKINoNXC1B/rfBH2MOgr4HgMD3u7tQq5Ues8W2Wbg
Xn5sEuF3j3Ikfyqa3eu5cJtMxaHyLkkI6fac2CKW49pZ/NfLwnaX56QGWIUmMbfkNCcdf0E1J2SX
QJUDI6lkDLH6+pikaxFCLakeFhfJ5TZTS35scIOx73s5Qv2t+LTwNVNQIwPV2uPjTaUCX8ay+iZ2
CQYWnKgJpKtIOA268ZOg3UYPxVmaqg4udjcVSd++kUNw2DlGHOR7hQE3w0RwMxMrgIhXsv/Vk2cf
y59XGIt/6AIYIDUFdhtuJA2Jw0/zSyzTqzbO1s0OXUBSK7dRQD4AJndffjdoyeNMxrYrhHVyF84X
RMaDKYtCjncRPWb7oGTcg7E7uhH184oXhc81uPGXL2604/INBE5TpiRYXQYRRTKv/d/J1Loap4f+
h+okbLqpH+imCnWHK59SotojnIXdY6lSAaOyNoebSXxRLBKPnr33tNtPRisgd4r9ZujvjJ75fDdP
VQLpSyQZaBv6vsJV6zjcmcSf9a19e4gwk5/UISLN/TpXEMcaV52ga2lyZbimabp/RGu7tx++v6Yt
h+UKvJzW+dGjjZ7uoT9ZUjsgarYbozXyBKij73emKpeyj3XQkuhizOQvcTjMnjqOj6rV5nC6S2Jz
cWIV2r5Y6s1O2iVUM5xaqjc07L98mpemSi0a7Yl1LVOavHD4lv+ccOwzweEFT6uG5aH6sS9UawP7
e3+6d1wOmZQqQiqhY3Pud5r61Y02jrFYJzKEU1kZytzYeZ/wQv66A9fyjeCdgrDg//VhLNxYrAzW
bgaFjIMPgQahFszOjhnqnBkJ9/kx6SEZc4MtlIT+AbvxjQNAHizul2W2orKs6CuzwtCCwySZpg8k
BRsivn8RjCs7xLapUufNAxHe/cW/ee4i5kHad/8Djz1pp3EGe0b037yF4DeEVsoyrXU6Rf0sGqn9
bUg2uWueuxwGitXT4LoWPealAGSW9AIurIRAUCNYigg3SLLoPlWWTsq5sYE6PGssKYB6lbB8lLZH
fkAzUfx+VS4KBGPMCPFQ/qaT6q9k6VqAAYLTV1gAohg9cJhtBKYiyTbJq3SW6tmZLYR3FRuTgo3c
/Tdas/z8n6CNX29FOs1QZePp7+abBMpTZeTOKRChCdZCMVCwKOETTNe2JI7rEO/dglYog03QHJD9
JMb+CPL3omJcD3LLLwdBBxBvudlTyUxINRxsXgxxwtFOe1hX5c4Pu/Iw0LVajkVmaBGDeeR2+jF2
KEKHKLTqSSIRhEYO3h+LShOV3IHgVVyr9yPlMhRcBEJeVnHkomXkfDeOGPjnX1QvZVorSfh6x7wt
kHeDWpaeSIVh245dsHGpcn/HKqT9i/+GyRd9m0C/JOMVuzNb8LSQ0aVJGejHC/fmblyvS4SzbYnw
gAMDkErUIwoo2Sne6Q3iTaXsCi08//ws8kSParVGYDv/pgM9tjEu1sqiVHiGNxlZ/9dcR4OepH8E
xfuPpBwoeGSfFJJZhEYGBL7L3p02IIWFZlckrQNR6icJJRihtTjP68rrs5kUZgVowZRNEkpqGr07
nd6v7RELtcZC1g3JuIqcqfzJXMZW3ouaXmnIFJfS9Hkutn8z+HQdqwAh9EJoetrupgwDZH7lQx4V
+gHa0DoKa5jDGgpls3cwZa5aFrKFW0sNgfrtjU+yLxa3eVFiCjHqmU9UwpzIZSPmJsP5Hq9c7FK5
RiUem74sApoKI8aYB3z8uKbgCz0N6k4EO/CJY7W/d9Pt7m5/JPWEXdANBiB1/JlEYzkv4CvJEsSf
L+J5eKQGqB75Oiqxh4/xxbV7E3qtrXt67DP/6BQsfUGM5QKM8URJmeb1aEtjNBz1I+neUGPCWz+7
naHZudyOeDxK0lEUNL7W+vb4+G90mD6pVyniIMF/wZQKf0ELlOjm2Mw3+6Jw92w1/So5ckrllTC/
kJwTaLn6NAkxWVn1hpCk2aduhPm/+m2xgj5Pqvot/mutc6DECQ4sjaK//xKU3dBw2Z+Z6W9y/fJ2
saML6G9oNRYmcwy2OBh2JiNac8aK0OjcWKY0Y7RDYvzs0bUYHDXCZxao4NzfgXJsFFLUF6LxrOa9
49dxDVEocEHIEg9OdISe3HameiFeDISnDHuqt/FKOJgQxvo+4YZOFCMF4gOERz8BSncwccyb4xPe
+mm7Eyr1HsiUp3Mo0X03RMdce3/D9nHEDIg0dVTNu9z+0rKEmF5eFk+WOzV1VM2rLUYkkeRwlm2j
uyJ/RXiSwUcWiNTnOXiZSFndmGfkitcy7+tjEtRe9y4jKKyANiFAiToVfe/++UCn8zvE8sfT1Ko6
L3PPrfGrUbXjkWqZ6J5lDkcsd4eokmGNpZdkjvcrRTjmDf3hLbx4MGzhsDeu6atCXRnkFgPjDa55
/suSsYbhW1++SrsWez01TChKPY60EvUSWULBfUkf+JzXuw2c19zsI7cfkrbR3aPHS100SwyidGSD
jYi8qspQG0PDUQZlxhpYcTVsBVJhBCv8zUT+TugT7WtS2uUKIjCWNL55fs6RzFeQwQDSxzLgu0Vf
FdZs3dXi346f/9bER1JSLGvMkvkqM7AK72usOGIaEHYq4LsIy1D6+ykGJ0WYzcbF34TSAceoMlIB
PJPgo91Jv1cMnR0UU/HRa+fi3bY47PtM2c1QeeDJltWx2ybesF8YC+mr4r8tsynGXhYXJE1hbAsd
0Y+s5aiDMYPAQ1E9l7wkfTPL4qkb8mLRbROeF1owOkmJnvFcO2vGplRGTTXcb/v771fg2GY23TIN
TFPcpdnaxqqG8QSKR6szCvdBqo8NORFHUbWPDZUJuiDLrXgmeffifvBUF4mAobzPsUHMr3F6WnD7
85vk1UDbNfPS2TRz1m3OXnU4poV5RvxgonALxsBUc2wW8eYWtksZfIq3YGMpgZht5HZ6jzyiGOyk
cQSF+QMJsPJ5FaF+fl+rsHb/oVxYBowi9ywmG4+MS0+ZtunHz6+HKPMhq1b5d05Djcvul4UeuH6X
4cdPlsUeUT8JCR3dZQ62pvO6zgzDbctUGaJLw7H+xtg1YTCtG5L4Y3BIhZ7w0F2/gUDkIOoW+ahi
MPeqs5vuTRUWlQ9u3KE78kTVIga/Vjw2Ab9T2rE87SKA//55hsTGLb5ebHHVWhijLhPoUX6I+CTg
qdn8hjvzzZmqdnASkUjpd3JraTgJMEf31nGUqE4UMWHzsfpVwhH6pKF5Fp5P+GOC3bt9stqLlEcn
73FejJ1yzTYjH5oHrvQVhMf+SVC9p4kr7aWdd16/DJkkMSpcUID5CmPpHQUKaM8CUiB853mjAjbf
zYfhkPu4Tj9G8h+hLYO2s81GcUCalgGM/M+C1Tel1austtc6/DKepvz36MeTQhdkeO/xi+Nhdb7N
3GTjW9v0WYK9vqmXJNt/qEgz+fZFeIksv4HcZh4UmhA6Hd0e67cHkP+GRtCiycJCjMQ+KwqT2p+r
E7fv3EJoXzfOJTfgxIlReLi/ZRhc9jZawqXE4lMNKQOuVF0509vXxyuOFe1r5Va/z14jzs0E2S9o
HR0tXtebTen1HksEXaCfLzJQ4SpCMEfXWex+5l9QQPL8YAXj1r0q4n/Oj/0fUSHsdSSL/qZ9KPgZ
AlC/+CKGsf5gf7JTEjwuaGiXpfI82SN4bVscPrZptm7PMgxNYoN3lNUmvtZ1XjPaiQNo4bGQSnIx
7Dj9I2NcJI7WmLa6KaySo/I3OBHqFG+q1gJDUjxj1p8k6PQ/i+Lxl4gc9ocww/VtaZHpzP25MSr0
C8j/urxueoJnQBPy9MgCdxmANjZeA47KCTF0tlQ8kkgRst/XiWTbcrZziV40tnuN2uRX8AKEIIY6
0zvLs9SgKWFX8Sv7zFLGGz6I9+MO0cP420lvypMzJb2YCjyFd0SCPV0p6wh0emylpMaWFzhXmTcb
3VthT+KbjVqPOj/ELVdl/QaGLKsQ8QJAlEZlba3am7CXgkD+m+8O7nqs8Sfm5FQ15Akcieu1CyMB
JiNgcD6HxpqCc720YDlPvMg2w9fikVWWIava7kEb4dWCDBpdQNA0r8NJHrNi5bfS8ieaSu3BLrKh
QyWH7K+9x4zqtBpOEharxy64NEtciQKJx3ZDDgSXnyYAmeC+5CyqiWhnTNJi9PyTlbZeV3CLor6b
gHjtaMRmAkvSeUthuCpfRS60CmwccKxQ5aiDLvuvSIvUwO67HvqMVZBFGYDhdMwbDx1e73kJtcUU
dwbZytt1OCFKOxHA4MovAQDjNEEXdZYk/gJUVsijUWTQvO9TDv+DjHLNBiBGn+/TnxbZoQLUfo/1
Gp/L8Kda6+OGS3/+I/+y59HfXAXF9Y+1MWULaOQSdoGOLUHFDQ+YSmEyoOjTPhRfij++0uQ/JNQM
Bv30xfwDBcYs8FFhBQlUIFPgE+xohVheQxCRDy0uLJG9wt2paRhzMZoBApy1gqo5KFcks9SmneJp
ELQmcCp2KTrkYuHMjUnzjBQGwhVdm4mQriue9pga5bHTfKKQ2gyvWsMyUOj+PxNV9e8EDfK8mSAI
KKBObuD2c2yEEVRQaCrpiapbc5n03ENAJIiaqUCLEEZPlatuf9kGA3BZ3i+wOte+gWMZ+DT46k+k
OAr133Pxs6WRoGnOqImxINb7sCuYzUA9NbagUdHZyrm95BmHprpmIrECjDHVXgAtbGrZER+ZdsUu
JDYZFq8JxCoKQrY8xx0Qi7UpWD6NE1wkNenaFBRYeDmEE12u42gqbYG7/OdBe6IFje+lDgva6JdX
HQQh7l8OqJ/udfx79VNoxDqgoR1cOnSGE9mfEJkSEHHtsSnkylwfOGsfuPIoWN9VF9zSnI8nhW97
j4y7yoVtpjSad38yXFRZt9NHRw36Dboawi+MMXjkem6BgOAGC7FSPblbwQfyWhuRKcqfbNvzKgcW
UfTl6rJ8KUWM78eq7N+HvTe6FuZ5jGuB4+QnIdURGWjkPudhgqG8yvYPV+p/t81tsYZijtObBIfB
WlhK/P9IsjzJjSmHwggjroGPdapsOvsR45dj5aHg0BbviivN9cALJFZdnsx/kkgrYYW4pSuX0iWn
oVs1NpaK+Gj6dwG7TyYZcV9BgKWntKoTn1wl4EhVLOiF+Coxvdg5+ICwrX1e+lhuLNJwHYYnscRg
Els9/GSy/BWchsy3Chag+PoEPdgyogON8JY4g25+9aoONabT4hsMwJ0PCdaNF8H1s57bVjOdYbOG
VZnNY0KhLcTOYQvORWM7Vqr9aGbiiT/A8IpjE9oEyN3VRPGJIxBkZ1joC2ip2thEHQs03r5szGWr
0YZ0d3FCHaW+ivdHh+sE5Ug+YtkAPXZIF5pB33Yg+CVHWWuD2bx1a+w+I8KZ5WI7jlxIzzPI1caW
cshVx5v4iYn4soW/4Hg1dal1CQjEKacilGjaMm0rOJNsWFa1Sn6X3dHimy00iIA71JHRyUCixvSv
aTLGvJD5YsalSswIMmSD6rkQa1N5OEmk/qTZSQQfqI8sBzSnJ5MOqmqjL5M1lLLpwh5R2oNUk23r
TYY8pz+CRHwCp+BYrXkEVwXWGE0TMbfjEyROyt49unaHYNCSEEU86CAO1iwKKTY7ZokBwv7u90Ha
tZE35QwkGlFJ8JH3dpyWsE/ZLhWkFrUoUPV71hDnw9IZM+ly1A/1nI2RHwP7fVUdT55IHlOH33JT
+oIz4YnTgVSk+aVKiTXO69vGxBN9lzBUYeN+ai7u4fkRyiirAkmn/wPM6Gu2rwVgXxApCpqKCkl0
kj48vBabPHY4OHHE1N37ZrjzrAhL9bH0DSuOW+20kpnmGL4jCASEYlR4s1EluDgyA9ZXS/Bu0GTf
ShbVR7Sncd0JbwQHBFhKE4LjpSW75GE2WSE88IMd5UXI/VgDhm5WJNZZjbjc1ubdyjX3K/raNkLs
RdYFmaF7JP72CPTGE/5/GMQS4E4yxBY9znst7+cZJ4TzDYL182P7YREAdbPQ/bFpQHmUnPJcue+t
9Ud+lXM6HGG3sAnSVdne2gY1PEISpJhrqJS8kN6dG6vdEnFpMr5Hnh7HT7ywUZIA3NuS6/MI3VTn
2PRcqj+OoiXLtcXDaSH/jELejq5l9BjIqERbK5MDqn4T70ufKe0PBshHKIb2FNHjL6tO73Nln5Hf
y0Eqgof4DO1LEbJKBdSsuI5HlqOUe44A0n92C2tO59JR0Em9lFwTP+YWlV0hFF8hNCrIDOuqvZiq
g2fNUKx3YdGathhUeuH4jBZK4x6sh/PGR4vPEshmO/DCIDa9IrGWVUuRUan1T5mdDgPAEgboLypT
LnqVuOjB0HvZVyfPOJ/ityXVAyjpDoX2abjNPKfCB3kGHpuBIn4vzN+Q2S5PaEvgqoHpsrO0qUpB
HqPSSQ34+4TI0Ka7NWerjTwxBkXyZw+zQsOxpf9byYiUUgolUDW8cXQ4BXI/w9hLBGxX3qjL/as5
6aBNzftKmo0t6MOf7KcNFpX+ZDU2S2qQZEgULU7JQwntv8u9TDA/4J8wXgf8ws+CtKWQy35aWGzV
qdTl4LjoHkg9ExZ0Ro6jR3GetXcNEawYQdjexGJwoWy+vWKlmbY2EUYV0GO6DqaIXG3omTEUEYcq
SwMhF93iIfHfrAzc7IbyIQe5mUwRWom/PDdjTGF8cvbLEa5yidhQbkpbphOb0vVbCSEHgIJQevBy
h2sjXSLHTEBqmONx/k5ECGgp8oOarTyp3e5wnXEjmcnQc13toC4SfD3iFczW+/12B/EMeZp0J6+5
W+8R0tqBaMPikl1zs4ZECu5wTl5rRzUrm7G5pnvrAvuAOK7f8LyNZM8dxEhZiCkB2oFC4S0d3IF5
8dk2Hablx57XdLQ9L/S4mbkW/JBSryvtzLSeMk1UX5+s9XG2xwdIMici8xgoKuTMeIez9I2rAXX4
BmajNM/kXVuLr8Y1ptZDAADWRDGNEAu5R8HkK+6Qsl3DnAxJ0u3pNILYTfpolQgbxbuVrGRsAkNU
KciAOnP0LYgnsLOBReJkNGfNQmiDJVwgaIp8lCDJJsYqwlw+fmTDtA+F360KMoQ61ppZDJ7/n1yR
mpiMNyHp+2vFEkre+MmfWmKs6HoeVslt8JxUdiiHRLPu/YAD0Mt4jm2mBRzkRKRYgI4bIW2vW3vS
dhPYVMShcjL96rfk5jT2zGj5WEQPZJsmlCukzUBkgXPZUy1YqOlBNZ2R1LC+uNxvSSgkeTFJAATr
B0aRrB5jusyTPf3kHcG7K1vXGR9O4VLkOz4DxCZTEXLF1dQFA0+FXOD2saHV/U5373VEmeI+pF4Z
r2e5rdRiz6hPCB6Y89ecgsFW/CAs8xF43MfDOIEqmkCaHcIeq4SocyQZS0rytdCUb25J1p9XHGOe
NL5u6imPxP/SVioDyzzsU/nB92WsYL624xTcS0p+Dr97Mk4xg2vOH6j6rOvMPYg2021A172dBrVV
XpoueQweczd2+lh4S82yhhRB1ucU6Udf54B7TNNB3EqepDWfktef12I862WZAbmXKUt5kJP/kzNC
YsV8jQtTlVxX4A8foa3+oUnuAvBsHMIQFmUPIecNhkZeQsMx4IwAhWOL+PjxTs8DnTJkIKO+4nta
g12wDOObYe4Gp2svkOtZj80rs/42Dl4yguz+GiVLTCoA+DQtOFM0TFgikISahyp5yObeCW5qdfNm
QAUv0bGFKT+PhpiyefjAQ6ucp8W1w3fCMcknUx7m6p2ZzTCz6EK5Yt0/RNTExWHMp1FdBaG5z2gw
jIqvVGEAqAbyh7Fo0f5x2W1GPhMThvxZbLS12FFajt3BBbdwHbjM1LZGYU8AyWWq3LosJZAwBf+j
deqdOJ1UTOydx+cYxd+2622OVQgJR00X9CRw2RMpscKgmI8Ia9vRN5giV2VhLWAKauxT59vLgCC/
OCdtV39xM129ucPNj919agCYZhTPxIrJXzSJHpwMF4O+0aNfltnzUfiahuO1TQDs7cuS5OTgd+AP
uSonv3Jw9WybGEqwy+wXEFhwClHc4RVg0N9sJDBH+4gIonHEcJ45tL0aeFfKXFq13i8aZLYKEQVy
9To2ZgOWyd5y4U6LGL+D+CmjenwWBWkHWV3s60l5+BNZMFXwHfjMniiNv5w3eGOQZyat8bSMrvzB
8pEEZyi3vOdRv3J0nm57l/ldEAQh5E7ll+uiUFbnkgnjVgGI5F066OwcRm2Hr0wM+HyNzQJPBsiB
WYKBBwaRAtDU1291CUUnU8qXBVivLu2PLqqTtaJyYSg1/0ujMKVezGk0ItNN0V+Tpl80W6Xe7ye7
2Xzxw3l29YkpUhOdjJYOkG0xmTXmeY/WHpkNaTjVl3pjXPlvhqoZWN67xbuwkJY9Rdd3FXojMLca
eJb1G3hixqQNqGmF7BN7Ix1kUXGD4Dk0NFJjzinyVzeKk3zgX/k5FxupWUqL6U+C+6XQuBxF02/c
byW856rg3495HdCplf/JZTZEks3ZrlCLINFLsWB/Yj3FKm3kYU9O/pOntmelT86zHsaS6xUaa/uo
VldNkixGbTUwdoooVL6NNlIRsFe1+hVROol6F7V/J9G3+Ohddbh4+qq9r5NhMmJFEJkTl064aCn5
bjwNmYi6ITdaGZ9ZHoV4LWQkmtRCXDT6IpY3+XZi+FN/gtS77dZXkGLgn7aSXzDI1wIbsoR0G8B8
zxPn/LKsxVgKynrf0XQFP+gU4aOZI6t+9+yeZ9yrfhJ/fvLucYsI64DguZigELqirSSXSoyODRVg
EoH5ZtSqepQK/1/dM8OWZkEa+42vjfKhWlevMInhZn8Yhhu8wEmImBLQY6xbeEWQwSriVOWgA+eD
p2VQT34SnziM5A7TCovgPg3orGDhS41KPQoqogCrQ/zJjT6IjIKV0NkRF4ACDQtHHXT4oW/uo5H1
eRG1NEbyy3qwQxuzV14boAFoP5U+UHJUP71hY9+82PU+Gj1ORvxJRgHVCmam1RxSo7mY9DOoF3j5
773/ubBMZJ3NPWJlokZYVxf+CijnNjuqk4EbaOyAwcCzbU0ugCLs8u+1gBc0Yr0sVEkEUdSKbbKU
B+ZeUwuONUaPx7MJBRsDK4fHgujiySyBiRNb8YK7vwydkdfcneF1H3EAZ44psJf96TnhIFcwXOgZ
b38W2jb53x7NQHnsTx7Cm4eaccueYy20XDbMfYOEQZm7cVDNo1dp6NaklehEDv3Iu6pcZdIqxwEX
Gv8beEbZXU0fKkyJInefJJuKm/92dYAbvOhb8B4lWjCSUKb+La75bubaeYjfZypX/Kuu1tTsWVmU
43rLrVS81iX6yIHiZvnrTsx6plPj2HpZJQ+YT0fTwIDglRF6QCVNpKr92a+wXWgfx81qtmqT+Ilb
6XHBz/x7gVnGuBj9yKqtaIG8ZIgiGBBuk1mjB+wbua/CdU4WE46LCy+rrhdM8OhLggUhLHGzu640
l5bzg+zq1xc4nYFwxbj/yuUNlBJ/bGWPq7OddqBmtgXeBgfCcMFYRbgNlapQQPKKqpIHpKho72zj
aAjql7OKEyz+5zfZxkikE3TxwRFD2KSSuGoh83/wSkz+q8e6U80U852yM8E3wgSrpu3siPGUnbUs
dvK2UC9Vq7lk8QuFKUmoi2+DUf8pLKYn9RZxBCkeBX3uL8//JJt2pQooDg1N3IzPFmFyA9so+68j
hiiF/YsXCTiOwZ/z4hkV+2yxWJcEKPmjiYLPeOGdPtuUl6T+p0E55nCDGdOYH6NFvGcF8GfyYZg+
kZL5iH/H2eC+AnTTalBbdeCplTUvObCqvNAUYhNOPHK8vzZ85TSqAPkaP/0+f+HaNJGfmOHDnqhd
9E3Nw3M/6jaCufweLxBFEdvKbPSduwHX77QMYmmTzH9Hz20n5SjoPO+F0aHgq75e1b8zARH/88x/
XbqhxyF6Lcz3OcwPVHTITjE3uxtIcrdHo5RtJH68u6BxVxAN30XxwfLIVXgy6ap5fOiW5rPmPupS
cLQxD20hIbRpqrDaR1ImoTc+ayIGr2v0Nw5Oj/96N7g/CtsXQqjsQ7akMrFbBle/C4EbyRgPSzTL
Gyf84tNpUL90lcqwFBpf+nWLZYCMno/JPqHzg2JbD6AVEw8jSMIt4nbzjZbk7W47P3h7Qukm6svx
QJUHLGaT4bz0P/aiXa/4KHLb+cxvz7RIXwwDZsBme7uSWKzC7peBl1gFIsjLxisy+6dTdsbf4A7D
u1oefVADQNOAg9J8BzQr+3449l6b5SCEEf5hrR61NwFCyoEpNGp265qd+m5HDCtlnF9PpiBHr8CG
aZba/T3QZcfVAS1Seqd2inw8RuD51e5cV/8vERoOTStpVLhM8VOTqEwAxLzpLvRQoN6G2BTJmIHB
Fb5LFOF7qbWimdrG6W5knPj8m/QKcMuamehR7vrBEbudZ62QcPZSMLEywcXNJqR76oclfYAhjWa3
bsOLqXTZb/Ua0eDyC3VS3QIfrt9W7JbQBERocltoaRyddRDZ56ps5OFxGYQLSX38QT771M3NsPXI
6IBKlqik8783O8/sWMDdD1qYLffa3eRrP1GOLwkiHv87xFHbWwkQjcjdNgBk0IVfwPAk4FeuGx1t
Vb7ULPV6rRc/mQ7dD2tbEEfhSWNxZlzAbCfnb2jO+shRzRSACoDvSB3pyzkaUOeVPVP3G7/8vAQM
jrtuQ6ZV4Q4O/3e5NrxCTUZJOCLrKqLW/fZZMka0SPWXLAMcGpUdy7or5g83SviMJPgmi0ISY60w
ofS44Ye4Fvw7gUpn7vZ7c8j9zOJFi5uhZN4pukh0/cd/99lmzLJB1wjmF0fXtTOafEcHfKrDqBiK
hol197sMpZSdAZS3w4WLtYM4VgrWosv9AiSJckbaNwyYln4dWRSakHfnyWd6bY0nnBJV/Zbzcnmi
rfhxzZfWr1GlFvGBl/JffpERtoqX4ipmpCObgcdKH3auPPHeRl/6U7YUe6ctUMedWHPkuGcI7avX
IEIbI9USkuFPT4URxbEoL8CF3ZUe6Wf6w34O3Q5xtoiw3Zyrb2hipEkRjIsdJ4wxk7B2UR2Lenf1
wkogntLTLDGTHOUyNZQTkYfNaYElMy7KdhCuZQZInokmC5gQIR3Ux7LJOiwwJmL17TKmbe6MODIe
XXMWed6jJghWrWXMgsYvBVoqSWu0vcuGL82kc0yIHEGuPI3OqIMNRMkybwC3O8BXyVg9FWy20uAO
hsrHfcUoe/RVoiDe+6ixl0FDUReDrIffuzegETbo25ClGSgmqaUbxYr8qUp8lwOP8loLz6/ptmAX
MMhi3aH+82gV+ri5/RLXbSUG3+miOj5zFmV0DuhWVz5Y7Bxf0X15qo+7RxnSKbTOaXZXdimaO/yX
vK1QEvVkMErb1awtD7WFZjmJYcJOslc34stNnliBDU28UJERCIDZCjUzpzjF7nbd786/vL6hPBt+
zKMuKd1V8efkhxh2P4JAgspGDUCumDChcKm6U9Cy9+Em7HwGoQEA2Ms74hh2aNE5gol2sNdo2ONx
1DZAr4M6+5trUFdx727pAD50ooNAtnTnecnvAbbieTXfScLNaNeu208wpe19z8K4X6lGIeZRGYiu
NR/ud3hunxHj7R5VusBCMRtr00YQ26+NCUOu4aGO63re6QF/IHKnEvZVzoTQADLqh4QCsWDz1uRG
RztcXGEc5PKp5JI/Y9Xa/A9YXC6Y+hzAReKrLiKOlQiuEdeZ9ephTXkoluE+ak44IqO6DRfxjr5z
FpD7BDRV/G/go/QWzL/HFcK0SMa4r0bs3IBM0mZM/AVDC1HN4mR1zlzN0G4xg2rnThGo0xy0LKdU
RC8jvvhv4ARO5L+hXPNaMFxMi35ZIiIzZOzQk2SAEsaimMrfvfp34nZiW22oKLbgv086XRD72hNz
82ofrpI0VkYMnqn4pqFUGP9mHzHCYHX0P0ZA9spW2dkO+wrIYB4NH4edOUyhCz2L39nKF6fKnX67
nEEYRI0Tma2WSrXYvH6plnzNxqff1m+RCz0hAYLr6zt5lMIa2d4sXbu7zh+2K+fPv6uO5xX/kA+I
3VDDQJHFuQm83L4oZlEE7G+XXdVf2L84CTtEfMeQatBLOd2r9Dsync2uLfcIDvLOZHk50aI34NA5
xkf2nA23Px8WpYFO/+KOYD/yUM5Fx2uGaZUaXlIUmE/Oq728mbYHBLjikDhHHtx75s7I4bMTsSB3
n79BUsWBARevZ8i3BcDbY97uGYrlQrmOVpc1r9WdLRDCMYUc6uq1mia6zO68HesxNTMMbKrqiy7X
5KTdgGC/GUlci0erlZAal8UxZjnP9oM1GxBAAiCRkzf1nxQvWZ5D3rY97Bn6kCOm2fxgCGr2ytqF
CkxYjhUaH2OgLqn+tim50DM+8zTSwf6A8XMpZnh9UogAYzWK9lDxZkHUrWo48wPgakNw4Wxlue6i
nydX0A1r5no82aVG5Vc5ZOteHvQagCGc+7Lg7Hj2rrBJ/t7t+JYA6bPc05HkomhMfp8hwu3DtD2k
KWFCW2VQ/afAziG0a+JLqTxEY34Y6F+/mRABA1YXt5nP8c9Gu9FlWNOXSYCLnbWTLahhT1nZhPEi
04iZ23NNeXsU9EVMykcqJAAU63nyN7URQFQ2nbMZPl7Gv6VjrWg7NBbJEa4y6ZWucbuWOkJgnYbZ
ride7iDKH1MTffc2Rsm4prF8dc4O/zHBWXV5VO7vLdN2GBDrAxGawNjgkZIlX8sWNb7IZ+W4S/+n
5UgOfB48q9yzr5tg/WV+IDxzcIaQCL9E/+I1i/3xEr3t9l3ufWthfbHgUPtXbVj+myNhDB5DFZR/
l1bGMgJ9YzFDh/UgCS58GWjDI4JyV3Z6MOq4nZBs/V+6n96dEsjc0u7ShkeLKcph1qClwbsA5GbF
EAWa1PSyWoToXEfIb8JkfPQIhYRC0wb4yzv8QXFPzXsui+wi3Q6rmdpZn+EMaVlM1+E+hyAHrUiw
YItXVMJI+DdZ7sHuiKyScLt9amLawlbw89Xeop1Nx5kciTFCU2vuxFFSBNRzrdSV68Zke/yE7NPT
ZzuKVdnU6U8BpStl6V1zCO+R+ICRF/3Ug6hnhr1Kiie+q1P8k7zkQVcVVzu24TWyZ7lpHXcrHJON
Mry4YDsoVbttHAEHkgfrqJsg10USsh6IgphrMJst+eoou1JWnvjnAXlDON+dhgmQVa6HoUZwRBtj
hob2UpL08xos6FuEhVdLgQimeV0v2ptswZPfmvZNVRR5kKpqY7rieKEawpoyR/y52wxZSKUFicBX
jjOvLLJdV6vCWB98rjm36AJ0Z5YGmUbbucbn0wYgjRcLLj0JiSBI+EtkknyEUBXoSXakfPtxqt4i
t32nu1g0fBouO0ivTZEtspb2XNkZ/7ZrrZGQC+zsDcCLV9rhuT8tdeb2gVLlS8v7nzETnApm3uZs
0nYlaLxfkILJvDNBsZm+tTpmjVrO4zxiShR45tNRF9o2WWlBfURLF8uGsy/5Mosq/cWvJ3KWVUC6
FppeFCWthRA9KsyfTytWU2+58J2jEWFujuxvg0Ok3oc/0DYts20dVS8WDXfwV2H0V5jJ4maxbT/2
OUQ06XmLSAI59p69tx2rG7sxsAxlH7c11YHcLgtVJVcBiC3sdlifw8OWpMCBGUKhD+1x62GhuswB
vYwATUZ3eiVS6iTk3RQz3vFimZkyXM2/uj5QkIV6CtMCtM0tP0HDFl9L/6tTtsWAb2V1wLqFP7e6
mRq+m+AV/eA8EnmWuqCzmYduBTNx6eqa/sDr3DlclbzDlSRsi6ad9KxenaVKtZWpSTD1AZZ+acOh
ES0S3Kcz8pzhwE98wTH8VzRLG+hfAhOSB8O+BKj8QcqXucvJVI4WGBHuC/l6rYT6Gb91Ox/lVpuo
6HXGymOETJU16ZLHMmjF1eZ6e30P6HmxN+qQOsGvSxg4W8Uia+8KvhuEEOmWpub5VMEYto1G4fMS
sJA3i1JdFxLv1an8C/T4FLr/HopLo2YH3RTjmAOuhII9wCUBwUFSaNNKvBZuhqNMTNciKcMGIDtr
SakTlPGDS63TSMFssewKK5XqvyxH4dERvRbYAPs7yXl4t5BBoaKJD6jS4h8oOq8c05ELhh16uqKE
PSbhZ57q/sS07BSBK+KaHUDgSFK1TP0AsHHij1vH14wyvRlzpl8/URK4OLoV2tIY1G1uH5hg49Js
NTsmCzujqBf+vEdWzD7RDPe0SiFhZxr1Jo3GZoqVY3jqABqn5iLX9y9+Pd5swhhvC0m8xRDQEaUU
kLZa4BPkHvQw9bPvQQhJq9xpZ4WpibW47d/ceQ8guReByV61h2B383w4S9XaMdd8tC+eu0xIZ+zM
LgOzY0ziiFEcYOpxCbaJp8e52vgrKzy4Vdblet6pBFJvxkICAHvR5vyN0LIQqnLlEtSKqA0TeKgn
8c9rpfMn/C7lkapMoU1wnwq9k+kXPARB66X44zlwTwbWSE23AFKfIslXCJTYUrFqTgNcm11LnLb1
MguxxbGXr6pcrWd88c1YeaP07cOMXtUv5LQnNAcJ9iABZ09ExVEWdD54R0ZHFNwahSR2Xy2tC1wJ
NIN2KHkg+R+L6dYqTiVBNSnpF7Tu+psodya7dSyo2yDPiyLEw9Yh3cczYh67g9rPocGr/sdmp5tD
hX8ze80d8t9csBSs6k1noAvxvevsloNzf6nlmKVUZa7jZj3iIWrCgMvVTEd421mv89fj+NAZCpqU
9I9sCze6ZZr7I2oaoX6leQY/Jt0tckAFzNYKciPLUhbd5nWxP/RJ7GVgsw7vp0IAg0B33lys2i9F
CKzntQ48e/A3fF24/QbAK6QPO0138Ja55OU8z6LOZeY/uqvoPR1XoJNIIIQgLOhBhcuJW4ZnR4EH
pAPMnoMuwtKRxOKZgUVp+fqoW07pEu9oJTG7N14WHXQtEKy8qFqYFj3pyhPqpCPM2HHO1G4dK2qZ
qNJ1RQMDa+nvTqrJZasLWBBnw+TVQ5YRERsPiB6mVkBPxWYreY+ksaeYCrs8y5Fj/pPRK9JvXpwc
2Q7YNVTnHR/1b0ncoOJIo3L1Bwh1evOJOlLES6wcZJAjikC74/W4TadHvT16nN3KKESPbjPsp76U
2XxXojNRi5XsVYcyGs7qSCLVDHq6DI71LdclR+vWZJN9z+Aprwmm/F86k86QIGU/QbKfZkJY7CYx
sesnk/Ny8kAPDrKpBlARsCmPqNDEdWk+l0AHZUjA8xQIU5OjcPQbPR+ZPXl8dl9ZibH2ZbKVrFjI
0hMryT0GuDc8GfNKCLHZMAG5EbfDIJ8QeWx2BxIJ0HUBgHOdVXvEBggpQE2v6BwDF3J4OxrWwXaD
o+nN2QedkfW4PtYKj25xuayEnVguYRmzWo98Go/In7qrqknO/ixaEPxs0hIm2GukhpB6snRw3a8C
ldH1Ui9aXoCuBAO0Tg2PDdJttcUU1MEG8niGv+mm7Lt1LqVzB005iNF/CSvSeLIkYEPtmXViBqoa
RimhSmlF1GcKzsu78uFO8Grg8jSb7nTs+bc9k83eNtqsNZ5/wVlu7DcW72tVs0d7QvWOHiVhYivv
2FRIIrIhxLMrC9o0HoK/lLs1y8066q5nEUcmqQTpT/F3mUkUsf/quSpSjKUIgEZrtUfS310cDk95
AkJSuGtL0IyugI/pDxG1qnSNsoozY1GdzhfThQDShCSS5DhWocR0QIeF705aZCtWoXREPX1wlrBO
S+2RETIIljpHrTwppBelNP6uCqS+TEKIP5PLtv4+14Y9B4rmcexvnbo60IJFdMbFgeyYMm4Sfgp3
T0QFwB9QcQI9iOliF6IKVldRm0LfgoiBsN3B3KPHiNeQg1XWLq6BZhUrRhy9MKkn+QWN7KrfZG9B
q6VtbEPBe6de9wFJfCOITvSULd5qgUIjOsCPUVuNdVwjmEhUQrWWFmQfHEyEkkMpQ/MK0E2xVvYv
7h33gsKimx+fh35oPrkVJrOBCy8TxLzmdvOsW3rn9BCwFN5AWoZWmCEtk/grhlQtuBYukKlETobM
fBeHdprkInNGVJlLC29hsguPvBHBEanNRW5XNhMD6H8Z9jD0KPeeoL93cJDzh64A4CeFFTDPdOip
v0yqEeSiKJYCK6hubh5/xHvlLy5lOvvn6wPDjEF8T06PkgOzNZMCU4mXF3zv0NPoKzJaA+3f2zNc
peSmq6KsWTT33UA0+hsyACmGTmuSh8ZpfE4fIE1XWh1jPwr1og6aFv9fUHsPqxpYc5zVekC6QICp
0E5tiD4JoS1wFxE+aY7092Kc/NskklDeGqTRAXDuBro9UpYV7owU+AYGSvimEmKKbQYWfc6HHUPq
H+hKc30MTdRxsJ2WlCpf7ce0zIkRcT2C6oD99+ftVOgZ/li1tfnJOJAgjCTeysZnoye+11dcahbx
cx8Yq6t2CRu49yxamhLSUt6RkrHzbtlMOaYUlY73tErNs02YXqfgxmBVehdiFMqJFbODO3gew+CK
eCcV8+AP3R9Qi6xvHnZwasD5zzY/kT/Eu+L3iCvVYwy6HS+baqjD4UXf5MdPVdTpV6hJ7CNSDh/8
EZgcCOtgJ+rucvegLzM34lc2s9zsgYU0fkIgY5zNFm9bI/E9L35GB3eiFphnuEUoI55blD0lImK1
7x1GXIShjbTtAuHmVp+k6L/MAlf07LZhQYylEf6K9ReeKs4PKHnSjxPQlhsVW8no/ITLF2UJRTjS
aFwRz3wROjGNPzXQNGbvzL7QAo4Eu49iAg==
`protect end_protected

