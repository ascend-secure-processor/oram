

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RddtphveL9BKrqDZ9RpPPmw6tPEAtSdz1LUFZh0sWXcWeTBOs5xpcLCmqKRTcuCUR9BMDVC3Gkga
BfsdHKX4fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q8qQusBz/cwQF/OzDbFrghMqvCiLpMgEbktU0IrwdhztSvwwsGm/jYfhFGLapkTF1Je0/wo1NHtd
gwrBquk/XlrM3WXoiRIERFGBZKjZnTIw1tdmO6CQvPzmX20GESsUv5nuRgIFqETf/QR5k1wC49aq
3VV9sDIFfHz4tWjx5OI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V62+dYzC2dsb7PuKHbaNG0RZnKNz6mDIWmcutrTstJAnTkBqZkA7RTQwL3iRzsgMuAOosqKsQZ7s
YTMfPT1Qh3sezeI2EJWwq4JUY8kZrdm+6jC6cDSarp0Opv8g6a6QAjL7yrMMOPIflJBSqNxmQdym
v5y4x1FrY49ypfmpSV87H7KTlsHsx0b3Cy4ODGNFyG7Shk0TtOdBGQ/HGIV/LAfA1QROOZKJX7Uv
gReovbJiQ6o45YW/WQomFeg/T+PbqjG8sqpxQrW5ulP/3VzB49x0AqE3cYf9EXfJula7JTf4SgvL
/QzeGSaGkUWTGIfee6Xoma7TZr3v02tDJpXNJQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pdX1U+eiDYC/2EdhCBJmyuv/s/+RXmgNvolp1VRFoe1FDb837aWo+JyY943Xwl4jxT/v2pW0wKPo
v4KjHcVjHFW7zcBAHrm+me9HxbNpUV9fhYMotIruCh4a+8+QcSDIFRn/czfIKSbAMJ9S6KNlp12v
FbZkQhZ8/U00bhtmSnU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jYhwoGYyD5FCbdAe9Lx4kvuqpVX+HhHsqK+FtBrYrBA4qp1ioPdmrBXzjiFIvAgxOoDaB43+ATLp
Aol9sKG7ieBBEuqmQzo2z1UGXVSOJXzDfRtJ52q8ncEh+tYDl/6SnOmx4QpPgvmjrVcoYT7Ygf8j
KhxWdj6V6AetMDWNQk0urfoFQLt1dC3R5bo20COQCfeuYQDDTd3jnNWWwFDKOQIzp5busR96iWqm
6XuwFiBwcoRI2Nsli/lGPFw6SHiVeTGUQi0ciuq0/qiLDiO6GRiqELz4IB0x2R9rdvhyCnCqfcb2
LeOuFFKb14DpzUn8Rdtyn4iHgPXz5n4PCSIGng==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9216)
`protect data_block
NjANS7qZes/Bs2iy8g4GH+84m/4ZcGS6sR+u2ubZs7J7P5KiYFQ1r7IZt0ia5uZ0Ztbd9vBsfEuB
VQ+bMQqiv9frVQMIvtlT78fFwZMjJ5XNAmQ7kyMzI/V6UzZw3tmTFaEDJ9yDQAN/xPb2YrQZ+odh
ByKYcdLoYyrwG7UiSbCbjkNqlFP7gyzp7jjurWlKzogbjBGL0XtNtjb4/Y4rkxAQVXW5N6YAlwbQ
PKUp7wvFKu0uQtsZE7BvXc5l/qNir5Yj7/5V8PJwrKSmSWo6UMmEUrk80eZncyCTKv3YTKS7WlAb
n3nojTrCpNDv9Z2QHDmezsA9Bbe9VA+tb/Biz4CdoV7GRVci6kDGfN5F21rtjyx8jEAC5zoGIfeC
rT5H2xdkkxIgxoOx6F8ZzFMAbB6BbQFjT7IMdNion3aEklzEREQRE0J4GN4iTXFGHvEVGBfZQqTV
NUaBeVjuUNv3ArhNyhbGyH+oTtZOQDZzvB3Yto0FkRPxEc9lZoAI2RbU4KyOecu5QJ+15ij2jW2E
dwl/MMhsVfurKVzh2jw6OwyjS/IsPPALvpkVdqJvsj3q0hQIk+DApItiSUVQn1ojKtKjCgImgkg4
VlyF9/Pl5iLdvENmG3QitZ9xBEgrIH+tWMptuaxMl3+nw2BvPAoLxIcIs14u+mB8pWyHzdU3l4NT
vA7rWM2LA9MSCi6EI1KOFah+m0ndDkPkPtmfCxMtbiKEs/kEpoyKFamfDE5I2wJCrHsRD40xnzgo
8UImfguF9UqfdJ/65o/xyFvHqKUNfA5h8uvZrhzVSMWwo3JHIcMJyg1SoOmMNdHTRQmJHz9mU9km
52UdDU1wlt2nfwqGBXMVJxWExJhj6/hwak6JFNzSRe3Sp6OEKg/gIIoz9ETRqsL7/Ta/W2Mqok3s
8uBZWBtrZ5382gRlRTflR4VPmPyi+VScMMF9DFcqm+Ef7ckKvMZVzuWUiAzGcrRiwJRm2+rvhOfT
NU/tEqOpAZ4AWiR6grk0oaYV/xp1RMn2ZxC+HNxLbXrOmhEnOyqU5Brwh2cvdnxyAAAtaqB/u6jQ
F6qpctVGWtlz8OCNfvfIxxtYvhUQcdhV/7lIFANjsvG/iV1NqxILZaqc/87CtOdZ4Byw6SPU9Pmu
nCzU/v7DUscRnbcnyiQk2Ms6TP97QTrzPjjLOWkbgHkuECw2NOSRkIYxjf/XUO2MjK5LOGVGeeon
aJS+zVrXLL53K+yhqV74CJ1ADZjhHQBmOW6KB8kvQUUwqDyYUXxAR/WTkq+UTojKj5kN3lsp0/E+
MLMCqO/utktjGnjnD/SiGfVMd5UTS1GaVvyLJ8BkfdmOmHDQ44XlK3Nng7K/Ga/oR9k0sxeLuXb7
hmgYX7L/NrQ1Jlg5z5J0+lsvSn6PCkTVvqVLwMOjg568uge9+3cHXUrAWXxxKMxSeXoQ3EBsDMOA
HpQCH7oO43OydPswZE0y8BMIPB1C/tGjUX+V3fqK8CMAumKVU8VitZ9RhoFpqN+tcGTcT88D2/QI
DbtJsNcjeljwli7vDw0hPo5Gqw5hJ/Vy+rvzaDUUZCLJNA9hTR8v10dVjSi4hUKgDTFuCu8WDb18
GfdXA3G9wAZHRtcadi4l/yqz2+7pDW3ygAfOeRwL35wJ9KO0UYH5s1eeAJd6fLR0BWrZAi7W7JJY
Et2cSt6VF43Lxz6OwQm8DrpA0c1+OaPjyCtt45HlHGno9Jge1hQ4OwG/78OSqEoP7ZI6gt6TQNCC
+qbb64aaVVsCiaMJzdgT8Bcu27m9ICjPmIPKmzj49HFGj5tW+70l3ka8k3t2wa176jyBn2Q1dX8r
Wax8u7xsGl0zWpeuu84nNy/MVQYdd/4k70B4+ppeR/gbV9htcLIwV03DtCcgApKZHsksZbUYWsM9
wJJQN58mkRnS8IDOB9l6D30DFPbyj2d90UYaWq6moe5Y5e/3pbU7BsZPwPdF/vFIw5BRR1RWl49G
+O1vRRK9aUlJzZmag7sXKn5piNL0q0Yhm6DIvW1MphU/8NxZIYeiilGdDc5BP1ZqvsvXSCGzqV/l
1ZW2/4YceA/ccUBB5UqzZzoWNnaoHuVTUEDGE+pxQuWO2ffXMNQISQ7s8XQ7o/x5MdLIjUshwKBd
Y875NoELr6/mj0xon7cqeK4JP+XVlJ1tUTBATQDRJt31bZ+zzWVdgD+znH1YiD0GGCUNgVyzieU7
G07dnXphzvpuaiQ2LbKXzqc7+2NaMq99eZFMeFJk/vN6CgwGzlOvN/6h+/N5v9fwnpWhcdni94rc
hLjCqSpJXtIzcX1B5HEe4pNRt5VbTg76aBwkV+19AJqtPRFT8VDcHwhh8YrrbYwE7pp3ZTeBJ6W0
0r1kQDGfHxjyk8yLvAx6YKNFSI3fgZl/ihJjvvZAyQJ8CpU48gwxnlDEVUOWt2pDJlM504wdi85S
GNPn4/Z5kkp3AlTeA8FXeGiA5QATRfTJ7CTnV3F1F2i1b84QJMTtuLZCzxm5EHTR73qEnr51cfTk
QUXgn3GC3gLBETwQJNr8equ2pBarLat/g/zH4ME18awn0Jy0Qzqa8w3F4gU5DBxI+t3n9yH6/B3Y
U2JZYPjqZ+YSP/g+YH+9EBHB91ARr0Ph2jsf32pwBrTes7nVYPaF3NFbxkyisDiwKo8ToqxoDTf9
Z2cY0RvIrC5Ib7/jpQs+ijBON5WI9iwl6nvEScU6cThfy8hL47QRFUc0iDLcztByyYIaH0ASCsvr
AcXcFcHYT4t91ktgIyrvmjEMAqW+bKpurvI3Dh/pufE72V6jLzng/tLEIcWUJYnZFNQNXr7bixvS
vZM3V25TMW2okyPd6NwQLeJDVnplNOFKVGYgBLMYY8kBXrj7+NlDsY7Hf907a13X0Fe6FvU955id
XQUIhH4nTcuiUNUQ/aJHT04zWTtmNQX/bQ6QbVfv3MtWWAVgmnANZIY7JkzECzj0pY1psl02Bnbq
OX4PxupBidxNvuIZBhzqbR5A3q31AYMeM9ldnGUf+SLyoDMvVe4vAB7uopXVqGmSW2z9BMkFYPGg
cX7qrn/W3T8V31M/ccPkZneXHa9GE+snKjWXPxwXJCga+jFXEX66B5a1rTK/b87oAM00Mu6H9RP2
UxvRa/Qb3YdmBKQNs+e9lfeJ1b24YWkOXIjItvqajZ1whvIXpAIsy+2EzfvMBqw2vw/jH+MDD6R4
hb2wZJKQQFfRpg+lk7m+sii0QZeuOk56l96WCJBz/f1H2+Hx+g7Ktvumu7Fh6RUHXTTu3vBLO9fF
oTUyAeZXiVzfNE4V1Ova2OB3J3rmxphDUftswjLV0bBwcD5MtwJspwZ628G0AHG41uYInIGsxwQx
Iqu3p2FNZmcmN8upSauZ26Cij2BqKgXqlltEy1SLQfpe3c0+NMqexNoR36Dak0+a0V27mP+ite36
8Eh8LPaslxQw4AmpeBldAwlcANHXKS4pzXooIPXQmib0yi4Vgnn2eLfx/iUM+rc9WOtfgoA2SnIA
5Tddicig8wZSXp8Jfhrgs5IfTN7j37AguUvb4yA+FntUxKMG9NGtnXSr9lo3a3iPkJg5p5PQL7ji
rUMrTXK60yTyJcRFUa48fhU1Y6fFzIbpoLlygpr7JJFEd9YeRv60c3oqf/RC5Ph44Grl8qaNPQeC
DkDiTNhZbK+6+3Qepnvs4IdWgTrS8G4c2VfuqDhWj8JP8bms78GgSmqd9IxcKpIqPBD46qjC4pty
zEwVMKIEgRE1V5hMjqMgo6P4hmELFcMgdvidDEHJsHk5TOvKJPhYjjHQl1tlo7b7ffUJkUT+xuKJ
/Zwn3eRO/V/Cq7YC+zqdl6XblEc0D0G14r7WbZTm0Uus+RKR1zYYC5t+WS3kRNlucwaAZCwssd+i
Ia8+y/f+gv01QxrpOUNzubf/or0CrFolgxQjuLdw7v6ir6lQwZwOJtaknygSai0kBqg0lBk2Jbu/
oXxY2oScWat5o5yNQ3mOpovT6ObgmjsFJXsUN+75e9Sx9zenQq8r2/OuNRVYsE0tkGV4G9znOvEk
M/+0MB+dRsuOVBryv/ytIdjByGYOp1mRX5+jlkJA6kWm7JIP7YArOrGI7PtRPSN/E5TSnFg3CN5V
AiIYnysNZLYimd+h+DUJ4xB88g67oMRwD/VfsRBlqdmRIrP4VG2d9K52nmZFktrnJ4qP8vkxgMMV
hMmGOpk6BDTE702uo+OVNggZ+O1GArxMYJm2t12fKiemN7qsmwH62zv3ZXaR+HT1jnNXPb+fqUsF
mKZMiM42TINDFosZNgbYxBo+fAtRpIXMOxha9IgYx93uLzuSgATO1/yxMS1UqepmBZX7rrFjqnbm
soahtjZrZj9tr8ALu30ugxov3wYyC8zMksqGxvKevmq/blg8PA4zj69a+SAtNaEH9+wk7DY1jZ5Y
zQhT3mvwxsYjJLy0QMbsvjB8IGckSuMwzJfnCGdpsThW9uf9F5tjdrAB89CpsqhbChG78iyCUpe2
dj1er/HIgYPXw3kUMR7D6/I2ofCIVQg8YQIlTNhGryq5y5aHSnvxjAL/sngXSk6ourhY0kKq78p2
xeBnibctpcdIGhrFkMi2nm21tkQp7l5jvpzbcgtC+f74eby00ZFnIV/TnJcTaI7dO20F3ub70AED
uQWf3JTBuIYmiDGE2I6KeHwidgabSJ3HgPEt5dslflz477SjNy+j2bkmQ17kNEP1lKgk3CvNv5HE
c7cIT2uMUDMBoND7Bn5MriGLNflpRjHE8GnWWmlc2d5rmna/CUWjVa9F8su6WGiyfdRp0EhHex47
8ier/xFFkb4EZtsvyfyq3VC8maujb/RL5FmxXEXEeTt87XcIflVzk6zK8toL2f3sNEiLy9GQ3vH8
VLEkr1ge4Svr57WiWCcXKpU4tukWynw5Unq+xVSufJRA0Wgua4QIfV0vSMfyE+4Ioox3Sb+Y512M
Ri/zuXJ3XZjuwvipiLKecXMISBYBXLNDMTo2IbbvsMRLttKW7y05y1ZWtdMEQdRh3K7u3Fsaf63v
krRPfCfTz5cNtcKO6Tk4N5FcX7gvHWNAhtaHylwwZ0rfujxynowja62V+6lQSipgQwDQbU4Zi32J
BtWRS1PkUSL4w7he2XtsJl6cD9dMJROoQ/eyHrR42HyErSG+fxJYlLBuwRVbMKWPPASUF5fsvruF
xyNuVzaGLclzJP8U1lHd/HVZO7fP/lZq6byFgQ/phqrQUV3tSB0tRq2DCGbfA5y4iWE3SYvKbwvU
RXvNIIDDne1FNIEyJGuUu8v08q6pq2wtv0qpYVvZZrY+PuWoSf6zyK9Wrv1nOQ2b+2blVf3ezFp2
/0oYje4VMvyTQ6300yPtvNFg3qigiy4flqkqXjdYXtG5rfdWN6Fr3jghNSrc7/ADgalx935340iV
/wGVf5y4yI4TlaCm9WRsm3E1xUcgisW6u3pgVNiE71jH9NwDm5RcXWzvX/NqVdnQKZ4C5zfr0GuF
ZlPzKGYB+kkTDKll+Ss3MOIvAGxBlYAt9FB0FaADlV3o/PO9JfPkCiPJYEavwhrSbsyI4YBxOvUr
MfTu7enxpDI5dIf1dPq98COAO+T3g89z6o6ZZJcQ0ORMyyopCQkk9+oTh0ACJ2TAbhWsXq0lWMxa
ZpsNVyvarz+Buq9I0fyac1kpWXyj4S775CE0Fgrd3t2iyqqHaiU1Uw49OgJPw6a9RUDWQlxsMTVv
1p5diDKWXcswnkoZO/50EQwBuB/Xvl/cBu+kDQkfcCNx6I+G5y0gw4+XbJXhgJqBvmHzLp/yfSEu
nNad/lAVekCDApRzX9davfR9vSfMRwSBv9Y/wGtLaz4j0cN46eoMmjncRdfwphi9HIc3T5UMp5bZ
cUglIKplomyzz04YbYqHU0rzs6TAiPy0PA/vvIbrM+W4prhPOxdxQwyc8HDUBGVsdaEsuIaaPs5O
RUrHGcVAGPm7TYP2lJCZHr+hyPI7tJ05WOVMykMiPD0OwFCxyeQehQT9Xya5oGFEudZO1yre1dvJ
O3nQZanPfbXhopIeTr3q+4eGie35a7dkr7DWrSljzxcY8u9paXm1mLEol1dhO/s7K4X2tF/2xLx3
UOEdGOHQsoTL3cANBgVD2ikJmn0fNflmEM8EWVpAWPRMB39Uzl1jeH5vqzlUCSfKSiVVK/aZ0iQz
WfsHbnci9smo09O1iiQTnbqe9vaI4KPU64VXoMv3/Zkr3zqZww6bdiN3v/HjVeLDF/4g4Pzf7ONl
396jrUr4ulCbF5+4M/aVzZP0+qf52Dqm9noCkCfR9DRi+u41WAGtAhjJZdynqH95jwV9IiT6+IFf
VKlYrhdHsp9BDDbnM8Ss3uulRRMGyW/3KZnmEWsjG3rpbdkSr2+QRmDyhVF0o9lfck3MaYW4je6h
ukMiOuSA8V7elodu4q9MGfDoQFRgjxx8/5J+PGIDwMNj7QzMW1N8VwvY+jlwYDYaMDy5KPDD5xWz
d3knYA7MDKXpqGxHRjC2PLHKUatg2gCirFaaX/DF1mRRJ/UvP73pJR5DfEbouLOIy/jvwCGhBF/z
I365BCchl6u0oPoKnOV8P8QfeuXgDhad4gUrOsI9bAp7P/N2R88hk981AkwLUaD4ZYCcx0xJuIIz
vMz16r3rQxpBcqu/Y1OGElPL2FbACOxEnEyVOKiUnkLtJ1DtGBusb1nqyos0VON9KLkcmoOQnEl0
+jppAWUTbl0Jt1UXqj2phHX5m6Yqqx8PpCPw/Fu/atgQTqENDpeSg5lzemwWMao9o7qf6maAH7m0
GVJzFXpXKRQGVGSM9++kQDEd4vr8hI5m9e3zYWyv4LzAz9kXW3mPkHDB4XgO6Q9sSb1gnxViLrNB
N5+Iup1rPhO/BOudsOAF+45jizb26muLpZ5W1Vgyvdamj+Fe6y59bEPaQMFImPD9UeSND/00rSTu
w4CIThlgg3oOKBJKK8kVi2Ob0NGxdmZhw8+ba0khvGMX3TvBAaceHRuce41pjvlYvOLYkwvPchMI
CShuzO3FafjyGXbhTwqp2xMXINuaq1+Vpi/SAIhc3TkqKPlPolkpvEPjyCbVWlpHhSQGHZ1hFfUy
52/Ppo3F+kd0TGlHZ0FRniRffOaFZ34MoZaQ5IarcSXx12mmKsNbzGasLAgj9o7ITo3HeTVewCLK
2NOTdMltrRHhA1WMXog+e8EQvIG4PpsQ5LUEF9PhGs/h97QJCHb6cmtwi8hWkBae7HoD+aFn7pkH
DdeaZRnreLXa4GKnpnazyH74L9DIZqQfPlZoMf9HiKES+EebBnpIs94ZHqBhxK0nfW4JHpOzAK4A
80MHC4AHLUW9PwBzBYrNa+cJ8ObVFqubzsjgSPpbSP7+C5bhHPqkObuYqVG+U5WdPoM6TU88IGHe
64UZLVW7wu+G2b12QvMOkqzJeMRlYtIoDfumvxhSwiNpmFH337UeK5wtghJJaLdPAXjbPP3CxRZ5
rtgK/L0Ok2sH0S6z/wMcbqj7aWRViPNEc1FH9INjDpHLMS+jUg39vlhNKzMSqhvcGMASAXEMs2RE
LVH8r+1ITkEPR8hlpN8KJO0nZ/uNEic0snrYsn2SMEUVGb5FtjrTVGCvNort/rjRwoy2RwpFWySB
QaGWiIHgYZpworyyo+d3gO6hOkNhWOhNjbqUAvKOuVGBiQ8ve1kUZV0Wy8CilJVhSq8h3/EJtbEb
zhcLbiNcgha2xZgp6jAa20POjEwE16GWHPAQGN1Ima5dFXzq8Gs7SDwoPqp1bFRyxSNwzVTTtlGp
k50+3Go2DElKwOcdUaHBIZkW7kGnGnqE/EromIFARbYHitCuc+eqC6L91IJOEuIYhQdM9sgLJwJp
WBq8eJwOBbYvmkpmBYZJn19YGEDK64z5TFbhBQHlC/f8rmrrfes73+g8QjN4/u0v5kAh7O5n3yG/
/vp70GTmhiTtMkP70VYMksbcoVVedmdAD4t6PyPQ1FeZxkY6KbMfl41bbTknW6eb9MzLtavhEa4U
chRXMB2zakBB3IGDYdGcaXDvcVHMUvTkvmHVGWTZj1//fRbPEN77jSHnRNNpgPd3WqP/Lcpy/1kZ
GfMCkBvcTvPKSWDujkUDDxO4l/Lg8LgrW7QouPvRvek3l5P1hJ2KT9GQ3GMofPIHePg4JBYJUfaK
ckiwgyC1xPoo+hse0ZNhOCfyCMW03xJHz8RtG8bU0piggoRGyELnu8/J1EArjOJDE828zln1zZDg
WhcQ0ER6dJX/OSHC9knLUgXiLnygkEBXe1lkeOAALVK0PKpyKkKf4ZFe3mTmE4fSGNqYaeL6mpu4
XKOQ9hGc+AV+7NYRQEMwPQ8G45lf17u7iYsHNnTL2pXJEjs/Kr5Cp1cmBpuvO3/nqMpeW0Nu1n4D
CPfGWUS9cUL1nJje6WDsyzKCNIw5E4sKY9uXQj15vUWUHsDobH4qgYZD5LY0Q2xlYHNgDl/aqlB7
CBeBexekyeH6LKEu7xUlplDN75YCLuc7Kk1lyHOa1dORapEY9FXGwvigEUZanORlh6EAxNovH5Xi
M741NI98mp8HFffvG2bCmsvv0qooDUfaya3yartSJSU06kNQq71LXUOQ7NPkLOHgX4t8k130elw+
dsWO1EeMYROErOSiCKKCxelrH510gS1JjvT5cNyxwS2pibLEzPd86SjTpIPeliV78N2Zq7ZV4rr7
xqhvnV627n9v9h55HL5wpIFw4fLaIx1A1gBJHRuYRMROatrjwlM2uCQhuLDObcSoNrFaKciAeCjU
vIpN1P9CaIaeDMM3Ut00opC4kQqRjOtdz7zD0wFWRfFrtxMLZ7wDGjwRun6Zf4DKcfWnsvdfVQwD
G2Sn6gUqZ/nozh6MnYVakZ8e+faq7s5whBgCa9IYYW0q+MVFnKs7jcSdyXj7EixDEk1PXJgJObqb
bcaLY+MPEsfj2918bGNvBvLIYYyAQoM3B5QONJvb7gXHAIL3oQTFSc48Ig0ZvB+5/GmIUbBEGNTw
QwhZoOYR5C/2hRQdX1nabc1ljcx5KWEqRQ8EVb875+qKDkD8K0k1IG9AM8iz6vzNBMlDKtU/4tcW
8oDMdlw279P0o7hjtsMGr8rroJrE3Vit+CItx70EKJTit0WZsuwfrYEmz4M2wJQAwECCmWZ6L51J
2Q2wO944tMI6dFVstaofy6K/fnLbbBVdL0RWPBrfSuYqCoGeMQ3KDNGJA1iI3Bpp0RX16CEqQ/pt
HlEmQKf5DC5MwNIGmMcGHWyRV3IFynJn2tTg/M8YM9c60AF/Y7NbO5xEBwwQU2lhj073BpcWX5/0
h2Ff9gcKBzvGoNzLQfDaVz0olkyldeFyHJ2gcpeHoCzxtqXba4LerEPuRcdjG3AKUl8BAhTloAs1
F6snfCCDNo8JeB3wPLZxcStMivLhTKwUOn/mfV0J5XLWtpdD9PziSgAoqz1j5DhJJ2sjtAHHeVtu
gjS1JynOoHZr/K3c7Xgw6IMzFAgBh+WWt9h2QYkX/+S05yjT9XxdLRbh/oGCBiV+/ZJRIMcVzlsx
C7tfDKJy1WGzHVejT0Y7SC+5YP1e2hmTTGinGKS9FJ+S0nZfqqx6mM2hBCM0tCAgmCSiJbaBc2FJ
kVBJkdKPrm2/MfQxT4EP0F2UH3CnuieYIZBvOUwz3bj2GsVt3pcos/ZunfrYhvDMIg7r0fsvl8K6
3TSAIV3SUpIDJEulhh85zpTHJo/HLfPoN7MQ8cuoqEFcerAkpwdED0lMYJ3SmmheoU7jc/ElUidm
itJZ5nEKt+M+u4wJQWIdby9hoBXRTEJeJZmMdaxUGETrgpYIItz63llW0rniIwZ3a7SZMGVHZ+cG
LDzOP3oR204YwKEEq8HtUTYQvnT589+iaZxtZkNeMaI9OYBZo1vOQ2O7g/XdZdnhlhPSWqVwjW/Q
K4rVrpkcoS1/Un2PE606Gf0sYUvSHSTJzszjeTmyX2+sZay7s02IUOA7BMt6l0N4errI+v2Hs2u+
tVqRnc7D5e/7X78fE5CcLOc2Jf4KEF8YIkfHRCZd1f4z+Z25fOdW9B66kfNBgO+/P9le5ESMdy41
Osc4eGgbnLqXN5HOzgLm876TvPbKk2rym7tAJF16ltHUXFTX9ro7FsQGCY+geVwa6u7iJq9ymm4t
Bp/GtOKF+jsjCF78GM0SqTKzjNVgSlwsQjH62QUgKmokTa1YY7D7v67O1pH93Ud4jaBS8RM0vYr8
PFV+I87H4cDO+Is/UgbBUyN0cKXV1brMyM1AQudIFNkz3bBiY6sh0C8I4o4xMSd2wtbtvhRxNLcX
+Xucl5/KyvpZQLCIc1u56koiMg8qrfqP9URX83AObeGa7wNJcDkI9Mvs/95hS+cgKnm656ukq1tE
bDGncOIPoMZNgDUX6SFi6gJ7gkhzpM+yPQL7Itvc7BPPMMEnu3HJO+caV3oANh2hQNlb3UsXmYab
+FQaXWrKy7NnfQBdYEPxuD9mYi4zxcWoIGm0r4XGE2zh5h4hNO5rKMGwi9ag3rDORQuFaIeMcLsH
dVoS8vtkxim3cEgahm8D8gCAF2VARW02PnyTdOPZW2+cUopkyx5ZqPbbdK/sJKG5Jk/Cx6DYVmkP
yFab/I4lVRgRuueXPCxb8suDhORrK7aDvQQ84jHBIx3zYVp04/Tf/N79kQ1xw5FvC0MSnzTB4ugX
mZX6RbkF6O90CLHVBZXqAy14e0paHFeBHP6+q1lGdvrMzb7o4pxlfcpA2qQvp/2vW4ockni5HsW0
9sjX7/d8onuenBLL3/Z/1fZbpezNqjI3k+FLx2weV/fIb6U++5IX+fCmqpoCzqQkGK6MZOqZQtOl
n9D8JmE1rNlfi0mG4XOuQ1reUYLXfLRbXmY9bJ6/RT/JCAjHfrUdQ5CA1OCwQJSGI4icaEm104t1
q6IG+CQfIHB/bQLPmbUbbAVuSYoPCvNz/AEwGvP5JTMwOXyaVLgmhnYEVZRIo8iOtFR6UZanpBeR
jZFqiZsTZYDG+q8fZhfIO0PSgCiA/dYMG9d9UKG3hKVd1cvRKGFESzpPzjFNO0zWJdUIXPyNSfZf
yspUgrYqA3eoRe/CMif7bWej+nHNrlLyxNhY5bqnc8WlEpfeR7atGyDkj/vwn11M88JFEt2JdVgi
wLxHvXZeEVgs0Iqy08tTG2iP6Sg42oMFb7/+FuQH7r8BgZStLRu9CZIK6/gw6c98eLdPr0WVkiC1
2uznX8mHuXq3eizBOjtZU4p16TmQU7dwAY1mc4ksPTbmvAn0o51aJ2GYwzLiaXFrXfmFKCqWqLAZ
naj1agg21rCBcMPF+YyEVzC7jArgKIzIRW4DjODAqXyx785zHJCmnV46qUrLJD//iHztjeXm726T
YUvf17ZIZdMK5Vge9vR8APXM36lIb1yO/ohrxP1NxPAH8Xf/1XDvXnMqjUO4sbIiOAavDCeFK9Lp
WbrX0IUBBaZSgLdjETMgGDDC5I415pPRNB+P3/XStLtnJGKLFouaPAkU8UHG4Q/E6EOSaKTpqXKy
/J4N0cnNsZKnmx7J7gMQ+fsEMvz4q3GXHZQ45wf405Vuc0A3euS1QyRT0cUL9s6BK4tWKAiqv46X
FMnQ9kx9cn9AIWsh6tp8d5AdskAbXyzyu3QMntsuBslBzYVYrluq4e+cZ03MdvtmFCR/SM/8daYa
9yN7cyVt/atsc4TCnNXlnyyV1nEIbso8H5AREcFofWuv/6R8vZjT1PZZPqkXT8cfnmbtkUxN/nnL
vxw1taGpuP5Ox4OsrKQczviQ8cumQ1OHVwYXULdhOpP20x6HCTGEOy0F3T1Y5j1Z7VB6wTtX/qGn
fgAO655ZNERav/LFo7MQipb8q1w+JKC3TZzUHvJm1slJAFdAmXsUPVBM1ujySxif4wFFekYAeVcH
wLdsi20hPkdhZzadIMsMKjVSsLxtC/beYf1Vb78vA6KeYvLlz7Cg7oP0AalPAIae7dR3yGIHARDs
p2CEswNdsrrTeJPMlV5OUnjcz9XGbg88Aj1acl4PGkygfUTLiaH3LHBq96G/yqAofClUtOdKKocx
7y+wKvtxfxfZ8MAyVGpNbhwaGsZIHzAzrdXF1JezAf0ChLL/nPmMsmBAghZaWuSApL5RiJbWvWna
CmCxY/FjK7UWf04oT0ckXjNn+Z7eHdqwgn6hLOLZhxAdFK4Kz1Ql+DascMnYEW2AvDJOb1MisemW
gA3vtjkh94BdLzM2JFIrB5bHwnoAmxsW3Cm0iMGn1akI+JLBCliu/fsS2+fMxptPB8kN1pQjybll
wyTP9QHlOqVFMunbjN91/rW3Dv3lV6ccKbzF89N01riK2gwRei+N
`protect end_protected

