
	parameter					IVEntropyWidth =	64,
	           					AESWidth =			128,
                                AESDelay = 			12 // TODO make this a function of the memory clock / AES clock

