

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Dim80MW1FDzDpMmJHDGUKIZM6GOSCOgn8n5PNNThmpr140IugqXlkEH+UWGn4GGamH8NcVHl23/C
K7Z9tEfmYQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n0+ILXG6w9aMv9XBqXuTeZFz8g7Thrg+/RjAvZBWmbMg33oLKLbuZvsPzi1c6p84VaZ4iWNrKG4A
vQPf/SbjQ+TcyLOuqm9h4jUs3NnM2pjLf0BVXBXYzfgiWinyQ5lq8tvG7wi7r7IV1Q0k/c8PHnoP
fBHdkGS2CzSWx5v3oRY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SnPwpHk7sYAL/6EZewZQHl2ygiC9CFTximdg5HEk9gXUzMT4jEgMEIm80K9R0p9tRZpJZIfGkF7m
yz55wwfEMxLlPJy8Yz/wvBY4P08HLFdUuqvXmf9hIjcJKa+LhUPiAgjxlOgN9rK4i+kxwkumF4IH
DvCG9+82TF4WUoh/sBqbaBJlM47bGIDa/gHOhk5YpLTMSYumkoujSsDP7z0DxtbO/qQrn+hggrHE
U8OAUQsvSr8vj9l++TNAP9Apg7aO901amzcZhqIsRUBaL+rvClTR7nPH+7l7oon/995Rukx6j+PP
5Idj002YVDUvnCv/1w+uMklYNp4V6wHjpeCxHw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EQsfHFU7HjRlXIWcOPv1NW7mVBKeZ9qrbOio+xjCwDvbXOd4blv0/5xUDnWJaGbhicjuwr0V62vw
QrPEzz4ozqQqEtRO5z6xsf5UR1Dzv1Z7L/Q3/sRSc6sfwMlgy8yye1xcESwh7O+yvgAORweWkhSm
AdL+wZuwC59tJi7eUS0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R6oVmCiSyuCkOjet92cJkHc7xLJXThwi6DZYFxvm5kxPtPR/UqKA3x99khRXxiTuMwq8Wh173zka
AeG6qHX1IGRz+dBw6LNS3vMEQVCfjs0Rr/3OqQe/J+yAXw04ibSNipF9E7L0ksryrGa0No7SywBT
+jLRh8nsmNEpqfl5+BDOw3nF5G9Nh1bVwm/Z7GlMi1PdUwWvmj4o/mHDsBDXfAEPNolLfjdkvuc7
rKoF75d0NiR1bymse9IBbI8NlCIQRkU5iK1FF3iqRKAiy2Q0ewT1+KkxgiiNFG/PFO04h3eDVsTc
bleZ2T9DNMLgVGy/zhQH5Vcfv2jReOagJFdrTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8720)
`protect data_block
DctkmlrWBb/1axNa6ZKh7K/L4zWf/M9GQRg+kUkJIKLWRDMHuyn3QZOlaZcc7FzV+wYNyb65xSZZ
msleT4M+EoLH0Rjz5j3TSIRjXhwbWIKM1Ny8vb3hHkp8q4Hv6/p1d2oLQXXTRShLaLU5MXOfR48G
TspiGLpsE1IV+BnaHRryeb8Se3DJUQo4uBywR9BapFDe8J/rOY36RHu7mRdWi+eK6y/wh90cYblB
ZQ0Ie/KArSEXbbt+dgOuQnOFO1D3fCkxwsUorGQSZ46U/3IkfAJyvbGUBV7TtFfOSpIjE+2zyrJ1
3Yf6fqaEAD+1oQpkB6tOCpSQoiVVYuwcFarYIvBTDLXRsR8t9uyq/Bz5+LGf5Ml83O/r8o/VToHH
zBkHdbCG+wA71W8RlbatJKFiMeeONVs8XhDOPbIxA1kAbSSo7W3QhcmAbPrDrKQLfuhoU6BQwxwx
l1q482eJ6Ki+RO9xfugn1iTkMquIvvQKEwYxzKG6Mrsg4gRTZX20LZAIjXQMOvPSMqDxdUcHkn4e
rdMAIAZ7cCDUQCGP3sYBGqn186M1S5WWL1fQjiPn903wrwInTyXdjK2Jc/f5Mf5zH948D/dC/4Hv
+KXaKTveOfsps6yeBWB4ah3v2ALMy5ZCsv5tw4OZpGoLL/7vqpWRvHZDtj4SmXWqME9GfriVCvdJ
A80yhET4TvGYt5a70h5VLsiSSwPXnU42fWfx6kDZx0q9e9uUvDdmFUW4YeJFTAY7mmhNuBeqn3yU
0K5qkAl+nq7L82TQRiiu2o2mb9+WZk30SAnmVTSgLxYV0P0I1VXW15WztKMI8TQwc/74NU6KD30g
5tIGQ3hoc49GEgXONptZeWv8o4crlBBV1KKW+w0a+5YqFl8DvkQitmxmw5DOr0TYs6sntxbsWOeV
hLrAOH3RHPWbrPbTpdjJPwVf8D2mtvFVpDQzvomKul1CmLo+ZS0RBFPoEdcE4N6zE9+xN5czmqaD
GuMWsXXOHvohcEvZRRN3X9ZrDCv9o+MhsWNv0Y25sbx0IaB2qG+qE4Dqd8fEUdIwg0lF01byAayr
S4AW5dU6hNNerAH9EdixtRxguD3SA/ZEB9bXGmpOG1pEJaVeg0vsnuBX8pBRw0lS0greRhVe7Qix
hMpeAYHyG/+PPLgWFZHT0v0F597w/HHP1/hsg8Mo8VY0ggeUolma9+/Wmathmd9ZnNYQVBtIY244
l4l/2RWWrxfpyCSxBCuS+ZNyLT4LBeaxWdrUOXrvPyoOlwkpMTG0OWe9BBipm5u9uiF2NiWdYAiC
R89L6FZUh3TGye+xsdnbMtDo4buGJv3YWAlR9SqrqTqrqs6cvVLIGQKzlm9VWy0Ol6qOzQ9ntgQm
wC9YgVxmC4TZiY7lP5Zejbmu+0ZB0yau+ggDtG27irU9GGKzdVNMNZewQS7Go/eiSA5yDIHb5GnA
KRBvgBoqG7H8iI18WY0OIizfRl33fjZtf4pamlNuXclTbgS4dgrVePizWRwtSyHPsOcLhfVpQJkn
crcJz+4jNBnYHG19Trgnu0lIGlh08pNkgLelCjC1tzXQrlEARKryCqtD3GpwtwBeXHLhSxZng2vU
7hUWA13F0hMBua7dyhXVppe2xSeAP+VBD5IqIAziw/BnQNfutpHpDceh6b3pZ/iFJoIUqbvsyLOU
b6uor+pfFQA0xLh81uU3LDWqGx7d2N92Ey3rkCrV67eALn+SF1/1PIShVDww4kvKeqC3FJixmgrC
KLw/5a72obe4dzyttOvz+ehsLtTM/glrS9RRyqUSumBYQoVpxeRRLzKldj15lG13okUDKEKiHQx2
0DJjHQWH5FkdEaA9OtFG4qqLw5+bzBlmnZ/4E8z82k+rcnyq7+KmAY1HNwV4QSWdkUENxKA+vMjK
M45VmPFIHDCok+PMEk1OAkV8NykuNDsWKxp5+tPMcd+Z/6VRLly57ViQzKNucjOPmdM33xKPLJc3
BnN+FoNZYV5eB8hyMDI4Tzs1smJK+D5gpTmjBIBISpuGxETtgNvcbfwSmkXEw4CJk8n9V2tn5b4Y
5LxOYVSMmSRGc4RShNyIjLf1prfffiz+rtUZYER9Wr9jRwZWmXr6hU72ZljmgbqMMySkaze/DTBU
7cOEUaVz3xbXwiU3a1ZR+ApO6Rxds3pL88L5vgE9Vqnd73M4EfR9AYkCKjXNF4S3bQ9UzBNHPdg7
YKqRArEO/jDFJW75N+0mEyQGpHiQ9a0oeDNPGN8fEhlT4NOQz7z7dKx3z7+8meHP2xsMbxZsRtfk
IVZzWCSWmvQe3g0UJZULqGolzZoo6/HheAtpxV0JEfDMqrB+yfvZlIazKMXKSQmObTKSxSlUOcSa
praFyLhGsIIdWW4QXLpv7hHCdoHBMrU61E0QUtiXLJU+/XkA5jGKK5nJ4pKNfFPb78++QW0V7Zjo
syfOOSBFxaI/aZAHce4tB2eM+kyWYGu2yqY4N4nkfag+ePxm/y8EXBlRrsp+UQolLJZJzoaJSVIC
od98VGW2LkJUgx09anZ6uWq7nJ6sQ9mDcSZa3SqxLo8POYYHp1m+t0kb49xwJIc1AU/q79QVjICS
3NW25GfHNnqLzM4uBMldC9v7CpecqqvB2ju0cyUE8zqFmERnfJ24ovsCXBrhTGQ9lPAqVNzlHvHh
cUEdJSJI3p+CdB9/aYi6voO+RlSk3x5SRUCzjfVyFwlrRkj4jH5stscN5Nizi4talC9X2eB6Da19
qzkziAKvjpnq1/NC0r3z8y9XzZ8R2mQs6nMWhFretAn1sV36VSWUGP/7Y7XlgwxkqOHU+DYWFgr5
fXt+5j2BrAY2HJ0gkYS9WS+z+Y2p2uvhs5U1aBxdQMCL+2Q+fnupE8H4ep/zrRhchNnjOtjqYTot
Lh6qZkLw6a7zPdifc8hTSXNEiTcU3t142RNu1tD4C1OEVnqlbf/rwY0pHpMBPrP0b5PMnzDELQBu
tty46RV5ExCikZL1wBY+byKNYvsxzptmbFznW3WM3U7Ljs489Yeh5vIZI9aIGjRQwJttZCIvB/6z
SCwVBJZ6NmiRIj6Z5Qr/Kvs8RMO3Ke4QWVIoy0fVi2DepIVtLpU4r9DUlFejvsNJ49RZMeNDT8HZ
rIK8cO70KakqXopPsQE+2Lgnk3mWEot9KggkLgS+pc2h7vJQRG7mC2Z3qHSowOXCai2fKO0ynu8k
nzere+CMYfqyI3tq5wKpaPZJ25TUr2FUtJLlqYi4H8jW0iaNvdaC5POwXNjgg6paueS5uO/oRvbg
UzM8QXjLlHNZigqwtYpuCPyE4ozH/bsZb+jb7Ad3lJiz33WVdfH1xdspbwi1O+Zs4d4XkL04hIk+
8Yv7W2CI/vJ1eW1s435h5DTE+J1oAbX/fT7v5oFX7nQP44WzEtxy2IxVtZE2JjofWdxuGdR5/VWF
m/q7x+r4/8PO/2Q9wVICE8gJCOisR81GZsmvccgeIdh1dW7MJJiVXbHHqU/ulBvtWTVDTte4hDkK
eaVmP9mGksMhmYdYOSy4EFhLKiCJ3kov+kXSQGB3kXHSzSMVEdlGBkkIVs2ZlpR8P1F9wZ0S2TBw
pXM9MZ4mlN9FqhlYD1I7/UWrpqmZ6sRTWIauP3FycvBcp5Ppu7w+ZbV+i/auQuzODkAXzoxNHzV0
/MEoJIrSMxA6Ub/P2LpmwM2koNdrqjJA+B8fc8HZiJinKOTc/VKExYWoZWMXh/VJ18QdZt+R0u2L
kdzP1qcRgqqrTuuXVbomLRbH0RYRYg5GLULlE2X7N8vn2XWHzUQ0k+wHvU8JLCoQB0DrDJuSr0OY
a/pyBcibZIN3k7p1hgpswKJeTw1znKtos8MIvk1JtpgnhTYUWVJ+vokd/Yl6AFJ26ozWFsGdIVtY
TygR3w9waJl0ZnJsIN8do9KoMXz8EN0sVcJYrq4IGEc0zbfG5IVAYdh6l6OuUuQMiDOb4ktiujgE
xqOhobg+SMvoOOiC9CoVrs2Pupint0SQgKxok4lFmGca/uetfvClRrjCPieNrp913llHR7kpLtMI
YW/aClJH78fjwl7fBFacs7T90T+vbbc7E2u+bznxVk5qrtV7nChbEcj6ff2GFY+63G/cFNx2CBTJ
B0Mk42L9FKJtRMNeduXdzwCaPiNNFv+fd1fS6zh5pVGlfQXN44MMZbj9o9vUGfc3zp1kCdbXPQTl
U9uhNDx6JJzPzsOafWppV67DEJ10V41VPtoqfM26FSDnNvPSjP5GZDIilW0Y6HGSmKTwXDnx2BMr
ChBIddyxLGhCF7M7D6TkrS7dtjwCzI+z+nTROa09rICv80YetAvXNmA73eo4Go6ZcI4cGPdgiwC9
eSPq9wR8nlKqTP2pAyw1uvOknYE7YYkM3Qpi7vKH0b9HXovhBrNn10eb6ipFZHKf2Q+6BqfUpz9/
VmPC2FJma+ZbHAvvGf24l6b9H/0PJJIPhNXnXBcQbqZJzbUgQiaFCyEX/Lxv25+4/oIgNrNaCq7U
qdMy9kOF2p3OFCWeXPmoCI6xeXojbhr2hIyqzLYKSd9aTfl7QG/c7/X6GVET2OZ4eToSix+JZGhO
cB3VSOg3sXjhEgi8keto6F5rs8hTEGcSSNn1vSl7rSySlZVPWSPdf8GlVEF5nlzVXIGDTeWoxpiv
hwjaMPQrTSZ/kGvmB1eYYDVgd2MTfyq/5BGFGo0eniLWeGtHCjgycSR22Jq2LTv9pFEcLqxPSS2v
uvrotOJy5B0nLPxv2+w6mwiuwodQwkh9exaH0p5y86H0gruaB8Ok48KaE+EvY6dC+TXHKYoSu6BB
e3k60/5+7izHl21QtHJ3zIetGOJJsgtmnrsbveo+Y0/NSzP2h/XeVAkQC9QMGKV5u144o2yZyoKp
ul3CRGMYnu3CMwwrk3ny1VrkbibgNugxy6plBmwj9YB/i/wujGR9DfV9MIisDcQbrH0wgz2TQeN/
vEJulnubnq4jYePR04k8XV+IV/NrV+/xcZo2DysWT5I9lvauwa3MUk0VPsRKrhJVxZK/DJCDoES1
JHADNWCt8er7XKM2cqr8Ostg3UtBytEfOkfPN0FcjLN2gjMgR1hskFIzwCEt9+A4r8CTwM5joQN+
BbAC2Pds+sBb/DVL024n6KFd9giS7SyEWKchcpzhFEFFJOxii68Z3fLDZeIxJpqTB7kpLHn6HnBI
+B2DRSlzvZ5AROqrUDjstalKBfZz/gsPtB9V297s2GT62brsYaofoWvyjik6p1xCODzlwPWt9Pt1
H9x+qjiu0BOh82kvjM+Sd0nMZYlb8as2SYm1QiT5tUYq18v69ZnDAMydCbcwNHgKMs+/t4HdAmyq
FDPwozPtJjJqhBE+WvEQQIBRuyhjZ91QwHgnrJzxRS72ei0TGTkrCpAQPVM45hU7iHWFJsLBxp/w
TWN4WpbjBjW0rthBdlGKH8viSwDLYoJbLJaHCSIqP54hjYWSzXXWk/7qS74dJYbTqC8IxVDLER+P
YB+9aYXmQ/r9kas4rJtdYK5fH7/Wk3byWhSOE/GZqJIuphETIQGvbvi6QCoMKveTDjQC6isS5vNM
Eu5QtD8EF1uswH2eP1g3FoLi/wf++NvvGL4q5U5BHzjvEyw7GTa6rpU9VEJEmZa5LUd8fKv0kNvg
X6tKJc52auwckKCSxdh0TzsIhDUeTBioldpv21AZ7ZYpOB/+Nhw/VWfuKxqoSdCbTjkc/RFo9Oq4
qypgrKiHOnv5kJgeJK7GVBPV7BBla/AVa1Ov9SE4a1FQSVuuuyqM6woPN/UzkpOEekIqkGDnej3H
tighs27GPBEkQu/4skjRwtW+SvD6ZsjKSxeM+CZG0KbxglhsisdxWn8BkYU9in5RhXcwJRcEpI/u
vPo28TYm0aqAzAYw6zJRqjzFTLWuzgQUCCHEmYvSipUP/CYtVHJ414RIFTsvYHEkZtsvCSOeRP50
npD+MFpTTurOXcp5Ez3DKsjJXAyREodjcEXnOUj3J9gVg5x7DkL0XmoA+zpBBGkAOGp+tzAF4aWw
J0PavaOczgz2m8fCoGu2ZutrT65d/PeEld32Vp5PRfmrj00mhSgpHDkaQON1C+ePN9Tcr2VcmTnb
hProdDW1zMzo3akZ0FtC7fcX2tQkYEYYkLl2Y0f4or9citthddWjisfEDJ2/QpDmZwSc/IyzKx7O
ZCCqy/5EVvjyIXzk6Q/kb2jtG/8MfR4QSg34gJFNyRb8AmbiB2iSzlHQs5BZ9y4FqMpQsO6cGFIL
CKJpboxEX/NZIGKL1WqgAxTv8RgMqvYF6LXYW4DdNfD0b7xNHZd3ESAbGKJpwowziZYgCWQ2j4Ap
GV2DQtYr0WAIKWjAFVfHwt6r5uI3GR1kuJVPvQ6yDDSUv1PnO2YjjlPuASJEkIMxKtQ5Kum7gTrD
PX8rdIRy2n3/l+lQVv/xier/W85R2d+Qzihgaz1YRmW2Ygd/ayNbokA8BREfcTimEzeMVbpKJ/dF
v/CZAmjSi5O6rmh5DHFctW6w5rZPecM8dXOIW/Fd0cGDCG7h/IOv05yMW+zUfgAeEBkrQrIsf5Ng
aAik/OzjkASV/OXfK78O+wbWB7R7VJ/yPYYucHJpNjvkfJAVrIkMXgdXdcuOjMolwWcsUPlNFsAC
JDAa/9nrbIKaQ/vrFIenLKjUqYAkIPV+PuM08mUL4eRwzdNWqZWruASF2tNMrGVcryyuH6Omxcmh
ymr6zyCucMPDOyJqutWZ3NQ/o/KgGi+vR06igByiQAMCbO4ccLK+Z2vs6irSxFvv/KL6l5sqV+K5
Q/jQHecI85i8/coMoyGktupuJ/QdbUNClJZ368QxBmX9ERPnS4mOHmhbSDXxY5fNEhy6/4B0MbjY
CFlPbsZ5KG3fHG/i5QrhkT7mrH2/3aEXZWIAdZqX3tJW5MKD0JNumJYoUukMkrckNgdnMBgGBNmN
WWt1RD/Gf1iD5zo1PT6Up3RwTN4iggPTtth8sqg6E0ibSBf+q76M18FyXSuPIHlTmLf1vRb8y4SR
LPeHxB07pVOyTArWgHLm8gOdEVt+7ISEzuRzPcbGHCaL4ph4zVr3fjW/3zEyiNJcKwANdq8PoMbZ
sbxS9d2G9r6ejgyU1bhmVpB0JlF7ioMiOBGJUF6Up5m1zI8NcMSjgc8aVea5LuuI1aanzPwiSysL
ofFaX+swpyeGZQduCobc0dN+uYnH3LTCdFGRLlLCKodWBwMJrML7vFLF7FOuCPGQbYdZrOCjIeeB
+h/6ZqaRgKO9moJDtRvCZiVhELY/06gXZmxQCPPXGgZmWndqnK66CkdQ9UQMy+khEzbBAuuV/6ke
UmyKfM/3xNTchVmvmAnD5Pdbi3w70zXRhMWJsROoGrK4rRGZi0naJ+86tJKPrat9HJeVygaeGG1R
Y5cXswOXVpr8lWI0T9lGLG1cAlMl7zj9JUN7SFTiT5xy5CRCJ9N7zMKo9rAqiFAn7/JYHFCZEa8e
mNSa9en9lQay7cXlh28mGY55GJfNOkl+5Ka4W2MY2DF25XRbV/pF6VAho/1B96BnqA4Qx7poH7sz
XxoXrRgWxqhJNft4uXlPF6BVH5kELjoTWVQzR4wmLj/ApNONhmT3lvhk1wqJFwAYXXWYXiMsX5Ca
aMrKWpe1uFbOXTaEmXtvqPC+m20qNWCjhocB6gnMVJbKmiLdChumMNlnAZ33ralWjo7hCorLnNsG
w48bjHj9ZUCAwScSPVzGixqDKVAUX+9LWXGMeJgs77LAQfTDyWsVfE6c6kHrDGIJWIZfTGbR6CYs
jHKZnQphhZN+2i7Ba0+Af0GsrUfX4wkV0IIT2Pfg6kd8E2WK/fSHJEk228yLQHwysoAIucTXRzZa
nqAfV4K5sOLzzJVys8FrXMiLhfD337eF0FynClozGxb550epfWbAKtU+07MoaNj7uUS8wr2NQmpI
W+HOSvGsisp2a8LozJk3+6W+Uebf68kIZIZ6T9lOI/ms3UYRYAjJTsjKSyTfrRxu3n08JkFl6vt7
1gWAmcv4ItBleSyFpLovFOzH0SYu81KoxyE8LWAXyE+r0AfrejfS5JWGY5JQy8I+w0jrMFsK1Lwk
xzoKlOSLaa+DNuynbzxA5EPNeMs0r+z/c+hR3NOS/Ls7xBIPVwIwFJ5pJOAHLMtDjv31nYRTmRCR
o0wGTrsS6qJRDxawZDb7QxdLNM2zdNU9zbqxExdbHSju9VHeogQRCWPQ+yVFE5Szqh4WVC5dlG37
W9zYSMJFYYAsFiJoV7dXCLUSA9HHGrX0LwedrO7Sm5V+D9q4ag9T7qo874I8rEWu6pnRn9JYPvcF
mpQctA03ntDxOmvzhWBg4JuUmZ3E+EPqnipRCOIfgTjNz+MH9L1BI1yAV0Dq842RgHgpMpVkLzCy
NehxfI5PQ1/u+aTnjOvF6UowcENQkiYyIqgZhHP54cxvTJCeAXOVE+4J6UBsQIfmMnfcjWb9kA9l
voSs47WIKXe9Hsd7CZmP11egqX+ZwBjtu0wQgd6KB9dvTyOpq/z3lBX4ET8h9I0/oiUBZ8fBexmF
J18VZRPCDwspSw22j5Jj24uYxRSbWPneD8YRAp1HzuU7DKa5OEfvRxG0Up8Yrka+9GnjXY3Qj2nt
NKD5AwjI7zYP7YAEN1iJxQl8MymK8qNIGG848ewkoPDpio2jnK1muegbEGn6I9KXmuEpT77kXccL
AyYp1P4EESUfoLyd0o3la51Raouj2xCamm/zW42kwb5tPO/l2p9SQ9FjyZAG7bBJ4VI/+OfMH1Bb
nSOE+l8X64Kn78/mM4KOABC3bhoa50FEeg4VnyZH9NlVDtxIVOSrlrKRS1LZTYgEpFWfBcodXI3I
tkad897VNGDFlAIvioICTppY7MJyActDD8f/n4+5Vk/gZSAQCCjY+tQhKsdXPN8UT89wg4ZygDyl
BuKY80vZ3XvAs4vAe7G3D1nT62Qbn/NWf08z/4li/MzcFgFB0+YvCzhcnFmrze4Ax1VFL8u0YLi6
1xonY2ak8SbDmgBqsIzcK9U8tm7nAtJwK4WR3jkI/iiE6UCUPW36EngGVz95T7EAcQZKRlkxN5HW
Tqq27Wlycwe1xllHinWdVp9/mq35rhcoKuDfJBkP7Lm7YJoOfyMA2+M1qlQG9JaRQZ4kCCyGkm3o
IkTpu3E7zU0jPN4txQDh6Xq4QdB1zRGjOzCpXczS8ywZ29/shYWGYgrL2WLAi+QV2CZCa1xipMV6
TMBdwlJElSd/wT+ZjRBA/lJAI2NCEp8hiBiX4Pdvo2Nm+aemaC+ysQJW+67x9drfqEJmZIUFhTwI
dbkG7mWFkTsGXTLd4p9s2IonI6ZEcecEYfP+zIidUFi4g6JANYR8p+BLop9613S2S1qyFdAzzneJ
UNKsaRDkHQN9+zQggMm9Y8BX66bCmcVzH5wBBZj9DTyJVxh7UrFtt1J4QEBbb/Ypao0NXrficIol
5hblcMXqx2cxxtLLy+yf7O6PzAOcCX3yYKdAObvYXveNvOahS65Mtx5+ReXPL8YIZVddHzUyt+ND
UhDxx3m/7XtoQYlh20rIW8VyhBiiXz0fc89nhu/xeL0fFRWF6PChjozxbRosanyPerFG+vCNq16L
RVuF1g98R/rp10sXskYBjfuw02hwT5G32ipaKVd+GadE8wgEf+1+Mi7u5rMA+S4rGi/I9MrN+3vI
WNABrul8ADRProHlO+BonBP2XPv/thskq0f9ghwFcUvdVCmvRefTRv3OIrGwOwZCrtyzMr9E3BjE
CMM3ENlw2JMX50AXHhuFMS8qvvqeFCZ+Yvm4wsxytKp06FseeVuFB1RmbKv01FECYU66aH1s+TMa
bTuQ72k1vzDkIqNiCh/wH1KYSlf95GbFqO2XImh40rruQLqkK/CsSsLFbJECoK+dB3DWFYDUXId/
IQNpGVK5gc5mBEa8XpL0GyyUFXSZ1uQuispWreCH5xY8woXjSmyr3wLw5FFVLIRk2LcHOZfkUuBp
bLHUYAGzXDufZUq3HEEZ+nMrrDV3O9gL0tW76OMqFouZMZT5mnMDzyqNHobrVYhMYY55LfVuAbZH
uNCQoN6i3ap+9DPHJgBUVJeTa6ERanKWaM0zyiqgKfzWT6xsVAk/q7tWPW3U8DqXamzIlO5mZpuL
b17nWuNgiSjSzJMG+1P1f2jl73O4bIoewM5ojAb0ogpJjk/cKsfmvD/e0k4cIN+28raQd50ouM5K
5HJB+Gyk5Ee5VOtUoA2diWV8geUHmFFuxv9fLH1taY1Iv2TQqxE+QeYUiQ+DfEMMDXNr9RMisnSx
c5kl4CqTMXdAg5SwAGd+yOIbr+AdDp3XBBZPUfncx24rsUDD0HWoRQ9/Zx9lEXghMKyOGaBhhuua
ornmYyHpZ2CMXG9i7H2TWlEDM+iR9CZ9+VWPVNbCWA9ADvltzKKFWrSREVMGRUz6zsYdq+ynJsbk
hKuYairttjQxh6EqyrQxhbCsasGabgarxjSQ6Fla/tSLyygKkdHoTuU3nLG1kNye2fMn3WOOKQ/C
eyjcisAjmiwJ6Zv6gg+zhLIvgmwlTxGE2qpZGkIGg2CUJM1Vzu9nDfNjS77Gqq7x8FYEc01fDhvn
X2Ir7wBUv6Vg9sga6cUHRu+oSY7GR7rc3LdWRfgx8AtNRhlfS/SmFzcq/LRT+Up4F/LW7zXP2uW2
c03qATVrsP6BpxvunnN9NPYifk6ZbnnG/peB/uM0Q0Fw1GPzDp0U/hR+qv8fR0AKp6jovV95SZc+
ZfOh4GnblRDkwyliLn/8z55SX7m4+o8rVDIk+PEIIYcpXGUU47vxMw4xcF/WHgSaOJpqyVuN2+3+
ZHsLiUGnEAZV5hewpri+Ow+Wv/ynb4leAmprumko6I8kE0CrnwNK/Lneeko8b8ZK3mvWmyk8amti
doCRVHuJlVyss6E7aWp6HaL5h2vStxu/sYLNzgPIdwJb4KRQXys+cd6JMymivZ8d+YPeTAtlVEV3
LBcsLGZ7D49+dPQFw0DxG8BjCZYpZUh270NNIhG4vIsMoK3V4U68I9YQHslgqLgx4TQnLmVKd6b3
3gj7/eeAVTJ59OKU29tQssVDJogq4b6TwXBTnkxfPpP14wWt1P7NtVrcUl2+tMy/BfNpkae/fpM+
qG8IIwmmjEEYVap/p7h1dlh0QenE5fJX8QbD67biSCvoAEjxJJtmhRTLYh8nR9hekN21kGLSEcvf
+kQk5sfRMACkkEKC2GeAJfYbE7y78sAqi5ZHwFkds7CtOrvofabkCyEmisnkckuYYsVYqsWRciCI
qgtrEx3skkb9BdwXgsJ5SsmKaiHg16eadgxDzhtvWSaUlOnsDizJhjcWXSDMy/hHDdlW8CLcDQtD
/ZjQRzFbJ6Ebn+VVyGNzwilvHOVRaJSwyIvq+HY5zZi9NhFsNqxpwTF0cD0D8OaVAzm5S3K1Ip9e
VBmOPDWdlH7crhJSEnLh4Bz988xgdYWOnKZNkfvQn5kI1ZShI2cZLkQ8n1OXwej14hD7dRnQHfxA
xecq3oFOA9jgzIr5WGIn5kli5BB9OljEBJIVI/uQto9NzYN9xPBDMQGVyVVemlJwQlD+tgVOP1gk
McpCAGHubw4EGWlCtJ+mVqivwixndTEiJLb3IpZF3+mWbWdjVlRy2hfRTfg7KYVchUj4Da8sEoE=
`protect end_protected

