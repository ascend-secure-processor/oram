

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRspnG0xisfrWCuXYUYBfE/AzbalbiiEOGLExCcnKHs8umjfNxjW4sgcsMHtGuQTpAUFhLn9IUS9
9iZSbM8yLg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gxnx7HVo5Yuo7PSFF6Z/GKHM+G1yLMp9bWn/+/qj4Jqx+BYVQHPZ0enMcnZNyMqSXGtnf0+GYffu
z2uIgsnJG2MlsfsN/3vba3Lh47LZzPtuTY4xSCB+iWk5UJr85cbXGY1C1Fo5o/CUWFkRyAGiRoWS
7EG+S+pN6eBV5Rt41ZY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lIzlfJyxTW6F9GTtPoNWmI7TjXFsm5QCxohJUsWCpe2DSzOumuF4WWj2yWDlJMOM0XxO0wIGDFfR
c55GYbtK1548Rxfw/dzma3A1tULJ7b+qlx1MSWJNVGn7UnyOEFTB3tDQ0bs5eyWvkxJSc2FmcbF2
idLYV9SmHxTN6Xc6SfshrDcvaJXcsx6qj9KGJUOUVgM09dh2vWjOm4SP/y6vNdOg+GnxiMUz1lvh
jx/7UC6i71NxMVGzkFKeZLZFaWRveWrxDliLDgFe42iCHcW2+Uam4UC9w8Wlilp72tAKKtwqpseU
wLiZ6SLLRddAMDliioDaeCb0SPLY/f7Vu4cH1w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NHusfgg5D9uVsWblrZf3PgUBJkkrMCeV1YWfgDBWw48FwlSpMJS25rjZ1XM5BaQ+YKHXab87QOx8
vz7h14rO0vfDl0N7s+fSfcjEQLtyPguwmYe5jrbBUimkwpn2FjtkIRhltE2HPaLS9ewETCeXBSA7
yPGc/Hq+uVYHArBAKoQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G9hK0CoJaDSAj3kt/ff/0yHYotq3JnOL1xOsca3zJ1VcNkDX7e6IxBikcItdKZY2WVs7NAlI7Q/g
Qh1Ca+IuEScA0X2p3XC17jhyVPdT6Zn3IBgLN5c/nhxSXXmm7GYTToeq28kzOSUm4j5MhVg2d8eE
rTD4NTWQtwOYvMMwFIaXJFsD+GiF4Rs/2o/5DsS/Psglcp6iBpn9R7ToVcebbRbrq36Q/fJqlpkU
I6aNzRtYLFWR33thUCHOkQXNcrZ7fwQr/IMduqmEO4QQSkfYvV6DN4e+9tXHRfHU/cNKhCCR72pc
dYAR1rD07V9sqLVotVVAUNuS7cUI/ouitsRLhg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23296)
`protect data_block
JbSMfUDJgS2pfy7i1xdJKBvUV3o2GUvOg/YAAaybYR9WkYOoWsZ4btS9xWCSD4hIiLwhE5N4Iyl9
gCjHGGCGYMI79oKhhKnDr+vl5LSUF0++7FkdlqhEe6YREawrk/VgkjXTYPrHuwE+so3L9diFGUTb
rZbs9iRcARza9gxG9sMjXVUJwPZauoH6/eCn6dA9R6t7zLJPuaPreh0HSmTKnPMEMgcFbAkG85HW
QpUao79z0ARO/oJbumpTo2Joe/gSz+zRXS6TFP0IdVg1SSWNM4173g4CizBFPcNXZYh/2RhL3lqN
Ovzb4D+N7ViInefYP+kyZfkpYQTfpxGK/StFctaGKJEqxaRerro+4WL3Tpm0eMHllMt7nIPMGpM+
2rz3IN6nzLXPpzIK9g/RKNDvP0RFdi0epRvVMuTSCUEajU8j3xO4rc1iAWcKl06HokZ3y0YurpO0
Olm866MTrcmd0BUeap37Z/Xv7MGHpW92T8BwbG3Qgn5z1lF5uUZUx9+vWbyS0ZarjVU+dvP4QaEq
w4/8SdmVh1a6TC68M0aXaD7K25crLb7FxUw1BIhABDAOSNnNueg8am2VWq23ZjJUqNfbznND4jJi
9n2Jq96D3Xg1HwCa2rU2cxe8jR2U73eO5le5OGQIgqL08JEv/b1xoJ/S7/3WhIFdHBYajfPRs1Av
lgyrobPUbgR5UCk+Jkczr1B4jN+lMYvbZY6cuwiCDZUptMnMSOgZ6ntKOL1R0ljg8/H4s11+B8q7
xKfbhegKcOZfXNcSDthql3NCYv7OKIYxa7kG39C0szVWAIJLOhH8+Z7Kko8h+O4f+GEO1w0DPh8o
xKMnAT+4ojfRpGcC5EngsUpCRfWAjWq8cpxtxgq092Vtt1nDideRXVCoZ+SMxscAgh7RyTTnDR43
La588veFEj+zNqBEpvcUGZuRXn3TOWFvlSZtKlG+1XknvQo3WVxrwN8L5Z/w7Pkpk4bYrNslshiy
AGEBvkWDfb9qEL9a/Km0aXpndl78Tu8nUkY1bJad1xq3ssc6+b/JEvh6cpPe3NEu7aljN70sG6BC
OO6o28p/RbfJDSL3y7N1Poms7/W5EfXnKq8kem3T2MoLPAHRxQxDL/yWjIxIZ6W/YOGkSgKt0luI
lWPQuFE4QZ2T+bm8tUizcnroUQgujIP46yj1pNVYTxt9+gA1dsvUkS+kgHz4yupJHG/J51vX0xGj
KfPj9SjVNdyHOrLLUYLqmIJ59MgNKdGkuEPLKp+1UnpYFpSLmlZ4YCN7yEnpEt/eK9hiMV293VvW
HD1hT6IeAZdsM3GVWbs/gbMnO3LIQueFcrLUd23sR5I9EoXb+BUD55aCcVYPfvW3FslIqqOLyMgz
qfJ6ma3SEIMPq/QTWJcAte+IcCI7eXRUvP4R3YUYxDkL1bQSFQBRWA7/3c/qT9V1rrVDNyX68tv5
M6tDTuUdOklkwM9glKp1NDFldwEKH5Luza4/LI0KlGFmBOAbCJmoAtgVpUfXkrJSlMcDdkuFV+gE
Cp+zhHYSEqFrpAmIvJydPxTWrS1rgUGWdOhePrv8gyiWr9ShhJFMvHXit51jtymFX12RMfyKO2lc
O/31NUQYfRaaBj08Bw55yw+zDvtKY7PMefcOHJqwFaHH9ehM4Jt/UNBJOpTIgSOOxFbrPdQhwDtN
oJRtdoUJvb1Bgl79cYjY5Qhc0r6IV3NtgxBj21lLE+hmtW/q8JHGG7aGn7LpY4402Ufia97jxmc0
Qp+tHSBFarEWJdppU///qno9FL1kaUHu1PMHhXU7oWkeq8Z50QH5HZFv3XIiEytzkYwU/RuHU36P
H7M7ufzQm9DYiaPi4hZj/0bLb996zwvVK5kFRO9caKe9YPJ2iS24Wgcjzl+F7ec4YF2MK970zE7W
uxLCPe/3BSIUZdxfIGyQFRxe/Wyeb0AZMsWgUdsJKz8qL1soB6f1dWoS5xCAKo79Ovf4F9FtAh53
7JHkIC6Lta+Gn74zwnqs8TAPACqnMTeUIPgLbvVv48UoCz9ut895XlOBgWe0dko3GW4XqeSAp8uL
mFJZ2Vw5yoal9M2dfBO9MJa1XM450813IKuDel3bmOQfwQXHcOv7pjDaSTmc5r0u6dt7UV1cImqQ
66DcmfXdRRHohbDgr9tIPQOuZY15vUk4R/UUEtscIQ0IfJVpLNUrEAlOB8LxwCH4J4ppq2tLGnRG
lCvy5DVXpaXrV08yWrquo2OvajsENvNhxfmlypRRc7BfE58wATaN9ygYPIr88u/dBJJhWCY1rXWb
f3ScplE2lstVMbOlGs0rCd8U3cNJCXuUCFySwZdWYUvDbB1A8LSAKjmGbM9517cjCEvf8ra8aZt1
zgHxf9mJhEzdGmZrXY388ZB3wVHzi6fkZfSKjxeELAQyMn+KSDlAid2YMUTa4SMy/zmOVR62n9GU
qtOOq1qXmdY8TSJSjSUeaVsdABH/cs8y495Omr2UaPhT0o8Glss1nw38Zc6DSdC5t4IBPCJ8RumP
hS4thqlHN8nc6tJH1eLvxh1jIXOSpCh9e2hwEkFpGD6NJX8oJVceNtMtyhI9lH3ujy5UDtyY2ia8
ENHZDxrXLXvaR9Va9+ujhx1gAiIRw7NGLm8AKpS6lh5Z8eDrHL2yQhtmLVuxkD0Kqh2FgUoSK6Zv
PvxRf1atHlbZ5dc4jA237UVhGUUO/CYW5j8YgbBigER0nIU0ZmGo8P9L/aOG1Ldos/ETNdAYT5rD
pipnDFiPj2fRDonxx2SwOAlwAlo8ZTJu5MVPXdD5zGYxJzFzyfpmHDHEpG/p0wFWAAopJrLBzA6X
i12BVbiJP/Q7l0Mlrl/OjrZehEaSdlJomKAb7/OYOgx+quV+Jd/llaMZEpPoM1Iv7eZS/Rmuif3m
THdRdJGOpgDomphgBr9rzkprPJ8OIt1TS35u3sIWMKaddQCYMbb72mOJO7MhYUx7CUCZleWLngvL
yFQCOq4D8Uw56YOrO2kFlXoUHHgqsFubFZbKCHj9Fa+aBSJR88t9Bh3MsmTfbFQ2KSHTI/lQ6D1z
pjwxZrtfvTF4d99uM5wKpLfPwpyLuKMHtwetCy6/2T08eQ1NgucTOWWoFdaSLZVTlROC8LFODkEe
OoJF3fbDR3/vF5J5UtwXf8zCP+PMyT3dtPBadn3ewfDgHUCA6V0zT7RkoaX0+KquZl5dJfb9bSm4
SFbooik8k9K/7pzkCHkF0nqACo1aXjGN2xol6MU+Ordo0ob7s+6ozgJxou7+WDs7wAgTEoKzjYYW
MJCGifR6vCwL+KkjS20zVKP2G8FtGrq2lqhJbkw9DvKMxlpedcbFMb2VaIrzRSHPD2HK7YscpHKp
M9fIwb/zHXgQdQwnLq4cNCf2fQiiDqmxIz8Bi7bXfqsczIRdtecb2zNiLnPukWRC+NJ/5CPq5j9a
Mq8+QON+P5x0ihTvbcEGZ6N1r30brEl3uDBK4DuhNw01yAbeNI2uiRqNWbi2Fa3wHX0SeVUcjFCZ
7e9bXSthfm+aUwQCltO36OE5YOOHhCQzzFsvIKZ7LDQ8v9kHbfE7fl2Cb5wZSvELOyi4jQJ6+UB7
tygL5sOKjr9sTKy/sSDfynv4lQ2UKr+J4qXGYDGWpJ5gYFutlGWvFLQguUO15IWu5BRJnZNd50W1
AJQJCKMg5rPN8ZlbFhyOBtK5V6oK7rC0URTbJCdcCRkuskgkFqxTVa09TkW7hdgmxs7pH2ez+Jg7
WQCHcJJyXMmnBpaN1bSCyu5uIu1roDLwq4gITJcEg4v5pBXlnhXI9KX+3Mse72wd+2/3w7zaA7ZB
Tu2GgZNW4H3flOyJusCMFgyAQuquqawnV03Uj+eIHscIC5kuSX4eArSTEtKwmmxCyTuRte2TIPG7
RFUGX9Nq9wUi++L7AgZOlN/8y7DsfNJU8IRKx6ZpDbAKsko7YjFmrt//fgUJHbdtA8Eb67bkQKUq
JGiCnEKCgif3xZZUERPEW6kFyNW4R1Jno4h+EeInrd8EXRugDnq2zkqJeaUz6/1YskAvn38iDIUk
RULArwkWruRfj54pRnkrAhPh22ATk0ukEiLqqNxevJ8b3XDGxNGCIGwdIDwfFPYlInu4adahpL7P
sOvy0I9dVe8nf5jbWMcC3ZPcSHA3AoMwIYl+AWcG3W/6MRlveJGsdZFlXxlzwECCw1yekk+wsSvm
aLVO+OBl1dsUWxrks3IULSS8Ct7HaNmxH7P3pKi+a/rd3IHsQboq26A3gstDBvlzhAS34F9V1lDM
/VYDgj0oZ9xF8eu3P+MIVehGvLJtbLFxJx40Q5I3HteLgyZw22IWqRdYo1dSeb0nkc1ONQ3Ov329
oMWUMLWi1k8nYsjzPKS3tKdQpS0FlWp5cZL0cKnVZ97rWuHhsDeN23qSZn+buGK81f+HmwZudWY8
DJyjvQJlp7jZm0WRsQDLX+tefSadcHnv9IERz5ZnfLAFlrKR+Ug/jOztEpNDc0cSCEY3vH5iKNcJ
ufoCcaHlSPt9rEaD7C35ER9hjKm7H9k6bYZFtHL7Z+1BMeSIbf/op096XDvntMgrR2zG+QxLSVh8
w6hZGg6B+x1rYgqceSLkXXU1vs0KI79cv1D7c+Qbru8/nOVnDlcq8IzvCzy+v2Uklc9imT6wW1fj
+tiQlVsDoChFFWxDplw13Cllu52Miq36gAqdypx0c9mmuSRuc4/MlYePV2LCckMEPW8KDYJcjRwo
ULo3a4C/fjgi4SzM0edGqf+x3YaF2ZvzLULXR4ok53sJoi6NOh3fohDaLZD/+aewYX4H9v0FQWLM
nMav9PUJuSkHeSnzjdbAoi1lSDge5+17Sn96ESHmzQZLJQbBFqFM2czVWNyBiwjWv/m1gWJXrUZp
QtZB+lPS+XsQfrQvsEPsCResEESfJfS7twK1npFil8tTbb+CVy2FfVOj0bc09b36SAGk/AN8gmVn
EpWnYtX/lp2pWpgoCwZWwmPjCd4AAF3JLK1Fcu7tTrl/BhjFpHqAB/tV1y2KQ1AOjMd5Bhm5ITn7
SqAYb9Xrlwt7+lIFHFc0ipZ2Iql9VJUV9uznhGCR8toz/vIepq5RDYeNY+AXvY0rqnxCE2zB79oR
i8rtGPk9czPqqjX967wr1VskSccfEGGdIN2F7ngk0x2/pGVLWKv18yGpcnAIpqbAJ+5qXNVrgOjk
B7dL36FbqFTbkyq5B9ntwSRtGragplQ5BkXipDhXmlF8F9eb9ahQHHenAI259bT2J8BLfq1/SH9f
WGGSb+GQyIQnz7heuMQpFC/rYKeO2aavXPZ+hASBA4XQ1s+BrUfaB2GJz5QJSbDUuTI4tizAIcf+
HFfAZ0LInWdRLwsXWAiCMQWmBMUKSF4GElQBc4I45fGHo9/znElY2b0S4e1i/LAAA40Nz54YS+wi
f6K7arm/aSifykyEyNBVYy8NcyAWa++PBjzRtkLcBc00CBjtfODWG5tXevwFY4MhIq8/l5h3syjZ
imKpnmAc31VdY6g063bqn6/S6ISu2d4yiYALCfjCsD+MJDc4jAtPxPKYEavtl0KlI+ZmCAWjXaLX
4XJ1ZY7oSNIL9UXFCEFAHymnNS+RV3XH+PvXqZkr3COGT51in+Ov12YUuzgVeKRBWDn/bnnKKeg5
aJ3NNTZr50xiNRP3jZLg7N8lPLC3gbv5L7yDp0cRnZrRiZtPHhr/H/6ZiksUby+raqcjHvG349sj
nJSl/wSDsEPAUByu7HTz61uGa8lT+nvYP5JmoLoTi0tuOy5mDlsCHGcd8QDVqCxMRNdDELwlEVgB
cfzm97k5uBAEsI0fBSJnrYhHtopy2GEBkoOk5JfdqcH+RO5lGTmJmpi1eUwYG5eWm86juTNXb6oz
cDdHgtIH2zLlhFJ6iR0JGF2YHU9M9jOKNe0LgEZjGPlMpwjXzERDwRxhMu68I9qJ3mm8O0fTTQde
u5e8vE7IdAKnwBj7pMAisCNKVXIzIdG2iRxQW9wdvCT5oUSd8sArdPeyqTlzvWkVln7BQC7r9X1f
s4LsOfnv1LBgXd0q6fNv5rW3IDbxzrA7Eqw61/Mm+7yzx3dDKfS7tHNT78JZWAbakwl9svCMIKe6
q3dSbF9iQ+S2EjnteLjLsSdS5XpWgQJkvP2bMv3HcyY6Dje2R9dUfqsRyWRemTrMPWk7FeAB87Gt
2WSgn+Bkj519BbLgsca4RP9HLcHyQZPF1qffbsXUzAYtY60Of12fQzZWq3NqIVqcHfpvRAYZzJTK
/IbXkFAGbn3mc/8CLbK0shJDdmelqtkY1WSluWjfzTAZwQp8GReHbjTWkOFNtonK4rCOJaSXAIFP
5oHZREV3W7ugFzGmkutMNt4ZMU/8JTsShu9Mc8RT7U7J6SNlEa/4GQmcstfOqsnCZ1gm8fJWxgW8
MV8eyNf6IHtBtzJKnthVFd7xGvjwqi8L6memae4XbsXY2msMjrOBGzNhMcc7m3I+YzF9xqI9odfo
iJn+nRN85t2SUX7Cx8Cgrpf4RGuX+OQwyKACBEtWI3gLy5oju2+4Js8Mv91ZH3bgxztDtiB1Sa+S
vKiLOntZ7S7pa/ly+Ngq/Sbla/2Obw/VqgF7oCCbKv5bCE8Mr6wCUvBhOP3AQrxvfk6gQQ2hvgMX
+S2IhBC++WlLX86WPIx9MlaW9V2n3yRmIHTjOym2wcwOb03jOA7goCYx2tIQeOp9ARdUl49pU41P
2aJdSdr7xVrVBn4f/BiAUHuqYjWW+fm9PkQrrlkZOCXpJ8mVU30zy/mOLjnZUOwAv4dUfH8fozWk
yeDxDeEeayQJCfU6GCj4OFlfvOIiNn9LRwTzAMSHoslSdMvYeNs2PaTigEMCX2cUz8uJnzrJ+QOh
vVqlazvwl2hMeSV3+huugVGgZo/8RvoEOyYxqnT+LTgtm7AB3gj6cPyVGYkYoGrgU/NSz8nnk6Fo
Fn8XInNFeP1Fk+nuI/GoCA8zMcBmePZXt2nuqLh0DxjRyaJ6l7mpwyUot7lmmhkENWlYCGjYzyJH
uMXjG1rI1iyMnaq44KBi4+4ZqvTbNxaS8xPwOhNQ+hTk5fn2oHO0lUd11HWhGk2LNHL9o7DCukaz
sudw1MBu6mxgIWZTfmPLDGtgJbfAE1MeRyH/++YWEd/ue8nUk/C0Ip2mIKoE4kzwGpzFFK4KdHRL
NBFzqfqwyZVGLduUgDmCkr0EOw48+J/GhFZzQulcD22JxiKZ/Kj8CZAfEWqKDEc58enbzhXHwDBe
9Yko10Ddp+Z1SUogzo9RQVCxQn27aaZs2aq7S4zTVSd8xrdr4DncowgqOI4jqCXl3/Z6cEOEe9m5
yGDKWMiMgSBdofpBR+TKwF5ykYIEz7OcA92vLeK7LJVcgWOj432iprtpIjBaTAz8YlRUpXU6L0eb
b7LAAHaJi0Vow4wqhK7pn1PVU5wxzn4pyorYB1/A4DH9TLrySzyXmG7/NW919U13HuyRCl+7zBke
HPj3lKbmT7DgG+QY1lHcQw6SVgJHINuaU+zVyfjt5aQkmjCAmbodamvuF17YWX/s51ZfKngp2nUw
y2cGq7QOcYkeeb4v79bn4OyCW1nb0+G37LHuo1j51Le17MQTVoV2wJ87RdT9PfQGmItp14bM2xjk
c8CH6mkUjUViKajtjg7H+LPh3ij1MAUkV0gy3y5mD72IyMrlDy9n75qXvnPb7kUOAu3Vf285YNfE
mSd2hkURBFhHLBsMRb9hCDPWQqwOx5I+7WbeFSRIsX8QUpbKUFD+YcNdHLo2mDgAdeRGMPttLN6V
6WCncQbI3cbTb2m3lZxrY0qBdh+ThTCpy5dSgaTNFojdFOhzGsDLNpS3cVzNfJfws7Of4jLP0gvn
flMsczNkyVsuHff+yruP4/0/CotN+2+4pfvNgoTU4BqB8Zua0AmM+F7d3sHhI0+w7vjBPB1ju2rj
wTALqBXKR+cpiWL4rKcyI4YSKfb0ZyeCJr12n9cFaogqK/4b6dfcOCCQ8wjpuAmbO/wHUGMlEPN2
kPmJ7UJwYsaktqJZtTTrqw4oQzPRlks1FBfXu3jMvBOciKXHx3sdZ1PqSGCXYYGqyenXOD7VVnM1
f2iwj0KevVFAdWNrb2bZFB9IN9AeiS33eMFxjEJeTHPEOAGKn20+dcI5OGpub6PuFy7psF9CMiGR
eBbFn0V4Qy2D9nJci9E1fJzs5iyGI+40Fvz341aE/QuIZwweFmrdfOOw0sPmEkNYfJ0jM4Es8hZV
s42SZtVMx8RswnfjFbJMMUPvR/VvX7Uwxd4Fski84S3XVWjTR8uhBSHZgmjiFsvL2ubFa1MU0uQY
IoKet3/GEkN7uu8AXcn8UX//ySLMOM2/GEKYzaaQZ8hely9zvG5NyNbK520dYi0MBC1Fw4w3YGCQ
VIBVx48VDAptjes49R9+PdYhtjhbT5fmYgrYJNu7UkmRb2GM1BFGxwpb2xYG26zjHxReYt+1A2zF
7Ou3JQA50ezXsvB6AXIvvxSFhoouW43UwxSXUJJj6ZoqWy1mdEaDPU9AoXleiEx0u5JwKjcYooNp
7y3k+sT+i102bQMlvtquA4dTAXbIl6pHV6RUFNUyNtatI+9vBkXXkZccrNmdTb40VB1fJ5Rs1Dhl
UGShlPqRxdgJ0nBS/mU/wJY3gZKhO3IXIhIhL5mG8mUxgZWtglaSBdQwwdMZp0wF2130t6dhip5Z
Qr2047edWtW5oZe6/EV05ddQ0V+U+k22KzZIf3GkM/1pQUQ3G54iEdXxRTHZyKdAUwJ+DyDybIJF
C+Z5ftgpKvD73vvpdYFGef7jIVEVn+Yeeuaj4R5YqyiS3av88byyh8jWliPHkojwAv56/BWtRIQP
ckONwJxLh8P/FpURJhLggaiy9liiASWkkLjKqhzy1FOrCGbDJiUaNXqmZt2YdDMVoGIGqKAVHD5Z
a4lbAKjfe5LlGpnVJ/PaGspqe6EbGcXu4gwWlWsX79mb7v8nx2Uy/rD2cp5EZLx32oK5G+YuRo4C
Qvj+y17ypIbnnIpDjH4q8262USwkGe5GFB1ZMO0ZjYJIorgm2I5qjvc5hwmq9Vg17QPuDAr/Xaoy
unZuWVt8KPtWCGBqBo2Yrmb7ngCtiaPeKoZeyEBAyj2CJ+j8wENVXy12A58f6NaHABz33XNfXz78
k/9XU9j3qmPZlhrjvqnjfFegsAG5c8JWy2MEf3wfTNrOpXHrXCqGelI4XvrQk4cIDyDPi9+QUl2P
akGKsn80uCgBv4WkfVw942EAY08e6La43nMrbfHvt9BovHVumqQ7lP8Kkp16Vy+bUpX+OFf07+LJ
p92VQuZyWFbkpX8yGr9H5vB+MO5so84dYVVMWsIBHY08A8ieO9mUY5dpCtbwo7/oZ4mvPgfG3NEE
DRv+s5Hi6cv9ooI2rbNUipAFlnGwq2ti0ahVVIKSQgpHrWQLOcqNiVPp1NUfPj2/9GTy1F70cS3Y
XiUfg1P/UnVEX8XE/20odMh5YyupLOuE8QL6uzHXhLUMp1oWiRTO0oHANsEGUO4Bdf9EhXQuRtVj
mJkwG8weTDoqSU+SpGc7gLyuS9pDx1hSvVPbMkvl5Sx7oguOMHlOZ27ZPw3BvJ24oisxBoURAQeD
PHkXwPgmsFh4+/J1+ahd+dR//4BHfE8ffh6xlzoKN6jJURmVxDL0c3tVT9LXPUHf1gKBHY8v7iMt
6AkciWIiOW1c2xsVepeCNPHdMfn7yNuv/NeF2/AYwYqc3KqpHyHYXv0DVwINZTbvPECaxJPzB+tN
ljgW2EBHlhHKPC656RBS9d0kKi2rHZJfPR0UnYsidcGx3GwzEaPoA7kv42Cy3DhVtoXYiWj0NFTo
o0a5vR3Rhvs+beN+78+F5EAlaerXUVJHwhVHeUTwk+aadn8/1mXFZ/lw5icvX4mNq9f3nu34gB5X
tMb7ZxUkHzP9p8ZpENDovtsP116XzIKcry9s7DfyIAFtJokq80dgj0zNqGL33lmm+wYCT4nMDcIM
9l7ufzTLffRSuU8ebH8GM2DKhK6IcWOY3QIWzr78GlpYpLBhd8cnhFMknquXBJUqW4KAFUyKwzL4
j9LjsDMByyXrvV2jpiN1OakLT+f1kwjz0+iSDCrZ8m+D7wxNoD7cK8CUVcj4009Xhe9WSujksKZl
W3WKlrX8Tt0f52solLOsRcUUU9aqSjc0Gk+L1m7hBOYhaQWnob8coG8zgDKvUFE931iZQViIypMd
l92nQEEQcvqJu+DhFZizNxH3Gj9629h/62EvHZM/h5tfCNJQFOMs2wh0JNhImX85Le+33aY8wKhZ
7BB6cKtz/cwNIN7PcVAAlKSCnFf2rjuieKI8Ow7x/kO7tPSEDKPP5Lu5LVw7NgmOVH0HPCDIZkmO
IZgSU1rXmEcHrJ7k81r/14VgEJFaJchtXWlu3rdcLyJdWd/Boz1mnnp/GLRgg6WJploSzapZ7F/y
iRmcMo3k5gglIqfLvOkW9MGchmLroMMk8ZeHdRjd0tmt1lloL/1Kq45bSzxfe8vKvQBfa1pubfp2
i2YveOHKjxj3AbZw82IzB81UyPtJUSsk3b7Ld/bfbyn3ivqnsw9hTbBEpHmtzn7iK73wcjY0+jdi
Yri/vqpV2m0fpHS937sBm4Zgl6ZvJJkWiB/05m+i1aPpnaz8lW9WTuCHxjzAyg0xV7fM9we9GFec
orvP/H1r/yDNaV/hfFtKkmMx1D2GthkrTyZqB6nSr7zrxjtDRV6YM6LLbi2ji1S2dexAYB2iMQEp
cVPC3+XJ2ecumsoncuBQc/5eYNTGgPq2JmGEg0m8SoH3AFBxFJvQz3T8t5mAdhRTQAkPUarNCj+y
ApnTq8AC0w10R3NUSSJxwdDvRsKFvY2XA0GIsDnu7WgJMPCkJnqb4fspJVoY2VsLYONPBLSCDFa5
85dJkNPeBy2sTB3Z6gRWbCpKcIYe7yx3ub6Cl1t0/hqRKJeePqMsi/CYYaaSy847dW/rv04Lo8N4
Y6SzJsHqFybK8xgaOu4H3Jku5xjc/8Q21/U+4QvoAIPMOMIm1BJrlx16dHSojZIojqOUga3m+VfA
oCzHiOgIqnKAeJztaoBIff9hHe33pUJePTclzV9VtUnpNmXZIP7PGfQE+/zBJTMZpccYF+sAv43t
aCOdfcnRYOix6d6pYLckvXEa1Kqi/JJKM+GIVPOG7ZHQ0g1QDEV/3k/HkGOshkfbl0bhrYsi5dDa
4rua1w7HM6pClU9JDLoOd5a+udjaQCJL2dOFqi/hrWJ37bep4Vti7XuX1vE2u+XPJKuDP5yKd4BK
6hWw5JHqrks2en7Pxejnif6tZ4hmiWmAv92iN3KBKStN941T7zoHvhD0SD6NSIgMlRSqG4KKlkdI
TAxuCcUlIvA39SS9E4hvS9pd9BJX6SIo8Isx9fNYfRm+l2bBDVoci6iwY3lkcG0PgVPUhhOCWlLI
lRc1b3oAMUhAHUVPY64iFa1b6126C7Z2yYmRcR9mJKNe2bfeG+XJZUwaIdkPgYYbskHnDefZF3y/
t4qnlgjvnw9E/3duAgm6hi9dLsXxa3QPvP2by5FIdUTbTR3CjrmS9XbOTPX+aWTk4MkEevzKh/0m
W0Ahek5l4W3htJNbVf+oaLIghENcb2JC5GRZ7qthTCjUAA5u2YCMk9JwDFHcELZ4RkMKGZYV6KIw
3dQsE0xDciyyKMAegYpF3m0QQwKbP034WDurWrIwas7eaPmb1yuruyFwdFetI4WCOxXUKlQ7v41X
8upazTeRXRwpfIbEB0C12YHhHNikPO2gMMz1m6Ac2OBOh8y2mG0vchwKnApPYGzzAu5Rs7jeSqqv
7G7Hjuwplgjrm2q9a72DTLZNikXrJvOjBdO+jClLNvLJSMbdroURiFbik6SEB81el34bGieaXWbo
9/EzcU5UlfGwGAoNS1Jt7IlfqEPk5wR3nwjqdYXcgkCikoj6COiUd7zMV79P1UCG1JR4Efvu3ZhV
sg/Yko5tkHdQKHanYMgaRog6Q6Hjz1ZwnrglC+SQJ6u4K1uU8jeqyJJRGjZX2uoHM8PFDmlawXJP
YTgDHIFuMvo5Rk0GJUI8nMYtR6YX2+6FbvLUUedRO4mBv7S9R4P5mgq92BzYZVJSMDrBnnRKdEFM
Mqtz5VOaOBWHj9AcS2w+0Pw+HwWU6bW1YNBgJybY+OGu69tQppxZjykPgrCYAZw1cAXIEaifTZGh
yfSvQ1ewmd/UsbziKvOEfHvC3+dc+Z1rqztf/dXIJXyefZC4Xad44wketU2PvcVQWOmZMkvtVAVY
MyeB+br0+TFO2Wi62capfcIz4he068hIFkF09b2zEaco2S49XIoc6dBw6bEl7V50Ohe19+uIuOaF
QTCOOfh2xB/BVuM7cgFzBXvWBAx1QgzFGa462kuO2lky3SJaZDGeiggGEsQW3IW70diOgMOuoqwt
WlxcdcuVgdKX16JS+QhScUJvaqXjro3r9dG/6mhmF93/BvBRBCBqezcjwwK0zQBRvD2byjPu3Kxn
J6BuBNQOPc82CNUkWUpuaL6PLEh9S5fDX79Gza8+Fa6pwRsYxQ6X+JXXAsHC5FtIsd7rc3hrtwj5
/L09en1nHKXsaP/fPxOVEYVhLGKDgs+S7C5NTEotVJJQNmRrwixaWBw5QJqmRbL9AySulbzM9lZW
BHdIScrY5iw8LIs0pc5pLRIWSkpXIaTTfiPR33nf2xQjqcXGOSSyfpylAGm5Br4Y45i+UfEbA+4/
KXel2wIQE2pRZ74cB5dcX6Hv2C/ljV/tcaWL+8sKTlmT1kygu87GwzfkKEwUNIm/txWRhNlzAkC1
hR++Mzr+pBzOSBreNcn6CYhCrPLX4T6GZt4z3EsU1soeOLTgGgXydtspor4OylTJjiiFYDoWxyHJ
h3ivhAb88CU1Pr/Ucb0Pay+4TG+OOnKrC89YTvaoOSEpqoVH5sR0QzYhQSpPjKOkgKxy2FfAx2l8
SqDEAASitUSTrguJXiQVM96MdzolIKO6ynA5caqfoO3gIhzGbC0GTorqE547rHfI7aA8nioJavPO
VIoY8cmjKjGH081DqZjOfS3TzpjVs+I8Au7E8+FOSsu/JFgwdgnotVf7Z9ZvwEEnVGRuqQiV+9db
V8KPR5y46oHsvZNRaz5cHGnj5vrlELmyoNfr6dYScwMliU6um9FMDPEH9Kyme/yl1vUZmAIlyFJe
LLO6yq2hnYUfW/88kVWmB7Xoan6pIuIR5n1uBtb/DtoyfW2PhgaJ/R8y1WJzC9AAdB+QQwc/x0xR
AEzt0EwAvdyLMpDQvT+UXlo5JSSNYp7mLTkfUYBBoPNxbc43FneIrCH70OnQSJgh7Uq6MmcsCOVL
bqQK1Zti9azxFQ2og+EOwerjSUTDn3ACaHXstF8iNQkyyrMzYVYqsfZpqBcaWYqNaUXC9dHLQvG4
Lx2Z0e9c2cQZxPYjGA4pXcv9GgQkx/OqIHSWLJpGrBGQOqT2FWZNrXzoMG8z4rTiPpyBRUBk6cWR
NvlwU9Xtat9xXj5QWefgrSbNdcXrCIFueq8q0WG554V7cif4EKrJbrrBAFyyDFaV4BE1rNfxBmgv
wxhk2FdnwnT5OqEHXhGgCb1GZIarg89hxM2lTYX8agUOwso+srcP0CJ7+I9DsMTARKO/X4BPnT8d
MFd4m+3lFUsbviGsPuLHmiZ+q3psSInCL7aWSnwh83o1wddEfpl8MEI8RwikQ0BWLjTg/IyjRZPT
AXenFHpnICt6OO9QSxXPeJR5nAgE2Eo0bXsJQ5DovaYHoZkgZANiWLwZfzAnW4Bpep0CSBwadhkv
puLNRKr5Prgrbdhs34xNjPHNCxp2zQMr07IKFvh3ArhsVbVdqRa4GCVH20x3089TVXLx20durKh7
g2SyJbqwe4l3fEjIyXBstLvMwxCxq/t+GXqHnUYrJgRtHUBPAW2nupW1uYpJe7jzFBxL+88LvnzP
VOpYrCjZRrwFwTHHU2u6ZAgRamIEpcHkQ1rK9VE017K6hki0kcyThVtRNORlB3dm391mEfE6YSkH
TXigTyzKIkUxG0opj2OSxZQuLkgtfI41FNdnUWYQ5p4ADs7WiVotvs/xS+aDm0Zy271ReO273PVM
zEXau0mWc4nM4r8maEvDS+9Y+r7sLlJKZTDT4OQqZCtdHbjD8j2Bz8wGnLxgTUaKRNix3z0kGnZq
PLtu8I0qvNkaL2tX+rUrcEUKA9XWrLerWQ18irGQ8K6M0M7hMJMNKIihCmAA70MI0LUvUCWSZhqG
D4cOKGch7Z5kA7N0QhO4f5ia54RK4vLX8XyUgv8cg4sv1v8tKErWJ/RX/eYh4sAbXD4NO54rdU6a
35zHTxKYN39S3pQUHzaLn3W1xMbALob0cdrCi3g0CZFXCtLDGlk6O7vtVbGwBNgtVqnKExkAp5aV
dh30WIked2qjG1OAw8hM4nzbS/U74iseeVosf7xNVUtKn9VtHtdGYCFPSa/99qecpxcjsXQQi/0n
hbbYX+n0T4lQTorUtI+E6V2Yms1TgDmJURBQgGPELsAdJUj7w8w8z2MHut6XCT0NSl9xsIdnmTpP
nDuv/A48ncaOTvaKoh+icwtw2TLbRjb9hUxWtnDH1Xd2M2k6QVqDrllxLfAVIPBEj2v3fZUzi7FB
fCsunKM3QTnYp+Xn5GwAWr7QQNDIz86Dek0ImMyZqxQ1laS5w0V3rqZexS+UJOBTitkCnK/OmitO
+PSJLzuCP8RWaTdHu/0Uo6H/tnK4OhCDfwdyyM3umGhTfrgVLFczr11R4WlYGEBkSHc+12uVGoCt
78XRpuDRXxOldXBANW2fq+KbRrrnei4i6Ja1XHeyR13v2dOIWpxwSNdmvNhvqJDodxriNQ827kQO
2sXcnSvkSAoZyhv28oJOIAJTAPIU2wjTxdJPMOngtNqaCIKK/wl3lkmRPSfHCnFQ5xPVwn0d0C8a
kOsvUCeuQcLMTYK/KTcroq0tRarm0+XJ38SvMrRC1HXnwph9a58/YxVWSJoyVqIFG7VQsOpbqyiB
RGqk0vMzNSGmA9QVoyPWpXRs4viSFsyGJcF1Gv3t3PATruVDMJxBLYfYXTFvqeV7tAqlwnRteHqA
/W5tcAPZ7cpaGftW6cPyQkLxYXv7fHyqAxxpA8XwJSWlA1/2+rEtzNfwYkx8BnHvn96lFEIi4Bks
xWUOk834EPD411iASaDgQ6xWjV782vun/QsGaDuIDn8+oXaVLxSUn4983AJ05U1zfwprNkWCkbUy
LNHSRPtxsyVEzoQSzGu5VienbzwXZ9mwdWxbnQrWkS8/XJ0hnqD8rpILo8Q1/PDmEf9qbbm4MB0u
R1DGUpBQ9zfBNIFsQ4vaxpLMTNqQMIbcayGftauZnsCy+/pckXygf6e9LnezidGNg2wUjBLC+1DA
9cnDG3goQEzBQsdY25CvIv78qxHRfpUnUiReEeTna9fTctRjoPe9vgLMGy42ktpfJMziOlwGGLym
esQu4mRBIkJrOrwTJqeRoW1NS2OEC6bLQ59q8G2/HsDXScBYkpniKHtZd+htDHkBkd37UsjWZiGN
VjUqlY3H1Df3VKgSUffBmhwT+fPX9++jXzKqK3zMkAb4SeUE51JpIxTxiDvjhBEhV/GutQW49jfv
4UZd3hr6Q0gPGxwCyzH/hS+nRi1vgIMawZrhUIHfI6NGPnnt7XuA1b2Sb3/c6uM9S29X2SFceDJc
YC1D+aPWoz8wWCKfltNE8YygSPIBLVQqJkeJpfPgDkVtxyMx404sICzxdsTvDtleYkVSDIJEAbYq
FfisZKuurdPwRByJ54i9kNDQ06HUW3mUTCXfHjj+b2BejvdPjZXt1Y/m6vfT1W5tlVQDR2hJuRMJ
gu2iM6MjcBij8nXkGShNNCZHCXCLfZ3+rLfBH64CqSXAdMpr/WcLuhafU/zJIwy02CQAifQRTE5y
EgwchAAVXs9g++HCzGfzdXEiYAKKoWYYHji5v/JU3VKmaGQGsJYmusHo1DgsJgUr91rVTTzCeXZ8
/tdp2jtxO/yoFVNgNCdE7zMKvvO64SL0iyiySE20GhRi6BTpCNYtlMc1G6yAl70cGXvRImpr/u8N
HO18GldC60w5/S2e9CZvPShvJkUXyUBqTWeK8grpN63DHMOQ/7ZIJWPYsCJKVSp7B3hbP4lHTMNO
IM7s9ZTnPYl5HZck9XV4xg5Rdw9+oaQCCyDb00Hj0wRMIQ42CCfnv1S3hXmcCdlkYiwdmEIqwTkF
EF9ErNXBguY0G5mJesLr5KnBay/MGDkIStpQO/Ds+cgBhNjaD7Tdx+o7emykR4KBlpFVnMyu7eGY
9pYylb56OJrdWPLGgt4z05u0IFcEliKKV/308F1kpyaKo7MYEW7hbDhao0M8Z4j+ZALURSntluIO
9QqutDGJr0qfu8TDqjykq84tV39e4Cjtdz1VJVY5Kioql8OCYQ4XUXz+Re9xevsJPZT9A4ZT+dia
dboslVqunB3ZP6e6DIB4TS9V88PNLHeIpuG8qYSBOcx7xotE/9O55Nl4o0zvbMASdyvxPTubtcWX
ug3JGVJM5sB4AG2TY/E3J8+ueK37jiD6AWhBuND00IP6ygjuNuC1G7fSO5UwKLBrwqJvA/JVt5XI
sTT/SQPYFXP7nD2qQdxjNNdw5vTmKdsE/ojwQdEJk19HOCh1YhSktNy0Eu5xMMyPXnBXOlSxo2GM
Dr7lvcaNY89Wtl0PAfmYeBT/Ljx1/nh5Lak0cAPD07pQzLZW/PYnWCKUyAfOHvFuN99d9u9bHGdr
nr4MJ4ZrW2Pof0fjGSmgOkYzmNenTHj79Qews6fOc9eKsLXP791wKB1nWtGa2N9IhAzUjAj0YLMs
FY7vOWY/DUIocTKkSxl+FtIZhq2pLN9dMmqfytGaCUCrFIGNYF0zp/8xVBS7KpVLRKmby66W0wXF
Dx1apngbozaaNwQxRol43AYnWtOF2U2NhH4YZLOp9cZzHdzGQjTEcG4ZQEIjpq4j3KgKGzU8UxpJ
Pw8b52K0TXKkN/qftX0VjOkyTeTPNEhoLZzNNAZSILUyJwi+aslUfhCJLarYLFcyV8h8In/sCznO
9ZHHDBO6GQDAwPedHwA0yTNlub8n6iU6on2DtXwVQxN0T0drzvId5r3Lu6Ewo0bbfcFvRBdtLee/
fazYTdR7aEzWCE8WQf4HsQsjyoxxIhsYr6AaiEXoAZ27WXeQ0TwYhtRIcYFpIT7hVBbMxqCHbZ0I
y8cP9NNQdWP8EeBhGvIObmF9zIQSjdDjjuBjqfuChE3Anbzh4v2nDFuVV8atV+Q9+D1JtMAmbr1b
ZUP3rNGsNUTCDhul/+9c6oHp7eEwSRGDdo4BwleJ6wNm8kzObPGGRJaH0F+QvOJyHlNNOWv+I+9g
M9kbRFJlhQ2zlngkswdslmAlDh2sKfkRl2mVw6N5KpSwtCX40mU7Tf8jA08Yh8l+9N7PRhgSubK2
gd4wU0Uh1fZQo3Ot/WYUHUAbXj+GvWEz+2lmuibAsxpujc1E3V5B2gvNyVz1AJx/lojN7jSxO33m
uEu/85HXIR4ly86nFFzwgld/qHTXwHrafQ+lhUP3Snbi9ROwZ+Ra8i4+y2xMQIIDBDeFcZloHjl7
me5LtYkOYnZM4v6CNgkfNZ6c8/DtByM7Mq6WbKUYpDUmcxFKgoIL4ME69xU+y8LstU6fTvvzl/tI
VAM4Qr972Lx9WwneeyeOmKg0Jcfzaw5mqV0AwKZjZUXDCGICJBprjhVxdyZn3UUgQwZT9Q68GCoq
na5DwIirg+SU763fWaLp3WCPcAgjw3yeJKVgiml5VxpVBP+Tz5abGt5JrACfuGdBa2qURGF5WhEA
XIqGZWmb8pEclpdVl08mfHg4CABfdb3SOZ0U5cZbTx2KoS2Atz6pWVEICchkUN/DEZf4bvWXFtFJ
bbVWe0L7ej2gmEiHo17hmWeTxQbf2PDlxCLan72nqK8xLctt+YpGic1RD6RJ6prWKZFju8Xlz7H/
RczXGhXQJmYfCdQ57kb60zWbUqdbVRCANbLAJMlDFwu8bJvOfNTE1UiXt/ow6QmvzLz0A4iY2BcX
knNSjCDwIrGIRbQw1W4e06n+ZWUgn3d5SrNSy2VuTr1bEilLATHoNZb4LxB+7z1qcBizNQtODvd2
pNKab9DzzTH25W4Lsva15zIf/v43jvrX9uemh8SELJyoEh84bVAUnShhPoneOH3mKX4d6VBKZ4OV
fCXGzmZIk3dykfUKkE7sH+qeCdsvF8p1qJ8vubblc/w53e5GGfnTUqEE59yujv/6rVO3xFW/vGqX
Alv+frKrHDORFHbCKfNJLU1vN1WXXz0ghu94b1MVgP+nlBfYuBVzvXFOEAofEs2AKHi21iAbyR3X
Okqbovt7tcv1cUhY2GUCkKJKGi3hj5IHA+vz0EBEntgE+azqc6BdFA2WjcKx9F0/zWwfsLqFiglY
qTCuIWKHTqx+1tafG+NjqQ/7z/Uihw6FEOXIq7jnjiE13XxXFhIlymXiRdUByhycM+ERzo0odsy5
MWG0jatKlMTjydQfoW/5TU22yJANJFm1JWdDjsthXicYfE6xR+A3Qx0Tep8ueoKaxHYRAipdsbz4
rWvLSFdPAQn4g8b0+R7Ry59lo/xS98/Jxsosgc2P+6LLhAYNTELprWZ7D58LU7VxPbmFo9Ts/V5H
f61EmLaLHSQwby1KJrcIIQbUVa8kaxobFwmYyUtG9c/UHuMMZQxxAd7FXmeCBrWyHTaNgpXNH4Zm
MVAde9QGZ+isyep15KAREUEI5f1QfS5s27aWCYCBrs2PtyqSQzhJ5c2Iu/7483NpPQAEGpKk15zo
SpW8+nROohTXAxEapvUUEc27hrTwdKAfRqTCBrfHHGJKRI60kssadOdIqSxVB+AgIC53lQJjGYTw
Ol8ARIvM5ih+niDmSJe89fTpWQqvRl9wd0KsAknt5XD1hb9bvdEje1hlKOPNovYw5yl8UcloydKq
PdgufsU68HI0D0+xqpM1Z1IdYcaj2sD3q/hwD4SCRrEKSR/0ujcOtmXQzYyf1ARyQZHB8Qz4DJqR
UY2IajkhngWfV6gGoA1sz964hz/gtBIfzglVfYJWhKPofS7bW3VsLGy+iOur0cfpjjY7FV5/BLpS
L8kASxNz2OI1RH7IE0betqOC7FA0REQbSGJ+XLQuRy+UfUdd3i0bnZnDzRLzQHkDsqX1xcuKDem3
LubQqI1F7XYRBTv3rdzsVHDeQJMH1yABlHeUFAD8j9KKOFUnd9bElQ9O1KZm2ha7sOMPquXf2VmV
JWUpZiu2pf5YqZ7VpVEinlJINDoLg5+NXkPI38sgCHx+roUgumLlyqz3ST9vuxRegDyN+MvTGqyp
B6ZM/gXLiVR1tjLDrMPVo56l4ziz5lWQu3vYmVNLbbHYGirEE3SnQ9sCQiKqwXQxw4Xj0SdmRCS6
vcuRRK2Ubn8dz94UoFnifBq5xmyPGixwnPH0tpV/bf6lFBGOBOWbl943yx57cauyy1mJ+kWYwY2z
NMS5Ah3U+oLb55Ry181lcaUx/S+HaansUMDcAw75+rXQbOhX5oTSNMCvptyPW80BKX/IoL3wsJCC
PL7fPX+CocbvG7oj3YTvxZus4nWavJs8Ti0pMx+ai7tyR8Svl+WiPa3M0TzHSc7+NqEdDq5QhP8C
ZQlRY7CKKgCh3bBaHqSX0oC6+RWmweQNoHhUBzGEgAhAc+3QztZ6sW9NMzBfrfrWiR3GNeZkuUbO
9ds8/WQMz7BHEvB0eiKWz52ofEEyt1O3dvBeePvGt4wwhtjbGmRSYWXWga7weRr/hGFzvuJ9tpkO
gjzS72wQ80xNrZuJVJQU/DHPQ5aVlYJLLbuWdyUTmtf6kZR3q55E+ExzuSDYuV5hxSHLe4kFpTy9
gDOZ2g2iN3SWhsiynl4XDfvqQvWcE5UKwu9oUSz5+NwCGW12s0WeYcK8pgdUQyRc05f2y9EZipSw
nNYtmDSJZMyCDqUuvvKoR1jtimHsu94XAcFNPNxRVsDPP1d9eLu/32ez2zsNnj+keRhzd41FPC//
ot+6z8hc2VpHmuqi/6IDx3ro+9rEDJfFqprPEgq6Yo+NVwJ/27QeUf3SPuX62BBIZvIjyfaLAc/2
ZhG3dD19J9H2t1Pak2Oef6iXLwCja9Z0tywxi6cicL7vJudQCRgq1F58nCPZXDmIN8QPD38PWtiE
Y/DTjNL21JIAQUIkHwq7evZnzPQD3CN9Y9b4Phz/2MQWNsujYRctFVVtU06U+QbaMc9OlU/wqL9S
KWJkajTMKJCLUrbZqE2qCvnX6J7O1WWim1v4W+qusKktX8QegsWBlbEgla5292K3v/F1FDIVwlXg
jfDfVIq+Q/FxIKLiVfaeLcYDpN7QpY5u4UKwqLSIh5wLqCdhwgtZ/Zz2PghVbV+g6m9tCfe5vYVK
Cku4qOSxfFpm4vc+Fs0J+L96rj5jvGnFp2xZu3cOO7pzSVutxxB2gqv74LdwbMiTi5Uz6wAc3XqZ
bXjGng8H5J9s8fRSB5YmQkjbaea9Cbc/Tsu71Q7wjBerjR7GJR1Opxjy/3UESBz+31Ok+kteppyz
HR8bs/Z31Uw5S1hlPzB4sLL6Gu31XeR38gxY0YNwNVfOxeVsDnUZuUYZNakhS4cdA8l2HVf+9/Lv
LKmXLlHT1tO7yD4L/Tobib+HH+W4a3EkWQwC7qHRq10Bmyc1FGvkyF4P9oNeIX3YFX6arFJ2Zmw6
KkNKkJNNvRIsvyoeqFovpUQKJceB0odiZxSfXf5E5nMXQDFgWIm9k0uEQn4fh2VnNvej/5KTMwqt
tY0j3YTVUurGTuF6mKacBL37TbyS4S/iCMfU2xqzb5KUbG5nl0JfEMugvyTK4K+sIV9lxR3aP48a
567RB8AWjmPc7Zk66IltaPJt826HGVG2pAe6RoMvjubp/iCdUGLXoIwmY9UgYKnWsi8nC9bBJkQG
8gIgWNYhkkxGKbDuQNTrFe7OGHkry1/NdW+gwkgvLtaioP3TX07N+WXdMbu612lRaPD2l8p+XmI/
xGumHGaj0fk16HCjPfbI3HbGwFij/Jb9y9jf8ScSaZW/Moi3CbhcIRn0jkocEesPsly1U7BRjML1
rC6ZWH5HXaVDGtGEe34eFRDvHE4bMwUEFp9A76PGzwwFyqXd3DpzXxGeehMh1rn4KB1N3FBxpz4L
Vhd4ZdwLI0fNz+Hy5c4uieQfrfaZNawwUzaW1CLdgdihLBIDOSxvc/N4OSsN536kVBoiEUWrtuIk
L3cyBmyRtfoGRnMFC/ScDhUMEht+kTHS3lMk8U0RP03ravnEPTqD8gS1mZRvhcWeSfRqBpw6KceY
vh1Xf69IY+yCtwtGtqTW9Wwtm0fGDzzKb6aW/BgGz9lxYPrkZZ/wXoiLV9+XsbQTe7q6jKxtqoFL
kpBTT7u05F3vPBch3gCPZlE3ta1hGYPXLiJiFKeYQisRcgkujhPKy8gs4AhnS2UQD9eqeqjKVFQ+
BefGKakr5ND1f30EW+pYtBP2GvNsgNrZbmD6q/ysh5xFXLX3HG0BCIZ1JLSW2hDHz9kQGBmkvWa1
UU2OYRslAuHEwupcxn9DUcMFgbWGQT6cvho6u71HiZea6bqipRLlMiljKKoyU62ETsVk25zoXXKH
omVS/MOO0xCycRUWHa3pwxTN+L5/CF88yEJglhdaJbzKF7YmNJ15SrqI3eXopMxWoAq+sRGO/lnz
hN/kHWzlXAVLgFXZINy4hLfXOdzb4lrqbkc1wMKMMs8/WddrPxwO7sb1Se6KTEpCcw4Mt2O5j69N
JWKqmUhBSEzI8WrqrMWwocvgn6f8qWnAy15u7E2s8MMeDp1BxiGwQ9MT1NgJ4vjz7UGfskxN/CQ3
WgawnhzGCAeLFDFYVSP28N3f3/2lBwD7p6HSZWyOuVg4jeufcdJo4wmgT437xRP0zC301ey4nR8L
o4NKZ61r8/1PLz8TdWcmwgfjl2SvgdsceF1+wRE39AaXjjxn9OfA6+Sl8HDJMetIv6oKqlAZ9KTV
oRVxhxVypBVcnGNyVhMnaTWQma4SWDLB1KXTdm5cTZueZqLrJGoHF1SRfm8ZTg783dx+kD1q9zlk
wrs2q5sUg03sSevKESdrW0w4EVUrwEbFSn869Em/cGrKTmwqlW7eEsPAEDc6Vd9Ju+6eAJ2HAhH8
1EdhFNvuxULpM9bIOvuQziddIf7bMiuQ4fnW1V3XJqXAJfufhxQesxBo86j2o3lyQkGnAH+dHQAz
4MdS0xRH9ayypku9Wp8++G+FxIlSHJNMR2QXrIkslJm5x2z2bJenMzMer5YKBglwizkKDfWTgHp5
aB1uyqze0JMAPMjYggjEAaxZ+tSeEyl8e2kE50nXuFhI7efCM6HLPCOn44HWeCPXHZFD6H4DW178
tEwdhCvKx6DDSmmu2boxg677/9ySXpuxxD2oHzorwu3CMq5CzVz581+yheIWE+GudvmGr1wSLxLB
t8oHqMpVmrIs/oCv58E7hPUYn3e6anEvyf5uKIKpLoAj6rllo1XkRu468EVUQQRvtCWsW1tb38nK
vLrhNw2QwdUsbxYF0TbwBNKMOiCjOeI/UXqvBuwB9irm9l7/DsSN41r9/96VlWZAm8PItlV2Desa
j2R+S7TfldReHtmf3fovfqiBFbjl2/VZOzFiWQxRle+kKyYCBKpPz4h5ZGbG2fImMv4+jFykMXSM
uFCBMXbiJ4kIftMcRO8sL+POd/27nJDoyyqX/kNCmjudmMXN1Ewld1exGxlcAvvknfTtsziX85nV
NfTZRDTrnGMPwn/YFAQow78tM92uV7mD4TZlx1GObjXGOSUkL1XKGjTd3aq6WUkB13CTryD54B0r
ONUMN+cPEpFaxhy8Vv4VyRPnqK+pCuOUWmxZv0CR3TVjW+FPyPnssyrFYWs1W+bd+qhl3x8xsx/k
yoiTihD591WC6nQwp2yRW2zmMoOPrpJb3/Babr2t8hc5uv/Slnmqm5bjjBCGGiMf7Rmwsm0gvvai
vQqVut7JAV2R8RirIGrAZfpyddMZL522tlnT+AWspok7SGDMx41rUrMBL5rT78rblVs84JixXsaY
a8/BpON763aYlM9LCLKxxdHlQXP5pZaU7/pNS3aXRbI4ePoEoH0VhSf8tkP2l1KmsSCXgZku0cEA
c/D7nm6DuL7hK6iMmvt1Qus6Z3oOR2533xOdz0j/vQeG4w8i9cHzJxWkvl9GFQzZOFcP+rh1nQ7b
1gacdkuHIKaQSsmNdBEHMf0gui2PEjjxVWUN90/j2W5LqerH988wLvAWguoQJ0PU0xARsf8ZH4Nu
70oYqH6iN2uyXLWEamMWtqopnzMaWIrqLp3Sl1dynesOc3EAOFNNPLCKebuqRFAT+L7GPmxM22bD
EUj2Llrrweo3RzlIjxAhoX2HJOWiEiHsuTehsoz5uEwYyFiZ03+s65fxNBc4La+RhcXb1V6h0sxq
dQq2hJNR3n105SRbr/1bEmGRkHfwgg0EppFlMsz8EV6Ezsrl0oZ92p8Hyup4e3169UPGx4+ZJlyu
1csz1546TD/VmgTAtPXizfeHXRKVJ24irw0LROUDG840x6ttYeqH36SUZqlEBSqGb6HxI83ClzUg
8fLueo63xrCc8jkYEqlx7wExXbpZzkbDL9ogOVpPUlLyDCqtOuAiwr3bZ2CLh4x1x7TZj25E4Tfm
OicveDyREH6LlsBNRLu7DgDsya6CaoslKD/Wj1gbSm02Cp40kgkTouqX4EJNDnGEVzD2J+dwePUt
sVP0hZQlF21VolaBvDJ5SFLapYnGCDumAmk2RFohDCq254Iz6Ap5+3K0jA60la1MQ1ULDGqsRqrC
fgylph9kUE4ukWE2eY454/FYOfUEYIUcHngtjOfH35DTeHE0JnjJXCO+uuKe7oiEN/qmIijiYnUt
o/LhFmf3JFZCtCxN+ZmI/igLXQJTCrHDllKs6cnL2+2t2ruDhghZrvHSq9L6kK2sYhjn0zxI8wb7
g/lEjtowA8P/UZ+w+E4m6BDhMMrtLry2q5aF8TNaV+d78q2EJsSyJsYclQXY/K8gEpkrNkvAqc/i
C2FtkiPFKBsdcj6cr2mtrK07hG27ZYbjFM84QASIJlV4lJkyDv7ujRVZ4UQ2J09A4elsGEhn8m+s
Jiqsp+01z3K6akXdv62Z+B3kH4pXxv6WaBopPoGKOHOksLBVvDNJXSa9/rFqnZEE6LNUx8rLx1+6
WJQRFC8r0Yq+94hvI2t92t+bbDsJR4wl0SQ1nOP3UYzqp4HQtzKE5Z+4XIWJfUt5XG7JwY04Upqf
5lvZ7G9SlRzGhesAncfKUaaD20Dr+bsLjaoJDVIGYMAm8uU7ghcezuj8frGQ7PcSo2sP2SAPbN2n
pFaNNJmDSYMI9Ho6y7JnYAK31MLKFK/DIhGlNr5KAt7PV7402Gi2SO8BdHkQwerlEVv/1kyncOPH
b8GS8aZ5LXe1WXU7RTlyMlr21RajQmngoYTTb34a4OX+08lHx7FtToi9rRb9pCLBzF/N1fl717Nl
nGWx+Mf6ky+y7E4esYUyqBvRlzkdW4cieuNLg22a72eJ8PmtKUCVMnjzc0rBwY94ORC/JPOnAJoh
/WfID6Z4Yb1/BnjD84QrH8ABAkC1zkxRdM9WSHoqxB4XOTVI+88vOVi+CLaQVCT7NutF9SyvrtBF
eJ3wTvjdYupmsHS6sV3+WmV3Hk3KDu1n5qa8rc+ZtOS6agkuJGZYcuqRuHIp6GMTVyi11ZV6dIJv
xHykltvZ+c/F06Xrp/pPAQuGsY7nBznnSGLKDwYAP9PnU13S/XgyHJ23qhJLL5e0km8fva8r9n6S
7HvSYmg3Ga6o1PDA37HTAtBFlqOQG+2SbyH64jDcB8Cn+qpCxIWS20tgrgvach+eU5+LKQHcQLAI
HWkRm76SXxo/3X0qyTvpnYT8bTpHliC2HqfkdCLLSYbdELRHUyQYfYJMYwxGdBfJv92/fVn/KdKp
D9D96v79rQDnf6QvEvRenYJzEQ/OXOXYCpUEJJRuyQIMRMJU1Sul1Zq04klS7V/ERoPKHS6YiNwv
YYL1HlP6iRyiPW0I0aPPvNl3rxv8B6dE/JqDMbHi1g3mka7fOibaC+EIXAFF1Euzcpk1ahbc6wFI
MHMzhKqX3kCvX46xRBbvDzef8F46aFfcpeW1P0IPTToHu4iXUArtrS3jeHUub3Ht6UaFfYFfmYRo
AvOKe5CGNwYFOP1gT2g/7eALG2OvChk7WMiZ6Ux3b7luMXVNcZFpEyOsIXvGE/g86UxUQBg+kQAO
PN6BL4xfYDt9UPEAIou+SWBF3TR4ZH+of81DYoLod2ATz+aTRESLjrwnFki4pmtwXgw9sXK48MQu
Qyuo6C9QAcjhhRUy/wOrB7d1Ghl9eJR4xlXeJmdhWzAVuTdZYfZIjENmLGp59bIHnPUXFanSR4Nn
bOx/vQ6cPg1T9TcygVHzDJNggzI7Gavt+DIZ0NpgAahqWxrGudQyi6JRwZQwDlMMADjqdlrmZn+6
6cfeU6BWuj0D792vOVsTT0/KcwKlPJUkmH9FIb6b3171jNgwBX7ZzIGvlgohWX3LnOAWS0CsbufJ
QtznaSvJXbS4Jj5fHq1CKumWQ+4WEClH7OPiwLWt9dVVgbciJjOcN1GW87a6/K1MGeYAV7TmDQz2
S5iZ/PsIqfI9/GAaluFfTTi8Pgy5F9oONORYoh240xnlSxp5B7IWNmSY2E8KEF83JXKPO2UZEi/A
yxvBWs4IbR2dS4OmAK+e2zm+s833zNkhH3NMwO+ehRDeoWHEQnUlMcmPNawnhf7awkEGwZlVpPO+
7q29h0GHXtdWukHuwTcUDZxv13FwbcouM9P1pKRE8xwVsPm/PqOueHVQpN7/USZAWhfRDe82Z7BA
hbNFR1S5u8oi4oZ3DXy2Swaa4RBoDHCxveZ6z0kxMx+Zv89dde/Zbk5SiOP266aH0QHEsWxR7MrO
NLo5Lry9skehE3Xl1AM+STjkYhHdanxkKPJYWTn5GY6XbJEcHRiAQHZNUOS1DOai1mM5B7Ppdr90
Y/aB4Q+vK7W5cWZMvv4cxAi20d1KD8uAqfr1OBO0ju3GltmimVjX6TtG15L8A38hkMyH+z3/Uasq
kfHgydAaSfHRSZ8j4HOKj5Np8SN9H40S21pIsfYWjJkAGvOOrLwwOk5oD5pEPza1VHFLIDy35sTF
PatzOmCqAe1k/WPQUMrHz10Ul7h4CTGB/gds4gcFsKbTlXPxjubg1nuQxp/+gImgVlV9bRNS4T3e
/jCWBCM65NQFv5wsHIjtiGPQRFp5F7XOV8aJnpFYi5IftZyWC66G40mo3+nP35R2YOeX5kKlU3AM
J5NhgTUKrqUDP7By7wlzXlkBdLicbC8pkKZ8C/JkRGoYqkYxU1FGAZdYKeH/4a+Z+omL/r7k7Oko
2/Bt4o73vCvUJVXiyUK0ndU9SpU7hrc/VYsXRrb5WedHl+81uWPGAD+k0UjJaLBVcdXxMlIbU3GQ
XZ7dekYLLSTRAG/83IXOllN+pn/V3T2fQuRftgDtwcaYfF5/2PBhNzfDk/jUSjhZaFnByyedvMtM
oU236+dXqsUFfpQtdOwxdRY35tHPCVBuVe82kpXXf/ZaoZJhjDCN5uGmMndigrrWQVGlBPScIY3d
2QOTH16mktjeSgBLGwQs8WtcI6DvpPN+PgP0BPPNh6XvsgMsHYhg1QxCAdS8afiBFVviuHr8TEb0
RRmQedegne+p6uDRUqSpUzLVnkx6RUXbivBfIdBeYjXhor4hBmaeC6QbGFDygQy3d8+PGQE4P+Yq
HhsM8YCLKR355/9UsUGt/R0wfT/5g7jF8WoykrUNzRvbPJ4ysNbqxeTPSHTYb1WMDtegKarzzNou
YQAnTq2vQF4z1mCYk36Uw3sYLmT8hk49gNdiEWoQ28p6WrEXo28D/L0lsxuBgspB9FGd+lLxejkg
ZwCDo2KZ1uoxkCHmsjjMMm4ct0cOueG4Aaq4FCGpu928+YPuk4a0g4fN56EHlszsQJ60XI5m7biX
afxmvdhUolbG3hsxUgdXA4ePZmwjvX6NMz0QbutUDyIs0QUB0Sc2YsCIUhl3wJVcLJXVEwt6MavY
3hK3m/HNCJJ2mBEJ+NTM/RZ5RSzK4iTVzr8/QPfLbiL9iF2wUQ4P/Fh7rYhWg6v7bt5K0+Wh8J9i
SNWlMzaXbQ7BGQ//9ekj8qqCXTOSR90fza0/AyNm0+xhbTojLbTYMGRnYr4QGlFEP3GfuLFSdv9n
5brIkpE6h/WBszAIBAMzWModTE+P4KrnRp/YpxXvUOVmbOXSKIFk6SBWUodUrKkIYqCXG9SlVCSP
RLa0GMlWDzU5F4E9xkSlVbr3m29OBV+kx6f/FMU8+u9pz1Y3M59rAaAgyohZPqPBTYw6Ogw8QQQl
ohxNDvbMAHt9w5EGbyc4xZ/lZXq1uW08B+pKbPP4uW3XVgUaAKNkVLCKMG5Jxk0i/1HcPrUVIZ1C
IVI6VPYq+pIvrx0ut6tBp90IYMojBcIHwexFcPhIWYLGNUVzlkzrEVPnTuUuf1/EbFBvHTseEpzX
W1XKnx+hYjIzNpqGzQ3AvdMiPtD2aiieuGaJuXUnAChkuPr5MISwr6HfthWqBUqbWZhNF3qa/3Q/
XIPfBmFV+a6zHdmWYDP/w1qPEGPwwqQfn9RbXYete67q3YFa6gVFhv8JgqHmU5PQe5NizkApchne
zGqjapah0Y10Gj7SZ+rL3tDBuQG/5P007C5Irz/RznvDOWVcEe3cgD4j3MiK+qBTgcjBaveEqiH2
gMN5If1Se5z76EnpaPGLrkrszd4eqEPW/YjnrBdW+55XlW45vmIiWrUHsdeLWAc/aKLU5Ma9D6+n
3+UldRAGOCqAEfo8xFz1hpcAa+fgdd5x7cVw8sbc9aZ0Bb3eyriQoS9eRcvUkGxjEj66gNc7Vl0d
5esgLnbEkj01AnPgDWgloat4yFbFfftHsKXed+4fEatP8BLBgH2gWpvgyzPz3M5vhfDRqUNHtehP
BeZB3ZZLDLQDQZVgNO3gCEVRfxWtaKM8vaUY6MOUDISDdG2KCFC3a5j9Hj7Q2lyDksBXCSvEntIi
9lF54slda85ehFYeicOgYAI4TJYkUGlRvBT59TF284VmE1MZpCtT/wV2HsML7fx08/mEiL/zahBI
Wse4OM35bFgULH8nSZKSjx6uNCktiB16bFUVUOTYWIwhh9G4gEUw4z09LY7PnchzRpkyp76qJ/Ds
RTiR6I7UlDSuMOgfk3DUcWRNSi56xK2OJj5Ve/Y/GPeeIExnPar8RW+3lgu7EC8DNofiwQdQotVw
ajrPU7ZOewbiHJZi8cr/nPImXL6cvbJymisIG4R2t2E8kLP4pSyRLSsRVnmS3HBO70Ycr3HGUnTP
DNODKoZqlbOHCi8VVMBMRKjMeHQdvIWn0+rjzyvPSkuXzcp1NcxKtrP5cmxK5hzLu7QgK/kA0Mdx
has/u4SwmDk7yHuXumluuIZ1YT4JVHZDLlut2qyaXmuZDOuyoesXfo1vcPvhEvep2oq6osyyKHzJ
7RitG9J7JBIycJDpGRYONS8oIDQ0yQUy6PY2+It9NNVdwcQM2OX/kuszVWf+lnere2mDyYCc9dYF
mUxpxaCVIhWUjPYkFz3CaM9K23dcl5Z+lY4yI2epgzKot8Ujy+6Qa0mYBLf6wiSZMaAOKO6r3bQj
yTa7/ELf3oI0ny4QY27PUeN1nNOoiG6WEHbG7WZpJlPVHkp2SDCkgIRQVIFbW3klDqegG4JK72Kn
4l3HVLL30bmWNP2Sd2qv7GSJBkV4jZmg2Zw6HAmbhsJaQOm7qbErJs3WaXW6ZEO/3EQ6+SxIKj+K
M9/ySY5m1LgVu7fRRUvNCjrhY87ASvumNIFdXDxvRjBiG+zeQrv2nfk0YwtX8FsI6irJhs9NBDI3
B+tbHe9p1z1pg9AcncNZxmdRYsEi61ZRM15kyp26NjKrmxxi0ejbzu1/tDly7VDDXfoLBqXE1nGo
oatE1tlrry6+XruXJF89fZvBLTCNOBCt1Sc9ue72HLGCg3J4HJVSL4/qV0tbedrbyRdSNu6+9Hwx
rN+ocDRwukC8Mru8N8uIZlHnxGxLtKMxnS4LLbbNVRlYscgYgfn2utaXEoY/G6vuNGt1mWe0OUXp
oyfK8sC/2LGk6dwf0F0NWYDGns2i7rz/KtTd6IpzLr9jTIHqCcAQox9cng7xZ++I1Q/PsyR+ctNI
R7pXsOJeLCrzSAGNku87LZKvkibMeiIBz7OZZEVtFnMHwevb+8l2Ntw4bOKCNYkMNIzWOvmPjRhp
gbEt1ji7Uv4FjHtaCAO/WVF2GOHpNA9nspES9tKXtXufvMAsxsY7r7n7VQBDH4RqW+IKRSTGP55K
BO6F/7fwd+UPFEURxP5cSG38uEmRgC6M8jqnIxoeR9VnZKzIwwCmGhkFfGex6mP8grFpW4IXPB1u
aejvnm53avSwlrvWPX4j9Ig5aHvb0je5z27aDUtuX21v+UT8o9Lbwo5zljCgPLdLqOgEomIa2J3G
kimxOi0/5Olk0CStLn/V7ISRr6TcDFDvpgx3BiUVL/LxRlwsup4ppVmXGtHk8XxVH3xenqVXg8F4
YpHHza4VWNF9LI9F07W8AHSUMUsUXmORwDa5VT2xfBtC5v4zDzYZJn4GD9EghX7kQKyF05aiJBpC
9sd5qKac8+BgGOUwUiyKcTgetozsAxchGdF4JAsJVsEgtOI4Zai0HvChom7lz7gqzNv7p2Memawq
ZGIBcsRHuH+A9Gmz8m9QPQaNZmSO1+mJCZOdSX7G06/aynNBvuypaiLCUdrmYtN2t3m5ys5AMJLN
oSpZZzuydSIxetmLNDgH8ewbHmDdfFwMXN10qlyApc+aSmhHR/flgm7xy5POGFQMT+g0aDSaTqWg
w8u+5EjOyG7b3LCRjQTlqyxhnUh2g/MhdACxbGEh2J1n8VUn6GpTcOQF21D1JgkI7707IBww1+cx
owSorMAnFS9AIv2hf2uXJq9x4vKib0NcEBgPQRKfdGVpe/bUnkwfYrypKTQ/QRkmiN9EJGO+EmR9
VPDXfjeoRDLDX+IWf9jVqDK6o1x5MItV8ncd9+GrN5/7lw9u0LhunKWIEEBlSOxxFvG2S9YQI6Ym
JX+dm2mO3X+Zbu9QzPprPdMz75/13OZ5zBo3DfQRDR+nLJiaqDFVLvH8FR6Ter4rgm50TfxLd3i1
d+zF6uFJbZZY5VpyDdguGpPpc7Eq51IXVcEScva8e3/C2NLwikiYpT+V2gVSeoPUCilrWIieWfeF
dlBusUk3EGvMjo2Rfd590AmbDGWexcUdqc5CcXZ7n5F18/4KeoQ+H8txw0plOeoafdyI60FWDCZ9
xyFxI9fZJgPFrflBT2TFlom5KNacleXrq6xvqpRG21XsTUfbZGhkQHSHTWem7muwOB35HlijVbaL
UsOEnpYrw5XDITjLh4oqeKRcen7oL2HSO3UREvXPGUetH2+TqhVMZ/OR5r1JOSLxHT2i0+/Zz5BC
G/K7k3THWtjHiuIW4i4GTaEJo0RzKxV6wdAccrGUS2ZditWUOW6IGizY+PhhONSJHphit1t7iD39
7LsWidVRagYY09Tf6kBiO/TpOgCBVr3q2zj7gpXFCjQFpUeO+geuLjrHBOK9qoCunZuqyDwyr2cQ
nUKkxG3Px4m9lUgFqXXR4yMcer4K3dIrLJldqmDyKYg71NsmdmFwQgvsifA8ZX+sk1sqCAVHmesj
qMpC/dZ3QbcA1UKxe5yo14nltra8deDiyr4DdKldCRZ5frzib9E82gHyspIoq+r9kvTZ2l8OqFk3
hKoVtYzdU7sMHBAiPcPLaXQ8QVORG/RXWggIkYZCe9XYCnJ3aBdB8ELkSqXRGuDJ5Y6pkHYjyVSm
lJ8eS/A5QrNbxah+rU5mIrUSxfCt0gBUFtk3rf4EzQ6Gpdcdh7QfYeMw1qLIuEDik2Hw/d3SvSBq
q7itLLO+f9WdxQvdXBdSn294haPRCVuwZol/d1BRq1jbtE9AvjUSFlp2H4eEq2zai4ZgS+Rwcwdi
oYUVazSmmEokjGyH7Wm44nTeTsEAA+0no7kXVgwdoK/AGP5kRxqhuw==
`protect end_protected

