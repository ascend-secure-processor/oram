

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gn4UDFBHe9m14STdgPjgnK1QV9pDhJaahbhFQJjSM4TnUP2HsnAmFCMvfE4z7Ie5+t4JS+ILPULr
Nbxy8y+PvQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
km043l1n+oYpPWA7tEivfb3CqLKhwRNSugzWceA8XOStjlKHOD+oReVJjB/CKL3vxfSZfEsx8Zm/
Z4XUnjxMlANax/2VPnmlt0BEyAPz1i6Rdg2tYbzatdzGskFBq+5QsSz+77c0oGHb/L6mDw7ar5g3
BfsYSpWEseEpgCyHMtU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W/7xlCbNk9yhiAuzUi4tlL9h4dkIGgBUzHonnZ75I5A/CF9E8fpBxhynFkekzWjnJhwUzoSDu21m
7dd7gNvWqWQ8/1gK4gMWB6qT2FtnO6vdFfW40rodimPdN8NzV0Ky2gM3KdjhbXLtQzGzrQET4VOI
CSkBNcCLnrN4LYpNfu8VCyPcv8zq0irmz+xX31AS+QGFVigl88I5StPLw5M27pzcWljs40A36Jfm
FB4VT1kEAZJzudhGOG7bnnXG7MRxdnQjipWipCb6qt2kKp+DE7cUKFAVVcpaxgrs9l5m/cFf+6pV
gQPg40q0XLVO9vqOFwn/l48zinneUbiZsdYtfg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DfAUcVfMxGR0rjYk9lhHawPNA8qHNQXYhkIdCdV6ybXqhh7MDLkTcHMlWvFxAgi3KnOyxJU/nGqC
w+lRbtSXyhDJcsl+0wsIpSrO7u53XczEsrgcoxoXDbR2tK1LZzbY0gqgWVndmdVTxxpgXqtZYvFB
pwBZeNrvlImrl9fS4kM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JxAbqJVcJZcDYaEEuVQUPIVBAunpw9UfOIZ7aIYuGml8NZ/mNUvjerWZ4yQsa7j0XEteeArLNH9H
nnWWs+l41p5sQ526D5G5uX9OpT8A3FIIJE84qXjK/vq9aCwTHugN/GhawvPt3kesvJHJaMvyU4dR
v5O3kNUijhQM3vG2wBVq0RSkD7m96rP+rDUyWqtAzN1evf3ksciYmcO4+LCXiXKixvcQSmt7rke3
UDcq7HedajqzH+3jFfcAzrlAnGjhj5I9LVaCrNwGBltcD5vMKuOKFDBYpK+2SmwHBl2FdHC/vNEy
l+TDLJ+tesdcf9ccgXwMyMMg0mLedRBLgYXygQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 144176)
`protect data_block
5X+O45+GWYB09Du61faukiRYAod/5J/7eVhnqWQ9XkwbQ/ZRJw+u2K5eJ3Y8jLGf971s0fAPFwmi
XfL5sVkBP2HL6nF1qKsSo1ZEf+Cn9rX4mb+UoHc4i/AvyJQsBSEom319M4QdZQBb91s8eNhAakgC
xFkGeK8weFRnHJT1dM7t7kncNJrkda6M+dKC0478rYxiEiMY6Y9O1gwJopp02yBbO1e/ZzUc028Z
2knWFh89+IZg62H0/K3uMQ1J+/E7NQoeTihTAu29uWPv5S/Vv+MUWitXoKvqfSw52G8LlmxYyvv4
8xYBVJ6sjnLJHMKUF6ylxb8hQvT3cZKD6EIEOoq9sjWyK1lETu+4opPQO0UWrhrL048ccPo7Kc/p
WAM81c1ItY7qytPysezuOTfZs/I4YLTbX4VkdHOj4UP1Z75oqI3ctePXjrdCs7jvE8yCCCJ1Utqz
n+jO/79QmlQZvoj5Ib848SaSZ/Urq1RQVRPrf61v4oaQzG1OvoeGRNwUs9GaMC6KfeOZw7S8L8Og
ECS4JX96lx4h6Qx6mZQRIwVTbIAbSP+MHw+TpZH4RFpqvoZF0LxNayja/a4ZEJwcauI9govfK5Te
H+eJgwESreffG69xuOlkD/xh8aXYgmFOMr5FSo58Le4EK5KkibwKwAYKIWNJ9HGR14UE4cx/kzbg
kU5iPpSzUBC2OqR+AkSi8nl6Br5dha70KLwHx5I3xj6at0Flh2ompBRY2qzugy5K+f7BEp+8nNO+
jDPyWTHzXsv+Y+SBGe6waat82LaojPdo13lqGFdrORAUnJByXu6ZeY72dQvI1M3mjFQRItCgJ1xl
NG+AgsQwdhK4ndCd56zaM/dL8HDJFUQHkHlVt7sUa640/DhsVvqiPZaSI0TTLNe8hsFUfpykDqpy
CgAl5HvD+jOlq1PEOfgXZb4EwuCuV/9z4+K8+W8KkMF727I/tqozPasEE4B69f9SsICP1jmn4/vr
HoCEmn64xyzgnP+6u95BvGoCNVzLyHMpE63rUlE6Jb1sdpGSBdZkFvw69S2ND5tNl6XPr4svQJzl
fTCAI8SPLljxR6TsrW9Qtp6NcJQbOx782KudUHXzDY1h5TfWQ0b2pFiTw9Skph6KKjM2rcrr4esq
K9Ga8zDDIGvkItVJ8U8Won17xk+HKD/EEyOnUG9q1FzKxDAGRYpX2t6YAl8a6byz/6frlA+Yp0ZY
iANMQhJDZqLsPZoTXeT20Fj4A8IBahqiemQDrzqTziOTSL5qo9ks9M5uhw7tKhQ0UiT5JAsg03KD
Fpi0CTBbIJmnbE25cvhi+kXoF4oWf2/xt9OPiKfc4UTYMTOei0y8W9njK3KW/9YDEfD1RjsVZuQ7
LIHmj1TqwU6twPSSO564WHhwdrAeeZ7oozPh4NMyggBEralB1faK+b1deQF+5bvA91RTDS3YNsn0
6AYvwksC39Cn2upLmgJ7k6MxS+VNk0ODwWhYyxU0DhMuaB5I8eEuS5ALQk/frw9Q4uYz597/v4Ek
mT4yO2WaSq3X+dGvqZCd+r+0EE9BOk8exfjzZEn8nKTjO9B7cx1WaJY445IFQZYJYUANF01yLQfJ
W7et+/6bWWswftMsznoB/ECpTMKyTCRC6O6ZfgSCpJyb53SseBtRDphj4MEV7saYhsp8tXhOIxpo
Idui6NmB0mCbXndwQM2dGT6Q20WThRJnijYhoOAxF0YcDsIbqwlLeccMPt2Ci2tOSHB7RciUy35A
zO3SxggLt/rPzK0fg/YLIxuUqcC4/jMvxBXOvTZQ7rO+DbDmE/1szQ4aPRWl+Q8A6f4/hbuBiOfm
mbCjnGQcFujOBKprqxRYoOOLoVx5DXrNvw91sAKDEGZZx9aRmVzjz3gjDtIIAVPaDI+lk3G9VC0N
XWxtDyVZZ+jl5q6hUvkOGt4OtH5lqC5NJ5R9biDT4wmsUiMgG20J7z/Z17a14EW471CDBZM7kaO9
ODFzgNc5w0Q2PfzzoIMxxzb3cb2qf7V4gSMHDIMzjFroCE+DGLmbAg7PnHBYyPj+kGaLHiJNcP8c
8/jOg4VV+S7LjZQTlL1w2qQEgWM2G3c5Usmg7jQ7VbB66Hk0zzTUBuTCMWTD9fS9fwNu4lT9HdK6
hEazw3bLIwuIMS58djZgpsVtamz71zDYT+OURRmnuu9pv5HZSr504gR4GoZKIezWW7KNOp9ZokJw
OQp1fTS9hBSfQkv33L3s69g7hQVRD2rfWPsfE1R2hlyaRGg5Mt6ZK8H65ZsxyYIIxqeMJj8xVUWQ
A2h+Ya2TxNP4cJKtX7mp2c105NxRnjbmH10oNtUb3x1bifKbOWMnNptuVJzstBge0twwB5+jNxis
0C/anAu2hEdfBq5wSBrSg1RXnZTNMCqk3WmQVRAKzWFMek1SwA3GnXGWAsqZma/4mDjt6XnSdP3T
Zy2KBfDeFXu2Fprb/4SXimkGEVOQnUKEHB7M+uq+lISoNmptGl7LsiVxB9hDElS3I63PWCvXRaG9
9pTMdMsrLaGyOsocz89/s4WXkFX2PIUvROj7Rop66xNVyUN8vMkuatl1yTM+tG4XO6NHtN/y75Qd
uHomKVIFNyAUIurvgUq0X2jKRPfNTrbqi3C27fv+TRS6yaV/XFbrxOkXgKOFR2ATMnp2Havjcz0E
nh9wnFoC69dx9FkGaDtDNw6NzNUBiKTYQ/Ga63ibRPTzTFXCbg8NWzrVdNamePBy8MJpl3ZG5DwT
txQy2RAaBK78gfcjD2EQ6LoN0C9i/KaZ6B7biMhp4QcxtTJPUAxH7z2bbyF4derTXae+Amvx16hA
A4Etl9TRmBApPnch7MwoNBXLmHM8S9iEc7e81HOK3kRQodgaYoA9HiLLZ5mMO+3QqmLwaTJUYeb5
L9CX1SIQBdy63HeLW50R6hUIOXYQtHXiTpciDEzU5GhM3JOY0VJduEHpJ02WapbmPTTJ/hMzcLKc
+AYNlPD16b/X7KQzytFjAG1mrPAZNW/KMaO4RJfd83MIrnzbjidYrpUPDm1O5BBe8+i0+rZphDWl
jbYFuTRab6dla1ayxSJBzWVqt7+N6Tj/Epj5FCUxYOtVrCuomf76GhQx8+ozHVch3RUIpGHVhkys
Gr16IjsXCSQzsA6ZyeIBOttc/reG4q/qe63tS6XOlQgmhx5ujau1+I7v2a/Sj0sfMjVg8zb6/mQl
+Y64LitBcNlkGllW0Ffw95OQOS/8DZDgz7OlgPD5xV1tpBPFs9tltPaL6XHaaHyyN93SK73vth1I
IVIDVkw1T3DN/tWmkUsXisRKhXDJ5+YV0RZnNwLn7B3xbqr/H9+O5MpuWefu+Sf9T1cWqX2H6XWb
2mDeVsA5jPJl3u/NnI+LCV/xEGyXQRAlUifg6voAUhg0G49fqqNRzxBw2nirYT4TyxiDjDCTSC2a
4wuROiKlQAWim8mxTJsrrH5dhVVu3auVEdVHM409DuCR/r1dKjLunFP8lSLHixZlDEaqciTCE5UU
TrbA6dysYmZ/0FnFUSIpE35NCKt/32ZakkepoGnqgszzCEEiU6u5KDHOvi10Q6WIZYPWsDtcx67f
VOSayO0V62nctweOTue3N7LgDLTqiuc8yFgBr4osYoJDQA4bfeOjIiB8Kv8PwA7djwT8CCVgbZTp
sg2KTBH0cLN4Te2ord3OwTrQ3QDKbfc2VWrN8Cdkpr1zxcNbSUGGg96r4ADjzP0UaMFUsUpsh1hQ
GgvGTWh7XgOpN2p+ZQyMeoelhMOtldAYtGMFf4lIu5qq+jMkefJNCXsTX2KZnD+T43vJkp7RSCB6
sO0GAxe7OZs2Nm3FXr3cYKgl9KNsGKjPO8mjHnYXVmrBM9rfY0kNTgoLnegk9XgkgeM8m9PSsMkM
oeyr+/hbPRBTvIc+gHLx1Y2p8WJebLgQGBjqZgSP+Uu7jtcMv5Tbm6gSD//+gKuqSiMNBKUrz2rT
DfXQ42ZVreZYDER2fj6UX4OeEZVDg1pNhh/8ZHWBxlnhjgd5LK/FigS1BMiWB2zx4KZGEay7v/tu
vlQ0yv2EqJMFRtOl/6QUJVuJAvpMXVXjxpS+Ze2Z5QuaNuPefasIoHksStucNPl1r7DEmM8WUvZZ
2vaRn3TwWcDf74aKzZaM+jKkLdm5suyPiRNs/Shyd3iLBErGyWmAsaYF6BNKk7Otl6GdMV1adrlw
O441/TlWNaNupMvd02wSFvlGDKJSjHqx/qflLHEIFDBrEAvsj0q9mZ2apSx04SOXPe5mh4C/bx6f
qmJSchQMRbOvVVPQpks023wVJPr9NcqG5R20ThCuAxa2QJNAmggKoHLSs6oFLQ3umy2NL/GmbmnW
2dZ1qkMuRe/Wu2AwM3V/pQ3P5ixI0xKPr47aU7NT1jFOZNO5bSGcO6tWHhHFYiNAUbK0vEC2JHZg
EFo2a4kKzZbYWsPijzmvweT+wjGME+j9tmX+D668D4UW9j9hxA42SsW1bGwj3eKL86ahIE/zsBUf
JyO5g4F8BS0VQkb5hg5MPjl4ppSNge58BRgvN0b1WtptwhW01h8XwUWZwVfPeHbWl6qyswjjbc+X
1Du2fh4dvG3Gb0dRZuSGyI323IvJEygFTdHtTi90iyN/+7KJx+gUylkmHfrqSY9QLHqO1PtjsF9z
wM95QTb1xApojJRQPOd5MlVf3tmnAnajju3EFx88AH8hyC7pY/Qsu4wls/YC03oBoKDttWe6jeS5
6yZCFz3mZckxoskv/tdq5qRd4TMNXbqeiEJ864vEnnFy+jh+WX1U8UroTnowb7WsuKnUNw15hpWS
ULkk50B8yldCulhaffOuRdq1yF3eDpYkuHINi8gwG3e7FY9Vi0xOOfDEDRTw26tpwrZExerGB+L8
4j2y+aTnJKNwOtKoWm4gj7j+vL84U7dWX/JT4FXfKlzkFRxlPy1BswTt8mVD+olXb1ZY9b6TKHVN
2JuShMTFTzzQVoiYy0NBhAFYVn1ah+/hgKPfUerwxo0C+vTQ1/XpuOm0m2D9tc9CEPPOYnWGwZXK
2O/qO2JZpl4rvwEeaKrCdPpnYNXAKnZNmnotMCnHFX29FwUv1/yvPPtniUG9/Y0iFKp5dxx5F5Gp
lUclZ36lMyG52RKtrjuZEErl/wW+3O5LUsIbbsjW+oLMjcJEY5hZg/v4fxu12UvFNe0a7ZuESovt
UMkU0g7jWFb7kQ+4tFQ4DQZ77xH7x/XgVgstA/DtTklviR8MTw9bSXfMA5rPx2azRA3bBoUJlFV1
kJO4SqwSbrtHVhUy04jStwFGivN7mSP08I0HxrBv/yf5zRZXsWt32XeDb1Ekt+jHgsx3owOmpDFl
T0qkbUjkeeGdccwNc56P3AEKtsztmHmeDdD68bIYJXm35pOiORo0p0csZ1hFO0onP5kHzHV5q8iU
havPIzuFFi5MVpDAGYJ3kNBw6eVD583Q4LGNOWao0Yi0u2WZ3QW2QhsfNJ+/UT2wOyqa2NgPVlpy
HjKAlWcgEKx2e3iZQr/ieVU/8/oXkBF1XmMPYcrbHWNuppmxxYz2TbzaNAfD/3tfIhaS5uzwIgkm
8SVr++Wc9IWPyyduky+S0Ld5lCZuCcE8vZVySpX4GF49GE7/X/UBnKPQshjb9u/fjdB/IIXOpy0Y
zWFD3GFUBVGGmVWFpK3wqwVSDNAt5kCWnJoZiZVtbmF7WvK1CqOXo+0BZ2TFG1KgXcrI0iT+NuyM
CbIhIiNuU+pLeY8C+ul9kXQ229g5fTOZcKGjLcr+Rf7PIpLl8m5On1ZL0S8xoUTulflTE/+2W5KT
ZUcN2jCvSiVNOpE9kxOHYSYH97FCbXU27qon5NqhJb/xlSAPgfWcRP72Xju17DOduc3JaTNMUq6E
H1+bA6LiEzcf4wsxkFEQvSN2gqdkep7oxpZe0jVmAF/4TSAd1SE8gY2Opel2KPqEteSPM3BG2lxD
21GUeP5ffCVjfUn6nrMSBKees2V7sYwyp/bcN4qnzQRsG7jdU5oUa34rhvuoQBdjfrwnfNdLAzD2
Q35puFSpWi02PROJk7Wc795eIKH9afvnuZ1NHyKsAHKTVhatj8c/lVWpoEqV+NM/Uue1GKRrXYzd
yY07/cDztl1p+RjsUmsWOZCnWtNz/zBC0ZORNSw+S4nRo0rjDHTjT57l7RxANturWNsPSRyrefud
geE0fL2+0FKRYmDnZhPhJqLf4j9thorSiyn1udPrWH5vxEElhEjL8AdnvTFfxLnbRYQPBRVmT/tp
fM5Hr+qpSq9g7cfonAXUXkKNYbd4O+Bsl1+B6i+O6trB90dl16s2np02YQAgq9OBLumJze5dvwt+
uDrhOkzTbXyfyT77s7MB6UBTuzhn1jaCH2wnclW5rWaMGZXp5jjfnoeHnoZtAgsMkpUqQxI2Iwp+
4Ui3SBx/8qsx44UX7QRAJe6/hNxEr13axm4a2vgP+yVheB4XvI+ZlLttMC/smVMU85/+vjLx+qjN
/1uA7i7rwF5A/9ReRz5sdthhSO4tZHmL0svii6RllLGA3cc9qi5L9T2GrA/5PmfQfQ940N4GzZfM
D2SoM58xRNTAPKOozZaNdSwVrXzhs/G011/CZYHSZlwbz6UExOgdnlAYDSAxildS2p2r+ofGSRkt
J83lbLPbUVBrKBYFeiF+RSoI+gUFKW9EChmnsvkQo2EEMy/RDmUa0MVZIzHqYJs2ChSvQ3CGNgZv
6mUWUPniTOEESTmElAQWO9tkkK39v9FsGnM0oDIsBxwM0CluyuwGlNy2kjzUYoQAfNVFEIkZW/XI
/IiDhdsS7A+PwpD/lG0RTc20ns1/oR15O1YStPboyxTPESXsrSm7PnTcWHzVyI29x5bF7ltZX24P
loJ4gjDCbVWmyDj0gOtGVH+XGTygH3o1OGp1qYnMoyH8bROvSyKrAZENy1Z5tzxe53psnyhZlkln
SZmajS+LPkSohnDwXxB2hKMmglI8GYTas1lFfgB1sE+xXlV78kRg/xljoyRAMPe0B83HskbygmlH
Shpdbk3kPDkXZXhndaNLoEJcfs/IizG3oXf6TqWfhF9MbQkrkjwglNbjIMeSzjfssL5QQVyouKBT
LkfWbwy3YccrvfKIEEtHMe8PJq8BNBmEvMwyhue/IcicEv9XTV3gfBKT1LNkk+uAfpI4RQJX5rq2
g+GrOglOd5PONv8/k/5y6YiWMXnVcQ2g5kZe4n6a/+hiSJfbrNVoCmeLvhWIAD3DBNG90Qhj7p/j
Fi5SCHDBsPnNBCgi1RQPTxCvOn7NK3iyev3fjB+/T2N+9XhGpNfSj2R0wLuxvXslHiR+6yamWCN6
HcukyER591grBrz895/QpZVF9gTtw0ZMSKsb4G54GULVkQN/KtRcNUd8bf5LtEIYVeK+WGw4/SbZ
qyTq5Mpflx/Zxdap+hkX1lqnIKWF5ee5MAg8gw4ZofTA/9bS5rPzWTO5B+6u5MqPBZrLK8zvPhOf
NOT8QDCbwWpD47rMYv12OHWzcRwFSK4FqeBfv+q/M/RIPAsTuRNGFCuXPtpVLpI1IrhK9D0KjLcn
ly8PQD1cfCyB7Y1+TGWGcNHn2Wcc/9I0kOvEuttglgo6GrNHWo3vullIzsN63SoUFUcinvdqYn0+
0z1/ojoMKPhHS+V0EdINXvMb+qJnYvjqbWxJrwaPLOH8HpxHA3eiqnoj1OS7Bl0DcYdhYErow/Be
RXXxJg9BlYZQqT+TGfzhnCElXA+It48bdOLDMMI0npv2fjNoXBkxadqhWcBei3A1iJZYtCPz7OWa
3kf+4gakuJvc05GRTdfNu6/o+6HVxFd/I65E6ZrNQxlsvyuXUfTAErY+7hzgYn+qiQMq1CUlWnnT
0HuaGurNdK7a5CcMMT8LnMJy39Fk0zOzBxkVsAxiD7bnEiva2mQjtWJf2jPU51EIeX4f4vNKBWFD
My1L1Xn80EtBboHDIB6RIHjwwTmvWzcRhCFAr5cCfUvAJb4H5uRysYKGanBTl1M4CP+HbGqW/QO2
W675IGFSEmhQERBZ6VePWA4C4Yn5kHlmth1keLoRPvg5TkpeZCsjBFHflvEgn3PMln69X4vtuyWZ
ZiLrDngS4/BVVF6kYoRxHsOILaFlENy8W+luGdrxYbkFfZJb9FrvWw7yU0LUbCU6NiLEb3mSXBlE
C5MG0GB3Hee0sBVONezlXRflsgE0F+ija364JEsUmQco03/rEHOxD0bJqfpLmQW/SVqfIswIFHdH
6puRbtsTH+BISS4RrkTTr5mPa6edSlD2Ei5479f5/SAp6bQm0DtuYUrGS3b/bxbF3KiFswQ4HsXh
fwsPnO27tEBoypOkM2Nr8Ejfa5hPR+QN/LduR8CigJJjyGvfbhm9/Mz+1skisngCxrQoSz6Id/lp
JyjQ7JjHe8/fNOlCixdKb25hhMeG5Xw+eiZVbOpRDA2gY7rPAU0g4tWMxBr3BsZqDhWUO/fJhke0
pzCtYE34luhAyB8p5eW+wLRbMgJfvOfChJZfSHsT4BOvNM/aM6zVzsYf/0AMVpbkzQSEcxYB5HML
9nToFOJHH7556Dwd6u28qqmNPjC+GJzY/nhHCzihts/H4Dxbsv/40D8xlRhhEtk1Jsdv8lZ62AgJ
uU47mKzysSeSUkc2OpBqzLzLs0OAuLCxw3ihOzhBZs+Mcno4kb++UnIM0ytnCTYMUTBDauzEjEBw
HZDNCiTOyKH7N9+DS6LNq1VEM6qXIbYaLDVOgU6+kwxWXMja0gPBrhoL8zvYfMvt51bTrrtSst+3
nzyNL2fSd6nHACGPTW2DmocVw5BmRGQ6I1NlAJ/ujRjsEMCgWh6dQTktEd68a73msqYf3R8vBnjF
IZpr+QzdSlgBrvoz//S+4ICTFVHvNP5rCdeMVF5JrwJMqk78p6GZBgdHJ5OEriwNmCHIF0JAkFTP
aGWw0mmKbVz9XTDCVGxg5YnW6LFnbBkJiWETUCYt8NQLs4fF8f/cAfWKRyK/bY4YzvSlbUyZIkuH
cLwAYR9zE7pMfyFBtkxNo3c4zkfdCnDqiST29jQEma+3+byLMmH/MSJofZXuKUutpkryUCaC6rNl
dU95m3/meDg1eV00B7kmVa4NJAoObK5+o2217VOncmoDhtUYcfYN3DpIGExssK/EtfcIqHf5EH++
3n6aYCXfw3gFay0z3bY627trRtwo0uDBbgmvn5hvr/Vce6+qjbTI/xypEuTwN5V9+G/1yJF+Majx
khW9vuRaw0AJEFyi721K7WeR2NhpEXg2dbl6iYwmz2uNjNZ5UenDzmoM5AlLpicpSG5UehViqk41
5Q4Zo6uVvUiD4ECfcnn0eJpKVnkLHUz0umZD05vLdh1l+F9zOcivVL+sGYvgk6YuSsCNPyOe5EhX
l9kcQSH1BMFU8kIIueM9LpCsf8U90nQd8r6WzMGaXlvGJUOPDM/Z52QwKPNX/Yllq6Nj7N1EDz2s
rDsgOxsPELHvE9oPeDB9Bt1QL24H6AFSIMBpicbO+miFZMq5XTVI/wh4p4/rXkwx8Jt252CyXv2A
hutXR8PME878bibFZZ0Bjb7UYn39O9nkaVczbR0ieceicFHOm1FXiOlN0erKU/qMp3iFyB4+1eAa
uq6ZilaAbB7lUHoTW/M/Ut0DUGjmH0UglpfGaX8P/UOxYl/H/TR1WdXxrX/C0am3jmfZx0DSINW0
6Ybn3241eUQft4720jvAuJjB6AxGpK4ISPxwgzcHUrwKUyczkc3mK/M3jzIuy12cXWetWT53Hu8g
zwgUSY4lMiVQvgfPDJoIye1Fsk0tQLJJi5qfBK/LVAbSVC0w6xWbZDA9UWHzsuJacqpKd5YgW7PX
WfJVbwpKEbNEs9e3szYLUoLvE/uiZG3wZgiblKHzeA1eMaK/t0LhtED+Mp3M6H1ih6/Im0aYA9KI
rmlbcU8OyYYtj+rTaWrNe38s73V14PnRKgPOAEiJba+LYvnmFGwzAhpxRoVz6/gTkATKCLb6SaD+
62NLZPz6ejENr4dvj8hRnbyuFRKrqUQAi80fQXz0dOGSPjkpznMCw9nEYJEj3cYPec3pGt98A/C1
YIMEH8ObP72/3WIWK7PfJVIMayYyCno8xCCzaEYZq5S+tbt4e6SzMjXhB+Am1R3pCobcpoYB1pRq
M+dT6N9AfvfS2ySawHjiucEklMOAkIJZGuXS2tDPYN529ekhpX9N5hVh72JJ0++l7u53Hxms2RPE
ERHTCeVcIkOGUcvSqMD2wjTqqIcXvHIY4JugBiiVgzjQ8vk1j5mCNsG6C9LfPjTgrr1bqycFoKCI
tLQ4uJkitir94dZ7esCL+hXmmx5hdnp/dztynNSrzpainhjW3SYUnI0OI1XEHhuJ1VBY3s+/od1z
fiZa9MU27RmSpFZPLfxMl9BbkMsafnqfApmx3/tQVcbwF6FLevlVPl6cwchwpvKO5F4NsNBeU2bA
0d9Rcmnrq8X/lP7d+eW0lc+E7ZqnIiCSYUKgD7kB9G+pAXU3Q7H43LD8pZyw3UwqpmZeVxfn4RQ+
yqwHRriqXTANi8ol9Yljlt0zZERVD2QvUVRqKGUlyaSQ5PgQcxj+j0eTFVptJKZigOb+60ejinsW
YtFpEumjXRLSyEt76t/mpjVxdsAiSKpQyJjcgE5mw1ARe5HXl5xmcgIsqV9hKSa+rW335mGRxeDd
6HJP5FUnL3m00d3xWao+PYF1p9FG17OSnkGznMGikviZf/JOv4F5UXOGsZPSnPJTPFPQXMKscg5S
n0ftNQS6nqYFNtFYExl4YHjCU8kQipV8zG38YdYuAaqhkYMsW+WSDam4IUyKvgbzzYvibfxyVrRa
a+2ChGorERbiaOkZZfhLqxO/mU3ZH3g/8jHjgKRLZjLYcmlje2uTmsgvt2XVe7tK0CLzw/JcKCLh
Z1eekohOfq2Xz/YXJqgZ/8GSDunpxAuaekwE7bC+JOycHYfLpomICeY1BoQiaxYpioYMRSN8ajUi
pk0oUH0+65KVBC2KLFu6lf7vun5ziHRCeigBWC7nSUHOBcel3TgdfMGgR1AHKYPs9TjwhnrwOlzG
emvyAj+4TbxAfBdt4R2teGeUzQRxEF+sxRwxv8hM+R83hN3dgupBlMEktrG9/XrU5w/0degwhN6Z
JvMh+Jw1O8dQXLWme4+mWpKlfsYPYP1lMg+LWNSBJ9FzLR/NZWKkyJ5sx+iAhyHWcGdhABceltkN
D5NdGFkC83GGmgdgXcQqji4rnfzGnAYbV7mHO2zl2X79HlG43Y96SFB1AzRlVEe3ejoQM+eQfprO
tNMIhseY2RY23fpWWIcV53GXADDf67QvABPIuEqr5BlLPfMLoazirsarFFkszUCT5JO9dNa0PIAj
TMKXDuZMFi8oKdBRCxh7EkseTw9GLYiB/vJDDeSKdRxhQMxK3SxsxzkpTGSvCzfAXIY++5PoC/zW
CUHXEG4dQxgNpgFlTpRucsstw2hg8KS7LHtgq6iTD0uUEocjC94hofqi+uJih96/yJCLBdSw/U+Y
EH0hNaIXYuWcloqN8HzMxuXRU16pHdeRtpPa7rJlZN4zugujLfSNI+zqolPa+S9WTK01WqGLnk+K
GHa1V0L06NS4unXJL7pK4d0ezzjgloaYcxw2PWGDjLTlgxJnC+WM0GFJFfRXJGX/rVI8FNJcwz2N
6az+wg2NKXbvwXjfHgx099J0U5N4nrdalLlIWFaJq8TGeo5waPwsH9y0UloUmYEgC6wO463hhW96
kqty5sZV4cn1qS2xKXoOnppHS28Jyep1QUxc1dn1uHlzudHv92zLXH5OiVMfgF2Lc9jO+4DMwJOb
FY4G6zIFjoYf50sQBHLDuAUrkguH/dezviaNPFROS24tYu0S7m0Gbb7zHPuOTCM/iiEzMs/w+veS
sA3lRKf+UgAD1n5wEIz+v4Hg16623OJaZmTKD8GvDxU/ms68VZz6MpHtDEoWGQYraGfb3MJZEi/q
5GkUVB2MEdjLh9Wnd3feW3ordR2fOENs+Zt66kBTtdltPg5pn8vkwy4MkdXYN/jLuGlpb7Qoxuog
qRlY6j478Lk+mBbKz2ypNL2W2eYkHsGD287JJe+9mzW87efKE+nXmzq5Tg128ePnVz3BNT8jS8fv
Uf67C1vfmLpQe1Si27Ui4yil44HECaamLoDl0me5O8NEhgBFh0gBHMAIv6iH8cRs9RlMLiYxWwam
QQ/KXXeiTcBH3bo8peHf3LCp3NwzPh/AsWmm2ioRKdklEvHX1l+RetkoKv5W83PElLFfRU7plyRw
fvf4SfpsuxrzKFy28ISAwQOcXx8rOg3mt0tGmeJMpqk/4XkofgA2LyFdGDKj45mInrxvRssoR0Np
4K72A59+dbwTStdFhslmyfVx6JRs/HK+i5akB+26eAPKeuqGvFtonIdVytdAjmGmVbUVQsUl5pOj
qFEQPReRs4Y/uTReaOk/eZGiKfdr8soPyj1pLlqp8iZaffU9gc/qkseGm8+tS0Q88HE+ZK84IivU
uA94EQcPGI3RVirW9IHMiW+mBA66yFSRdofRnMTavfihH3/esdSmyHdK1y0CDnGZFVzNOLgltgdM
PqxdVFo4VeCZpaHBSejNW5yqZbqsQA9ZPgEzO4b3vgBV9Q+gze1+tBa9F7nKsHU9Tkmho6Zlm3eV
4XBcY+avlPuOZVeZARVzKOkFwg8ecgrw306nMvEz5P+AFt9fXtvyE1Le6ZJ64DQARCIBfme2ZHhF
Wlf3Hx6I4vxYdOeZ1OKYSG5P4CE0iQMaGlmaImfjIh8VWaY3eCF4xshWSZrsK0IKluGgw90obb/t
VDrXsjOcmlsVjDw4idv5rFHNn44WFJS2ab89tC6dEJQ1Rrf/KUAKzCW6tmsWz9cj3E6hH+j50xVT
dR1icN6y/RnSmJSUDiiaOw6F/680XCP/OatGlm/DxJaMXPTSuddLjjBb9LJ9+Rq3MtPRcbwd61iE
3mKpvFQvH+G5jbXQnGYrxKWOxUNs8nov3pB2jr8NUlrm7psfz0+3x36qInD1q782g5qKqooFMq8L
BKG6rnLXee/WfixVvQJ6p6njqSUTV46O/wg1c+maiKxSt9J0R1wx1A4aH9LoW6XB2qAh2lx7nARn
KpMO0kDFocd+aSbsC69pR48utKubYUtp0udY0OW+HnT/eH2M2968eIxoibc8J9ip4PQPjb+pjDw7
r9R7ZQ24ZFrVkrUyr2LTIXFKNqwyS5apeDnFsRSZ23L6jYwBE/4BRlll3o1Lc/9rjeGtaW2AdVjI
NajpBhXISaVaYPl292B8jum/1kRFXPAUqf7Fk6iZ0oF4gK+9j6uAZFW3raia++RqKBSCQR3/euTX
wLGZX+/2CmX6eCAnQuZ/eMl7MKpcPwjdxTg9k8a78k8Zl9VvsrHOm31inlAGAsIDaiW6tssT3OBt
0BqZ+TcFQchP5dI0p03bCUulm2c04aoeuxrvvz9LUg0TKtDStvO9ac6iiferF1qWUbirKmQJwARU
z0Ia/FbwiB2AzMiCCGwjBqe1FuowKXFHXU5mG1ZA+Q8aRtC7bHQWEll36DceQEuThcaL+60aYi99
xNb8CtsjUVowmVPo/HU38VDKHErAAxtAKpCEvaOFMpJ3Pc4ikh+ZkqSQvzlwetItR1w4WGAQpLpc
8YTafQAGsRhoFPwGjfonxAHUQT0T4gewu49VjnooaJvoNM2GkWTgfSvrH303HIKijBGiHjnKo2kg
S2kGUQMpi/4CD5+GAewWhdqXKgjPJvswqiz98hUUT//X0qcdJOjv0URhH4DkjzLdrdKlk2czZUjy
KMh2VN/KOgaxvPhRazVm2U8sOMh8cm2djSDkaar2+xxmF+0kYCTAyTVM3NNCRyl/PPNebXOxlcb0
tjUq/58DBtBDPvTZ+0pVkkFOozZC+LD0xtBUKPl9W+JfgCzVj0TNB40g4g5KyfpHahZk4Fb6ho7U
yzJZmImzJSyEcjpQxWcEj9NrSwkwua0lqyZeYlx0+96yoQ4LPb8AfzwoYh9bMz8pzFSLkGSwEkc9
DLosg1Pk8VpqW+/XU88RDV78zcXcBjOs5f7Vz9yBuXNsBL3NyNrScWClfuM/yaxyQN8KX+rXGW2N
Y7aN4DuFJ3QMeGzqeoAZKyrYQehu1Ru+UYucon/03/XBi9j0ON7Babf725S/lTlb806aFOkfTIQ3
gXWwzRjLbJ4rfKLtLoD49Bm0ibC+G5FIbTLkjlfQiAPECAhagyFJpwMx/ZZit3FMAGMkAhzSBLAp
DiOtSJXi3LrnlVq+NmtAkIJEZcp7ILzPMppSfYWzg+lH/Um8L3G9Rncm/XJDu92XRYXlM1MUucrP
bQdqmTgBWsrm+jA4ibf8M/bVvK/RtO0O/cKuwCt8sMq94hdHvNMg+2lzpHe/rrP2BDxTEiwU4wVp
UoYUF81B+f6CCe2riBTf+1rCFRXSs1pIl5+CL2hht+8cOuXGxIhkl/emC5NXduVS2c8R8j6mnpDq
w6DU9qk8qkwBBZjSo6V0P+BeQp1kQ9wTeVXjd0oyoqrNtH3lo4IrWIJEUidFwqlm7/8gDdfmRfPU
nsCKOgHiu7tEYxlAXws3sy1czEk2DRpvRePUN+Bv+j+WklWahBplaQLRQXQABssjXU4PCpgW1wIe
CnPVvm3jQWuBvgYi5ozl3MPv9jHSoKewrwhlyKk6mLIZ4TMfrnAnTtSAVHS/NaDpG2lycBWyz+up
KuTExjIhARVI2aUbzi6MDfPH5Pwpya9W4iGYVpNGquUFyrDav2jtN/n0UfqFdCE+aZVXbAopQgb8
okv3FRwSU6Dt6UA6E+5tiYKBo3QuYPz88sUPc2UJRXEMYHQ/0KfrfRNiZpkVxwNqW9xE6Y4sIUIu
IJW3QUokS+/YayVMHDI7M4j6LwJMxUiRGMPOjD0GifPcf/y+lYHZsVhfU8qHpk5U899dVWcjnkdw
eUeA8shfY3kxDkFVxpZkeespsTj7o2mmjwyjSvIQx7d1geVyI9oSL0tzFy9K8aLZp5fmctK4fs9J
b1vjVGZ47O4B+fiCP/frK2Nz+B8fLduYc9V+O1py/2LL2yIRpstTjC5TiRV2PJSKp/xzsVlCAG2b
ka1Z3kn6VH1RhCCN+a8aU5sqv+xt5TJOuqND6rrG6gIlQ0vXAxUs+yzQQNxj8jzovm46ExRAXQ1e
apoQdVoN3i5kj7aEs+8r5uJYwTwlkZ8Uzx8+tUKErkrsRQXLsZZvdFotNyMmX/FQQ9w8aHGZEjqf
IobHRSsBX7fg/SedqrUXcmG11quuKB77xJl7UloynN10Avlzj0ihs0KvmnpAT6VakBsAmQZ0Pse5
m4FF3NSUayfU1Av4rzyISSdWt5JpTqwelTlSagGm3X6JXLeePHkL7UiIR3RKE45TE1hCPdgEbcfs
u7OkASDr/Eb4TL/V38ABeWDqnTMGQKF+2X9EGF2H2XDNZ091RWSCiyuQlXQ2D15eWELNP1nLB8nq
gzav3rZlGTDhp6PWEtGw9QdSRvfx47KSvB5EMVYiGVi5nC4W6N29SK8ATx3xV7T3CBuniTrQ3GyU
ZY+UlnLQec766tnHhAi0lSZGisi3DLuZ8JqoIpns9ILUV+XcXQ7RCcqQeHvNDx7PRwnbeoFnCPrA
6VjS01f3XXXrcXZG3GTlGdrQaIzoM8NdESYp9XiuCVQVA3QNS8l71hQBFsFOyJ5NAmtfF0Wzld6N
v8WqJKs2Nh+jcrA82JyMi1wwLR3+Ikk5I9OKzgKiaSGMY/Vv7OcZDK/rcF/n3OdP4X2KSbrWUWtj
I2H3ftYPlw0pvneXtPerjlctGoLVlgRcRpOiAqGcRFf5C7xAOkGXJZ6SKc5A7F7ryRBxOvsv6j+n
HkAcx5VclatlSp34X8GVmN6obYXo4++QOqVKcbtERa1NY972W3BznomDPHtXnHkjsqPj2IkEQ7rv
XrzjMqfA4c29k3P7XZfEfnIODIpBK2TZR/uJy3AGdLa8XQt0KGEX29HFGBQ6lk5pmj/AGbnihLHs
VI68GAkZM2wWfmeE0rGwYMlhAIu6BvcJO6XWAh2Lg/vgvK2P7sPOI1r+x6kYHHkX+cEKQVCb+wSE
w811ETdIg8OQPPnLxiS8VqSLL99vVWLjQhhp/5GH+41HetQhzO3XoQINIKNPUxl5tfnZRFUyjtZ6
VCUZiKRcgGDiP40BNsLMz+ZyxCgeTAEoDs0NFtT355uz6EfHctGyvY3fiipywgzkc31KlCGYX0di
ucW6vOL3NPCbMHuHWIIBmXlIOTfpXH1NrXlqT0hO4nBG4kJvoN5JUqESlgOpXMgf6bYOnukma0gC
O86L9uMP5WfFehYtU5DJpGS82RtcYdRfugi9Tl7wMhlnHtZ82vPXzMho1lTwmzTlsGW5iFf6cDvf
ra9fa0/RXl1IG/tPp3mst2f0fC08ng7zphTqlu7vGVcySV6RHn+JKxzQaMzHgqDhDVSCbP+b+/sS
N84m1Lk3bBwJZQfp+7t0cpg3UFNh0zWqFbMn7GgJfoNvOWSk9sng1ya7n8CyFoTNLfRVhDNFKMij
uB/HgIVac4eAuzE9FopAZO8EMRAne7TL8ZF2Lzy/h28qY0/wAkszZ/8taTLDL1NNxr1piCkbixyy
b0dMwpEYigVROVETj90X+iMgE76wIG2ljekdkfDB2cK4RITxBdv9yppOVU+zfZxKqiu+2butEgqk
HY2dqaBFgLVCZcODx5VlX5EpEAb6bLJjK2rZMnneMX2x52r2JHCzIvlIF5NK+wrodQYZ2mbHNf23
FDZSULuzwNQUD/gzdcKjB8SV0pYs71XpMorlEumri4/4n2ytWO/KUs7rSuw4rYVVw9FmC2ZkKbOQ
qL4Ds7C6sNPWSfcpmyEpx7adUly3gB+D1y2Xjrqe/t6JoTwoABY/5oOEKu6koazYWYKtwM9feGIl
M6nUVhecqrF5Kvcq+TQbdnqNphu6/Ev3mtaRTIS1wxqtTBs5zkKcHVGhMFCxQ//mEipbHVEMUwvs
I6/OzHEokh84A2emmN1+qD3yotkYdQw6Te8GjT/4NHyErT3sjz+ofAAr6YS0Qg5FPs0BvjD0CitO
eiXS3Sg2C6v5Gf8jcOuS7EA8KUcmim88sXJ2WciUvQpbMEv+naL+EkbsgM7Et7Pc0xX7BcdadxZH
1hF06P9sNCTkLb9j/cZs3H/TgTPdUR60B9gQVbfwFqlIpuKOOnhsjFlXf6kyE5L1yR3urI1h734Z
jvHYwKjKkXhjE2ek6VxEOjs4mDAEYLMzdiIzqERUzEkuaqKnDs6F/C/TmPM90Eq/H33jhSqMAb4m
YKPZRxX38M9yTR7O/lxLxtkRecTrhBPjEad8ZtCcMbSW5ayBklWA/tAtVDB4WS64+SDymTWj9Lk9
34diCz0wOCDuxv9I3Y0J7owYP5jc2eaSJUj8/Ww7vY5f6Z8ewwhajvi30bKb7/hvX5zsrM9HqzXp
FlFaWHKO095NLOqMFHFDd6w2dBgjKg5dZ6IxrN2z65Vn6RQ5PoLeWNbrp3vw7o37w34hdFC4UHUE
06ZPlWn7f55uvc9rMBty7cL3Mf4a5+hHAR5jXA4unYwG4+xUtuafU4ie2GUfPqf7+K1JtOA96ecE
CrxqRIALv7aOW7DNJ9hxCVSJ7nk/uBK8YTW8e/6xuMNBnnaCAAZuYIVIqC+nPv3VZUEaPdEAkiKF
uxcd2y3oAjHGEGjNdyXGSzsPDkDHdk5OZb2rRR18JkXw+YCbiM0hBwcaXhzhMBqQd3AeUk/I5Nda
hRM1xMw8DLzl9av1MihM+ud09VXPo818ry3U9KrZkPE3xiPKygGkbRDM9fh8MgunSt18YjgCW1mn
lbiexPiPG08a/haQsebfewnQLvSNiAJP4LtQqgicO4/gLkSPhvGuOzhjIA7ZIhHPl0+YVLeVyDTs
IEcmC04Ri4J6x3UJmXvrUxk2LPjyQ5n6OrPUzRZfThL8ZrdpidIetg9XZZo9rco1O45e1biV6dJR
Mt6cHbZSVG39628TEmHE+lPVwFdVrly4E717IApxJaXBEUIVlc7P1mGw6EBdrTlH7awBCn+m9CXK
pqc1+ChpWuP1Xrru+i9MqUofaZboVOki1plIK1uMsmVHvKNLu5uC/Iaz6WGFYGdLBH6BSYb9Ubns
hFU2KeRTHoKF77l594pS8E+KwBhN+Ew4f5zLYERwEz0ESVziikqedhKiwEPYvy/R8XZx4vwim2YG
UDwl9Oi972T64HJwj/EJIwYtnAxrQWdfqiuj/CnvCSvz0gSaT0LEM2G6joMF9Wlcmu34jpIFmbFx
ugQol6MCKi2oiiuql5A0O7IzRN3LgZwAEAn1rE+v3QrDxd6kjz2Tvrgd62V3ThtCG9ohhMvleiQO
YlCRj90N1N54WHU2X0Dw8uvSWYE153InE8HaYAxiIP5SVPsJl72QCOFWwwR/BRwHQFrDwuU5xc15
e6DnsOjrXZiy9JVC44PGdp0oxuFSdMfWyvXt4dP3zr9EOZAFquyBdLmeuPSvt93MTDslJ1ruuVg+
FYOpTS/K0iKCSONqCoUuecmWFmHOSFOJH4iRPA0K/hs3sZIZfZFUqNtdnWRGf8dfQBHYMF8IRbOc
LfOFf5yUOFQXCJLTIyKSlrPX1RsPtqUSv7xms4oS1IXbZs2nfnUG+b/wmwDxRSTWlEFBZcE2fQez
cwdeRsJbpwhqR++Y1PEsqJppjPgxsF6wTVV1anlSQPHlk/NRYRvuqKl4ymvABo/yrm0ISc6VUViw
wKXt542rCV5TmPTKVrkAFIQgxQLR9EyrkiGzh7zF/4/rwuATzCRbQbLAhm4hfrxr5Gg/zw9IiOAp
uCIAkpacwtMMMh5J4g6d8hV0HnGMcw/HLy5FLgwBTTA6i7IdDPcTY1H3wjSFfyGckbZZkSoOcvuu
i2TszSBWLMHUAc9uilAF83g5aSp4sgUVduFFuiS6cvCv7QTjTIGFv1HAKlM9sSoW1ruoyqun0WUJ
LCcceVxMIHguninARpp678g046Uw5XA0QGQ/BLiFIGiY26BGrVjJXbj0EhtBEZLZO2ntx5ADlLhF
ttcIxqRBzD/15x117dVcdpMWRzN7UWykXbJi4jGZPRIoXZ8W8NEJXf1uEVvAH81P1qTPOH8mf2u+
YkOjb5wlLAkwx2Zc20hlEWR0zEmT6yBAw2OhFtCZ/6Yt6GiL8jzC9k98X/0wNOSCXdhBQyh32/Jt
3NVIjzRUp8ylcKUlaJaKn1kd5Lx2qDyMOO75aW4eK9pOzZyVqRqIQzPHglaaFOm8ysj/qHE8a2Y/
j3h2Rn89TKrKNPHjYXY38wzgPZmmy7qiJ7gmEq7fajYD0hTYkpxwNI6WAdRzLGNoecJ9jzyDV26F
hIIDYiqmq20vtz/5AKmQ/qVDp9igGER1laz90eK5SDBmzP5/uz2uUtT17tdpzqphMWgTZCG9Y9Q0
5hrUdlPsNbZkamxNOcgT+kTH8mTVXcPWhR6DZKZ6JFAqqEb6WORKTBaNi/JjKCfXtKysddZpDX9/
tEk6yoe38PoNAOGw/8ZNpn6INk1pVZnkbbqyJ/wHysejSBOMgwQL9ViT4BPbbSpoJ5r3XIRLXI6i
bLYkk3Z4d0ufe+9yrsBgj//BHX/ykknYsvraB0OKiQIgFh4T7tODBIdC790D921RKsf27UVwU+BK
ZmD5tgks/a+8y92gwOQURIKeoLhHFzjtHlI/DpNMnW0eGlYH/5KYKiqSHpyHY8A+CWqAM3hQaBtK
vhApxSBeMC7lxlkf/54FjuJ5ZzWJvPc8oOq39GXZ+haTdL5Y6+xPltonJKedJ7tusdC63SfmgNNQ
GyJeQ+mdOka85rb7/A/wBWuM8rMVO90REffZEGEYoIbpUSEDy1OPMbDMIJbM1cWjDtLyWq67na6l
q1g1AaqYUjcsNztozxZOLfaoAsbtec9QeXkOq0zhhQwsEtiXT5YDLweUi8uqo53dmO71MEWZpoPO
OZsZDtfkXym3wS8ekP4BDMnhVRx/zu+25LJOpXKAWdURnazzX8dfrw8AySmQ+6VBo8whhaqk3qu7
MkJV3htS+6NJldDkaPF1lHt4Xgwlp3I+hyCIKagwalhYF0H3OXpDV9C/YbgeOt9mUKbHRvZJlviW
ir5QUNP435xQM1gZaXSi7GHDL2OE4PWNFMxjWFYEUzN9t0kGF4Yge3se4jeytnEh9QLgHJSAx8lG
JjM/v6HapPCex6eT3vPifbygWzbsdvGD3FgsRbmkUWDOmOCSMa7PdZlKcIU3Qj4CFxWfMHjXGWkV
ND0YRhuu4+XdXeCPoHE0zf7r9lnjpRk/KiFyiLuoDp79AlsyrF301hihJFfWIMJEnSb8xRcbYCRA
0jTRuotbJTPz+35Zg+DZ4etgnrKMyrVQuGosNMZR+HBwUdqUGMXoz7CKmPhvKLX7kodhpVK1RiZl
Vwl3AnUxjSRecPi5c86nCwW390XpkRjoVgVjLc4I76gZ/7LtrsYoE3eNH676ynZjLejTiE44PVwc
8BKnkm+ingX9P9ugNBloBczvsXd4QvPkPLQQZGYgozipl3ykvIxvOt2UUDNBaHWC+j50uOR1C/ng
uQk3zLOBT54oV1JAhLm1c40Cd9JNjHgdFLJBK6xulqKRAviQ8VzNgMHkxne5uBLESMveG3GbIoCt
IPCOxjeoPWBzqXKRvhWEiAGxIkv2l6VQNmqG7e8tQUCgAv5e72uJaOSKM31/6AHJu13QAbp3Iq3H
lNkPFozS46UJuD6F3zolKItV1TFNOpoZ6fVBxsItCBTCDmPKKrideUHH/xCAK+Ldw+EnVtmgWBgB
iS/eOM+JmBl+Iz8Dq8UMtjRFWT9bgzm2JVxvap6nQmehnT6Qz2sCME1TfDc7kLczTlv9O6JaOgA+
/5JlYgXmFF88R9HQdXF7NuzFEN9aooxeLlui/C0hRMSHCRXICHSDVf0P/0X7n+RwKaG30as8Xjh/
p38ux77FQdxQDe7jtbyM0XgBk08rDY/gpJXKrlnUG8M39fPa5LR3fcOSBjHVNuxfg33Ctc/s99VG
8l6LVGPUHbwxnxpPsAqFO+J4m0LMd73U3bURIbKzoeHb8apPCkOHkFlmF+DP46exmazpf+v8ttvt
LXOkGmkcNBrpPhQp6/uzzAh1EWoUXoiTQ8EvwTFUvXnpHBk887tsMDqJ3R1+H06GPPuNs7Ag8c0v
SONz09wB9+iaZiVGFcnG8FszsS7HJLXUR2a+7F+4YEs8X0GtBmREeg+29KK6OyTrPNsyzcJNfzfW
BTmSxyWyvxZU7QhiPAOxEX0GDhxMs1YFhn0dN+a2bd8mSegxvE2COPDgDFCxCoJHA9kdG7m59mhk
qOmVUlOKF3qqRizXi+h4UwCkXBvnlfxV84mUh6DdukYRYZS2hHQgDREAi3Lh1sNfeE6hZfsTbNhV
irjcyIf9twCk5OY7drkqsr/ALquBVVqr4+KaA9awQUOXWqjprycjCBmKLOnJvCL/35PGj9eoyREQ
BxZ7jfBISFBMaovKVWV+KhcXvQo1+eoGQA5kvJTlJPEmHEuF3NZ8pQEaW5V1Hg2pre3L759TpkYL
3N0Hbx7AHuGpKDeNb8rjyEV32xpPKmpj13mg09fphtV+q1hatBZ2Qb22MbI6UXEGC985R3mqXMfq
6IPGcXfCFsMu7KIFGZprFeHbvkBKWax4Etgv/8LZKtiqIMGX6pFSNuAP5PjLSXxj9Y12Efv+Z2FK
mDB4k/kDvhzTzx6RV9okVy9eXsGrWce/giNGLAStm+4lU1691HfklC9XVQEnMXYseQV0kLg7fG/H
ebc098HiNIdYBZHC+sxHY4hIh0DovBonVBYsa4+V75QYlDUsNyjRLbI3y7XbGW/RUr9DRuccINUR
CQ1QLOv+wicXx0bfyR4DYuGHmnaTaGacYqpzYfO5wf3yRQL3r4zrbJS7SJXvtF3IPNQQCpaxlNNz
k+nNwX+JUzsUbdrwcRyb7sgV2kORsCpUsCKg1X2kVftDzvQ63OsPCzryR7yyZH8rM1uO0bljh0oY
YprCK81JzotCipvIPHWX5jmFQpKrt2VHM6Rqg/5zJQU4AzHWZAih+u9ZaCNaKh/e4887/WX/tbAO
RlwXN6OBTUiemu1dH5lgcwpP5deskwiIO6WCTM3kImTw6n9AnftIUJWER8FBVpwvT+AzhbCAX0Iq
HUF5b/Gq72rmnVK7XYkF6Y8tdS7U17qrkrg9uWFAVjExBLhV10KRC1bJxmz8O0Ijt6bNtAy1mrGg
QhJD1tfcM85pHoB/HXiAuTY796Vsfd+9ggG/oxH9QfB33dCHqqpp3RSYOL8YGg3WZqjgEO2lYR/z
8h27TqL/xNQRsbqWnMLLz60XnkVPH99HXuSiDgaWf2MyAApUmPgNmKyUeVrRhqihEs7DTr1jDvud
KNI/Tqk48PpZZbKJS5yhBxDtHSOgU4fRdcvMIHAdofgCcP4RzIc9vA4jWqs+cigWzSFjUh/KVOVU
9xGDUdjrcCjpK1brxRGfGSAQUE5pMLBdiIz2cLKJf/xYxM3mWeQHOCErKUMyAjjy2LnPx/54KX1k
+Fez2OWc4k+FNvGwMIK0/9G0+9CJndIHvRWTkXjKcwJS9nYs8QhDgza7ZzuZY6cH1NB58EyQbDBD
mexXMYicybSa1M6XysKWXclyPmfZQAZAGF/ass/oDHL+6+OsJUz9N2JMja0QOcblhWk5OLMY1SH+
Pv89i3Huy0qD/+U9gjE0zu4AOhvIpUzaAzyFC0e8oX6Dh07dHMZUVAtXTdYu8aFQvpjrlyProJM9
4XCqBgr4NtvMAyv6TMvH92FDqB/jk7TuyqjLrESQUTmPSsSuOttMBKzcbtq5Iv6jGkkNY0zx/0zr
4mOSH34Bw6NcqSrJExp/PHuh3fQOA4cjhKC4v4VgryeHKKTD0Q6VjPAs9qqrUyuiZRhQaz2G5BqF
4nQiPitbk0RBWkKmQZaffsTP+S8fVJyn8r6p3E4E05WY+KyDJof4kejEiV8zupg0gESN0e8yNZM/
0GJj6xg81H2orYiNGg5QP2wgoeJx5NIXXbLRN56th6wBSE7c2QP/HKnDf3Snh5iTxOBNuLAhZWKA
jRClHIetvi/aP3ZOJcovF8Bsih8zGD3zRgaHWqSbywtMSannkwIxDYU+TOTuyhLJHpajOtu0xHEu
r1o2OE3hwUWO5vwr0wfRyxdD7q5ZkM1aPF310VPoh5QDFraRxz0tsal9K+mT4hBEmUQlBThp0S/h
ZvXP6U4GE0uyPQ6ACAvX9BIkbTdMWlmiXxMSf5ktMjFmQMueUwM4MO1PGik4HrUs5GhXjE3bS3AW
9DOPs5cPiUmn0fiD7q+acsMECDvjwEo7YvR/l9Ez9re6S0k4iQvp36AgdJj6MHTgWGtqV7PgUQIR
5Hoj2/1kljwExZjU2S3i3Sf7vqHWaT8BWssTNNXAimwnmiOmujM0tR0TONwSjM8jngYTjI/YFe7a
h3ZZXYtLpa5IYQMlA4lsnckOdUOurLFK4bA9+KCh2EreZpvJs6WlwR/NXLFrLfFWEfbjcsN3qULJ
fo2sSvLBV9qNgCq11+T57CxnkJDKackKCbxBW3MU0/3BAJWg4QEV7Y4TMx7ZP0CBr4ADfG+rSe6R
1ImOJyuHMFPJOOY34ubjwFeMUs648hgolHVXfp8hmpKaRHaDFH/etfIz2e1J1wBja1FOnZSeIgx4
YLG+PtrQAI0TrzAHcgiyyTkJuPcNjYdrro+q05euwUA7leimt8W7ywZqEnB9dKEYGfBSj78mReNE
l5ArxXslazCP3kdxfZCHlxyEXIyzOMo2V5vAhdsRcvENnNtJh2/8bMl3Kfb7x/HESOS3xXs0iaVm
I0dndepgcByM2wYrWrzwNK5Qa50oZV6lV0UF42swTFLGGVOUz4knlMLlirHELynrbEbiuIV/ZMCr
T+ir1jeK08oW+7vxPjqjFXuZSrGUR3nmjTlzU1zBHNX2usl7Fry6vUEwlNoehnVfQ28/a9lDkrPS
/QRryU6in24xTrqGyMzPJTDu3ptK/ipXM6eg4Qe/F6Lll7X5/jHHqNuJ1xi5lR2XvenFv0E/0sSU
fjIZ8oQp0R4dsrnwqqK5YxufWolw1WFk9PmsTWhCijtN41Z5exyR5CTCu7cwEhcsIGjFBsTYL1s8
RBxs2skAbtJlJYqR31ckb8sodsC9NpPXS9fEEP+uhdctZMcm9XcpJRXi5Yv7eagImn6nDMXB/FWy
O70PQARjAgG9CTiTdYehKMZg6tjQhfK584w93ayHJlAaLgSu7SzcKPZwMCpLziSMo9gnXPvviXIv
tcIyekmJaf+9oHVigBwRArwDbjoOqUsQLrzW72FvkkgrHcLaXBwo7dI7oMmWsQVczPIdOrb31eOW
Y7c5dKDNn8aYSvkFuGVn7lRunpwrSZccEa7QcPUA7GjYpvSPEBeNUqoXD57ntCdjn0ymhvEVP9fS
IC8/VSqAWRMjdruTOjDZnksY/d0IIQLj8Enaf/dvOakjMMUIQfS6Bw+MoQquKBTaIwQVupVTEXum
jaVxH07Ry1Ru3XbXtEbqRMEoSOVU24v1PJZgJgFbSK0L+NZACA0gjEGNzPxTfALXQmhCocW/fZoN
cy3Dr1X22FG4q5RQP4F1Rze6JTqgBIW+NxQve5OjMHITeczWmPyp/cKqbn6tYY/BYBZzASZ7IJvR
CdDmj2pKMM00D/TQHutsowJRnC4rTvJStml3ZTOnMC48Rqyd/NkRkNEYhpk9c1bCWCf5zkUMbahi
K28UV3WORG1KoW6ilRgm1EEIpBRtHWwopfNQShVaGis8PLF+3sCYB1zfgL5Pn3jsqomR4nhWH4WB
H9yQiZh4GoqNWxgvkM5AFM4DEee6sA4quY/CGDQu51US7yCol9PHvvX6PppcsTJXOiQyswoh2xC5
UprGFpWYNr/poyVylEYzAQ5kNXzIrrN7ZAM1SoQpcMYNHuSf3Gp87pI7wkcnm3MaJoCu8zF0T8k/
2tOchFg3sdOzNLNkNFHl9+OSTtu/hKPg2NsYLvCY2FmPvY/GvXUojESnzzhw+BWgd2A3s1GGHJ+f
N+ONKZm82Vu+m8smfxMgcSO68KK6HWafe4D9ze6vVGNwJ8aZG0PaRgfaWVwHk0MTiLH/g7O3X21W
TROZNV4mUXQY9jv+AFwVNXtb+wcOdokQ5aef7hUWP8aNuEZHq0Xrn7b4/AT96+qXWBL/kGVJLVAs
oWGopW3EyGfPiw1wu2naS+E3OhbXy9XlT53crW4fY9RYNj+tlbIj2toEGJMgnUiy9baIkixDYbGR
TytbCeyg0ORV2Q60eNLcfSLjCavPm613KptnB5j6VMZrCtPWySAnKKZs8MfnNA+bTpw1MMGVw55+
ifR8yceeBJMrhhxSM72wPMlNSgLR33qPo6zkGCgPf1RA4jm7OT31mO0X7NRT7Bb6gbgSNA41F5XZ
1rmrUn19u6OFFHfunwJwlyfGOH7C5Y+isJkR1nex68lXbPRLrjOkD18NhFThPaqS/RkhizRICPer
+yeh0WtPI5N3QwIujszJbdSMEwRnHYfvJ7c9lpOyYYqVYrg8K7sKikN5cULX521MAFpn0vvvvLRE
LAYtZF43kpob2VgjDHksZfdKRuZvSm2BZeeZOolRqjLJ9RqsZh4c0R2yWkNA3SgVeo/V5aSss0Gh
pm91mpGgau8mi3n4GwK51Tks5/53g3AvSBqjarrMf76LBy/hEomtyqMb27qjGomkIeIcnDPS5AKH
O/hwtarsTx4EGA3axFzp1DD2oi9n+tHyL1B2wS8wRspuVwPmhgB8mPuj2qWyCzF8KepcLA8Nq3wX
dQLEKePkyGPgULy45POLtxuoNJvJeTRT/JUl+hv5fncDmJMb2KHaAot3QiXCkNtTdgbdxNQQuPdY
oDNVGdjU+jdVXdGio4u/bU9YcTPUC24N9IRLkkWeVRnzHc2LtzjyqwA77p+zoKck/NfUuyOwzAng
2XapAI18PIva+5oOukwk6RFDfwgXtEbK06wWR/OsixQMbwiqEHF11REf5uM4EwmnqaS+qXt8p2HY
ZdfHDoRAnq/mCwRxRTkGKfGwKVPl4k4uRKdFhcL4NnOMRCphb5D3yNyiz4WMRTT/Eb3MMJM00ndG
Ir8h9ZpgJQvst12GSEKjLb0ou/OcwUGsc3qkCTVtocJlRIkQnsT8tASKwnZp4nsQncCJRg19IcK0
J7nazZNbNxMoaNqdlzwe8bXstCnLN+Ssdd1hjCSx+MMrx47tFSxUzBCmSbBuSNi+JmgOms8/QkUg
WJ+0kmvSFrh0FhKRryStMmmj7WRgylnlWMovLYk++/drB9xKtDqujOChUJtxvqJtS1ITCEEbT516
6bf2/HX7fOI6rUy7wSXFjqupA8E2rLeJrZA/cgeLSPFpfh/XVCc8BitD99NBPCt1BmkAtst+zt7D
Th5etAOxjG0wWqTutkLFFFwEyFb1LKVfjCyxQOwQMIPVrrNNMa0FEGop4TS+nZREGYKAVz4WLraM
yOXYrTPTRWYnIO2eQkkJ/ZYHOJ75lfewwqcm/esSg6NxrZ2UN+Z3XiYsPzy/o0OCqA/WHuOcvSlX
Kn6qXjcJveS3U4kV8bO1+nS6UhdCrdL/EB08Ir+LddlfljG7FZ9LIzOJZOSByCsZYTkduMBSC1ld
FFfDQjk40/cd7GURhHwhBLHcEsYXq6VKLCpMUoZedE7m1+5ENFx5t05xsRfbwX92TvYRopPJATWN
ecIaHmowWLTgrMgLApCtvTgE0YobwPW+Y6ciafsJwTXpQ4CCzwROENkGH86m5VST5xpTYjhHvelc
l13jZpZCsrvL3uoeaW6RYqOUkr7I0sJ9uiSVP2x7vGdSmyCGw3KqnqfeT6mn+jvAtLehcsFwcFJ5
9uokpo5kMLMhUjRYR2U1651bhjNwlhpuxC41BhFTBcCRAqWZbmDjlDZ5h8hpr/5JPhFQ35ySuOfO
U71CHG7bMxgwMe7g8Vo8w8p1WnJgGYA8R8T/yz5zDItSXvZZpQpFQZr+JYkSEUU4EaiEn8/t5+sW
+1kOg9rZHUhC0ZTIIddw3j5NCE1XmPnPTOT35RgOKH/rpvkvW16sKgPElDTlbt5rQJ5u+r+1wm9K
r8zNBFZMkZ3xpzJIIcMtjncOGmBqpm9/b6od2h13CzmMvMWkHrdjNHut22BYLRXCMuUSeycoMCN8
74KLKzzpjiBlpxwc2hgbENp0GyzcWFAJXRTDzag1rBZ9QcmrLLKMUV1M0kXRzKzyLnb7L1T51dn/
svtgb4BFCcGk+YVpimVVJLa/T5PRj1Ij9qDOiv6VLyfkOU0or1WEmL8cQ3gTg7hlxkvkeNZOJROi
4naAWMUYjMvutBJ6pNPNzpq/XIdV4PyjQGSNvIqE+7p0ULCUXP3AFHf4jDcN5ujMBPeAK/Dn97OH
21Po8DTWQwCqZIIUHGSxd8F9XLeQPNzb3Mv77tQk3jWlG6XAe+7FKacoOup2Q/UkkNaXNehZJUHk
HrvFfk7Zdysou4epjAVt99uPM6xps9fGExobAJdzj2bgnuthppaveQUb/zX3kaYclhXKoUZojpbi
OPYK4cGhqtbybyOdqxG8aMlXLDXpZwNd18/xXUSR6cKLroadFAkEx9r27qLeD9W/qRTrGXBxc238
y7WvZ8MIPZ5uECxEZDtdMCfGVXyAl/7ASBwQLDNDZqedDjukX/xjPdUQWkibZDqe6IhlSSAQMDXV
DyfqMa0OtnVKFtbVqgeMCCZ7JnBKyAkOgLexdyuF5KfUdAIMwOXJcuMGVMnvrc3vBcaYvcyT0TuM
L/zG/4ztYtZ/VnzawhYkofYCGchCgWnUr0sDUawh0hDQBBEBPFidYQbPwpgMvihH73vWF6U3ERDF
U8Mjcul7b4Y+S+IzABO9fBgjlPiEckjMZsSi9GCoZ5yRolQNEZVOK0QGU8M5hODPG5/I/hM6VSym
nnabzUwGUXsrQVaWWxo2AJLZ0E4U2TJ660ZS39XTRXol4auIltF90Aju82QIVak2lU8fGnHfewgf
e/yY0SR4jjQxjpNASYTyI8MYAQCdocsFEhC57qTHaVXR7htCM9byPfosr3zZJnheRymPQnMjBHH8
V/acEYue4wv75AjhmiNgzTKAnGKBNKxxIhfTeoUm0/O9gyRdMBhsWmTz4dl3DNWkfniNVMDvGYIf
ak9lyHk4UEBZx3p44NTQBq4k7Gx2degzhw2XisJZe4L5c8Bj4DY+QRAMJgwkyEmkrtAHR7O+9PvL
00EkAI9Q4mzsl6zsfHWvSysra0UeICazV1SaihLqRoHw42/CIakiYq9Oc8hOQ2V7RUgn9pXp1oOl
4nkhyMYjDKmeb+5l714PhOuLocDwASbPdR9XHhMa3TK430AP8juU1h+9SrNvlqRqxXNqs/Nf8Joq
Pmv3lC1MQOTY3NBtn29ebuTt2jHtRWEAF93eB0P/IpOpW0cPpCqQSXsyx1ZuDo9ENhF3EgOCkCm6
5JYnRJ3fRu7t8Dx8AnXRzxSc1B0yQD+prxO/aAH03tp0esd37QNj1UWRMsT7LWOZDA7R5dEWk8SW
UOOsiGeKh6vdkwcw5FXuh3fd23p16tvNt1JMXwRE0uzvt2kozkJnEZcYx6EHux9cMXNsbgSSQsxv
22Qb4pu7LRpkTDqXJXNo4fs/jjZK47wesEPjcZOPhPqCj5h05JJlNkvjvsXk1owC2zChp2mRdIjq
l7y7YSGZKvPmp+dMYP2r3/xvm4PfAw73jt8rXzx915TXSB/HJaw9bUdwBlqFJTaiQgx8nHgHeKfE
zDOPD3ADCACmqPajcfGYuWJRHW4vP+LvdRVze2ePOncvgXfqcpx/oyhN9txVF+Nn3LaFu8eIxktD
1XAuScDhT0JIEOKZQ8GWYf1eFchDZ4B4wbpwKPRn5zX8r16YVYTZ7TIB/T8snUrI6LtAtDczsVNE
RRCgZEY2piLT8feZ4oW7W/eEPSDGaXexcbnAK3Nw36lgHwsjc00icXXgs4MInCbMN/Tdfq6NW5Zq
X41oDtrCLid6FGWxqOTw8T7zBaEEdDlnteBdoSdIPIAmlleMJ+SqV3HD1Nftn2bpKQxdRqBj5UZ7
hYtxwDrq9nEfct/lJ0GXopWraOQ1nT80OXgTwKu0AtmI8EYkYGVbAFlcgR4eg/6QP2lLmXsIcuEf
8tVo5HZGRVnDZ1gWSb8bZZ6w7FyMeskLq4rY1vkmcOFGSt7GOUi4yOD/NGTdNDIr0Dy9esVvpBLz
RKze5f3OjQTfyLGnsj34NVHfOs4PQA8euQPpkAuPbp9DYQcnnGMWMOIOAHAgFGDPT7jwAH/z451S
W78vtbBYdFEV4sO1fBg+p8Q67GrhpeUxGah9brfgMu4euTyVTObwy2vfyKx3Ke4BVQO7Ss+ahOjU
Zi47+1TJRElg/P5E3sYJCy2goBYGUK1PNtVMyIg+x5+ZvrgFQP9Lt07ecO6VDpz+dCTsP4qxEb1+
uhUCO7QH7C1gCkyTgRxn8YAuFtG9o9Iy5tTZlyiQt2tLBhu/StBuAC3qalg8VfJw8NKjAK3ZPSBr
Izls1BJsISCAUOTfuox83tcKIaMdTPuqzSeFla6v/JBlKXGMsT8AaPmNx4eVUgcED+OPjELdPhZZ
IDS6j+dJNvuZdvryCTKiPrC0hbqj/3o8mFnVGmJXyo/Rx1trQsXeV8VUDV+COX12O1c32jYJb11Z
PThhe0G3jvxNNPn7xoydVetYQLzAjRrwba6PKd97ou5AJ7k2EppxWDS809fh1QeqMxvvSJcTkOy3
HHsOG+xMyOtr6FS0P/xH83LyvNYC9+Gt7OdXjdys1NvyhWLuHNEJS+UzLBPmggNuXE49o3IR4oFm
TpCAOqF/MIg9pAxR9LZ+yADKec6LnWObCMgCca1UFDdfYGqjBRnZNyVuP8pS/LmfpPFCZkCR/7K6
PACuZC7hZH8D4q9FsNFQ2BtKvRhPCuPU2FlWuWBfv+sfU9yeyTm+c9rrLWw0EL+h6wjyOSaQYbf3
FWDCfSl+kkYklfX9sc9zvAH1/MtH73tj4MRpmjBAliHCeztqCJ20hJkBx6QmTbvBwYNxTGU8Va8r
/793Jv4NFrAmYssJ30fcTAhBZIxKwaobag2P3Zq9aaXGC/UsgDVIUq/Vn0slJYb8sm2jvyZvgTaW
QHgSejFRWCjnaMHyec4q0stXQRUtDyhIVO1KiRbtMmysITmwAHYcxGKMTcNpA8e/2wMuSJXOOox6
PERmlXu0xfkvzlZCMzVoDozhez/reWxEL6kWUKB7F/Hh0rGdod3gCLEbw6GwZNkfsxQg+hbv+8O8
tcBOyGxNSK+FsY6wSMTm2361/zNhDZ+kN9nIPWIyC36nj/kBXtb14tELeCxWwcniTM/vjZNZQH9g
HfqA6ZaSfcGafKTukQ9GCXeS6LpMxghcWy16C7YEXri3JobDzA6xc61SHTzW9AjtlgJY1GgjRAGv
3aZTU8pNmGSmpb5nJtfCmvjfUNqXA0RAQ25Mooen0oPNdOrtGOy/s8tcpiyFj4VhH6OXcMZC4V1+
xua4/VsVjEE6EeTwLVCOTK4kha1qdssFNdHcfIk0ScQoaNJ2Z8OuGg+KIPg7rRkOpM0moGS4btKt
1p2rzv2zkwBrfXyOl+2NSqjO57O5jpY8NZU2VRpYlLymCskJOiNgMoDVeiMhayGWeFvZN1opYJn9
s1UIMpAXOMlgEAoZaMr+U+IdXdhWf+/7IEF1gX+9Ml6bWLzz2ZXvEQlDuwC9xjm/o3ph2rd1QG/O
QXGFjHdXXwecGBshh3dqzEbonEDK0L7+Ubxk70iPIk7xtXaLRfP4vQCgYEo/ZBww6F5XhqwQQ9F5
q9nh+mIf9dObRZ/t2eIVq/d64gnHUpCk4DywxEbhuyIbgXxcu29pLjkaWgN5Ebsmketw6v40vgAV
7tAzdnK3itkoC35cLNJK1m1dXXsZYE9C7eagKjtMVPy5PTJHqIz9ABZkB6xe1Qv7akgwFSRYWon+
Tofju97wDYZnoEBcgTcYXSlSNE/yuGUZd8keZMHAcpE0ML3VD9SJB9IoccUMHOuRqWZXgqn1dE2R
e9NszppLeMvAXzleqRP9+h+WUK+7T4444NyXrEKtyr5EWt20rsGHcMc7PJKY9vcnCschzi3JoYRO
m8pSFgQZ+npAaxUZ5ct8KnGxxADdYF3aTL7wThmqFJfMffmwSawbpD5509jn5t0Pzr49e86fEPer
enK9S33VqN/ZG05NuPlRLD12cjgvOJfc2XA7Utpb7K29mrwoq1l7Rxsq8nVfYQ5XFJ+1iU5Ay5C/
1bTCc6hbHS1wlTLQETyGGbv2YXU3Esg0AClKalK5jS8neLA+RK1Mk9GY6x/0U+VVnpRSmoI6ndJR
k+l/UhXDKHlBixsOku6CRQ66LtofIJpVLxnAyyMAcTeUgL/YwfpyXNhes+F0l9SloRF5fgM147yU
f5m39Fjnu25sgfYkIToPQ8zrsKOQ5ShiGpWITg2isiAP1wPy21BhffBR/jTyQmFgP0Zo1rOlyNEG
JoT2OpekzVENg0Co3DSaurgC9etFvOLB6ipPuEt+w6orJsAW7rKln0+y8D77a76XnYj+ztXn0xOD
oK/uKnRqvuTn+GA9PEsgHataAK7RPjZt0O3taqeKxb0FbEXioexCjqeaaXtGgkkGiC1uwOWtkHFI
+4GuLhI/nqkIpQVYL6Zo0tw5W1fGsQ1WBz6XHnu3PhnTy89fiUaQJEuaYntNddAqKKM+GrZxYfXf
OEdoKQgtSfNXgAxGlOEurTz3T17xc36UoiPpkq82LNGZho4D37jh1z/htSQazndOTzoQF14vVHGB
OX5oE5gYDXUgnOowJ9kXamasJHv+8a95tvdp3QOJeE/V/bE7BzH0HJ9C/Jf2A309r4EuLdvzUieH
TrNyj0AouZ9RUIr0h7vMBeitUyQ0hiemG8Bf6n6ujNxnoey8eobHNgMM+OZCT83uyxnrrkb73SCi
ffNE3cMHxHl/BRkuq+frwfAKft0DCopLk0/D3g4RUdlDPZAHiWUumMPl7P7mZ5dq3Ajwzc8bp5AN
NhVbjPyY/l9yC8RO6xsCiCMMVn69iI/1+sKv38SjHaqaRMho0UJ8CVl/ZQeZWuEaCWTR0fPDv1uQ
5SflE1BshPZtrrZcTJ+xf6ypiaFIgZBRftf01O/OeVt0cx2kzq+NZlN05HE1zR9lhBTZ6vIq93wU
HMpoa6bWyoG/EJJ+hFdtSkprdyPRhSh6t2XrSs5YDEMhJUJ5oJd9/fCmyF8vey/XZ0/fNQ+vqRjp
zMEg1sWFKBEtfdPNCwdUebfD9Vzr0c6uoucShZ1ioXMZdwXDQ1ZfqiuhvM8BStXwa+L1L8YWQxbU
WFBATAE3HB8OTMddUuy/fQ4HHErCuSVyjnwdy7x8mvkAjJzpzba7wz1nQQnFP3AyLCIqpiilyUUF
AShcJDnjdwVB2MJQqzIGjfUaLFouKo+eBaz5twlcmPWaBDMOZvwWPmK0uCv208en4ZPyKooDzIha
pIZ50IwwsnPX51De1kgl6y5zumDUZLcJoogeSRz8EHkkfEeIE9ZdpEVpkfKkzf5WZKf3X/WTgUZr
d9iGyDuEmntdOqIv1yWN7ELIiApnUvz5VrUQ/snHFzI+QTREK8Jt8E1+xQMAg6PLMzFzykkije4i
VSsuSDpQmBX2g38KfPH8hWZsU9n0cIBhyu0FibbYn6ZMNfkBIOFG4wsnExWYGXPLEGmQEZl+d5WF
P8rYuah1s4aVIJhhXcW+vjijy7kHDjz3ib20hb5DKXXtU8apDEcbs6rl9lT7VVQzumlkew5SOIVX
Cj1iXpaOVJy0AfSUJ+ISygWc6S7l76WLlF7oVONPteYcGy/ZLd00/5MpxwJenMy5IQY2m6f0jklh
VdECeyDaCPLaf/TSfDWeVutHNbboev9TFkTQbM0wAuYILLIjF5CzoAwwvHnhkanLABk1ZaBXN1dJ
0A4+vxaey9x1yF+70+KK9aSQV9i4Hlpk4voojaakyNrShgpsd+m/l1DbVZJYbd7T7Pg224bhBbY4
OPTPqaODAYoCAhaP4tMTNiuwwRmF9Tkk8KRrfa3BeRhFMGqr+N3j6w1RsoJ3ep3SM1fQCTLDq5iT
bfzS9MN5i9RJAgeJBbiFPaaRp+6tP21NkevDhI5iKEWG8ApaTfRJtfXq/toDS7DYpAuHageOlYXJ
j8JaEcUAOYa36XdYBPcHWejT2IBuTFozPC139g17po8Nz9JUcuIEaFTE2ZeRo3bVHNgfuawLuN7W
ZZ1dwIzsNyurcv5i7q+LkrNFoH9EPNdySFTwKM9xeAtKFG+Iw6kGz4dMYejmAU1RuaaJgo4tq1nk
xuraXvZ9aH6b7ISdcLLerIhEvCpJstFEeIv2GFRGzDBpL2d0kOvrGhYYamZ6ihr8NjvXHxnkYNSF
cL5MX19Weue0rvmxFu66DxQ6y9NcL13P6wWWX7likeCnO5P3Y3INNYUw+iOJqoZjP1Qmvs5C/4ZS
A/PgtZnDd3o3GfzZqpkBX1+bFTCVK2ycLcmYXE2qIUG82WBDRFUkOp9pRxAIubABD+jGbmVW38cb
b9f236n0GHnZm8x6cQwAo8bX2v5RULVEPHEjNisAwnci9JsQR7t+eAhgTlg3hAbtrJcDE3LBXb8B
7SPzbRNBn06d6OZcvBfv3oGFEhIzzjeccE6m4Tk6RaoI8Fr/Y4cb1tpsuHRihiDP5IiieSpS0p8Q
MV50GVLcRLJ3b65u+r40U4X1o3rwFKjsD40kOY7K6nQmeMA1ka9x5DMdkhPvtnz9eM6zLiMW9XpY
VaSW6Y9kzuSua1Nfxv5v2v9DNsbOZHJNVbRQ9MCp0XXulpIleXWRdOXSmjQqdH3JlRY4Rj3rQoPV
AJvFfN7upAm051aP5S3g4eCgkAnPIKHu3EoOZQ0mqjQI+a88dr3P4XvU3rp5UecqmJniLwPxlJDj
39XL6bAaAemXUThswiE2rEHqQK30EvaIhwwI7S7Dgu1WIbNKAh9N0/DlUBEwVZqrizJLgBvqjKt8
aZ9OlbvVb5BMujmh1vowgMoeUx5bQtb14LCyTXYSIAHBHrC2d3EPZU+ii1ByWqPli3XTPmaqVCqP
zuzTHFAZPONJZRGJJ4r7Qivoyi1TZLkXqGRsLUDNdl2Wqogcd69pSpeS/Y1q7u8KxDjPVr+BHV9X
4QgM0KeO+o5RWdoFaIRLham7WY1zYTgzepjTUToQ6bIXy244ES9cT/KVnc6awPCUp7DVEIG4gA7X
FPPvPqWAFUwmU47Q0Tn/ewMChVYIGUiJoxkuv9QNajF/rp1j7/fzft26N5gCddzvEmgrAWt7miZe
gmnWHFJJmcZyUd69673UXQyY+LUG9KFll4cTnumZkiMoO2bPcN6D0To3niE2EYpobsX7bL3kah+p
VXD1VHkjO3YlingIQ/C19Xsr1q9JTtKhVbtlQS4PBM/Nvuk/CwOx1V7gm6PaZO537q/fHaNFoJmh
9UHW1cZgVYkGe10cNmrWH0w3Ykdh8ZlJ72erZsWLiIsS506IuSZayMYY+lMjsO92WiKdOGaJ9kqa
2UpQNJaQrURlB8JgkLudw2ALqyet6x+L7VzS00ne9nxzY6oQSRXmoQQJJvQg4vRKWLBZk4ypk751
92BnTMHYWB9gB/a5OO/i18ZGF31jBOvTP4extjvpUZ2lmU0wtKJA0ecU5G9ZHQNl+kEwfVYnF07R
7jl6NBjX14uQujnC0oGJvU0jqPX1pOluAevnFx2FxquMfcyUUqrTvH1sEfBT8iTfnrzNsPkbLHLX
i2Zx96Zo6jQSDlYgOktjvhlYyPoRtdIopzJ39jReOt+qwKbevx0/Do3cpPX/FKgr/wuEeEOpBvmE
/C/NCjqPTMhPPm8bJsP3zTWbjvT3Q/8Ik5ubXAtjA9Lz+CsBLilsoLC+kxFxXi4IhHWtA79hFFZI
3JIOAftmqsUcRZkKRVx4VzwAqmejqcA0OBHs/l4Tdlzdj62Zg0+GNJBNN7VifTzB25yc3AwaiRNb
otT/80rtZWA9NVpN0252kyAenD4JpvJSRthHvi0VkGPPS29qE/IJT3w3tqpv7AFSEP14gXEfCV7w
KUYimyuax3PTUdh0iHULABFSd28ValxC0QtYiXA6tVxwJkdcGsozBlSNT0H0EO8ytn+/ebY/8Aq+
wD0liELEwLmN4EPMImM9npX4/ElJenNBofexx7xbAR0uKCd7un1/WjD40vuWyfN2v/qlMz4cpo+m
6BqRjm3gsZFfF9Po/tzsbjaE1IAF/zKsl1SI4rVKn70Mpxboj/wIhhmi1J6lyk6VWOJ9cp2MMOOI
M6EJZdly2UXyYJVUPrVfIZy2FSTRaTguQGOpF741zu73aMjTsUDxlUOdJJKvs3TEbwSJ+fJw4pvl
MtOruSDA/lQi37buIACbZbf3EeyxgiYTkQsZPDkfVWTVGqXIMWng3m/ZxiOsL/gi0pPGb+LVxdBM
N1+jecakSZPJwfFmxhW2g/0VdoeYFkXxmvL4DfDgyX33cDq/GOLZBHVBUb9Du9xds5IXlmeWNIlK
E8CbiouMNbSOczJquZBpLfcLarkef2jNqIUJUjuoynXVljzV2cWoyA9wRjN56Wz9dMLzEkNlWhSC
bU9jJelMVj/ta+oxEevkDqjeAkPXBBIMumGlCP7ermdGkQeu57f+XV6zaa9KWthy6llxwUnwCgAi
b47+byhNeJhkp5AGj9QYdCu9vGJ4wNcSIaGJqko7yHjyxWg7ieRRn1GsLitq8a0BdrM1wJUkTkWf
3rGRvy8ql0A3YKILC1c2cgMG5QVXc01AzCyW8Ace+KydSsCuiM7vtR3cx1nel3RgXgKXP8/HcfrW
LA5mhmRkO7rkXsrTkZ8YfC7+tOJlm7sBO0Ugq4H4HsFmb6cRKT1BlzkTjQglP6m6ZiKZO3wAiwK/
rpbNwcjlHBHJBwsjbPognswFUcQLmJkqqi3mx7TkBcpJFrXDVc+PW0I155JKti5MWEZhlVwF0/cG
c3kJp4xDD92O1srZdOaWXzmTT8c2OZ1ZY+LsX3UWZzo2Xmcbt1eJyYvJ42ryj/a5b3yj7yDPwAna
arkviAgxFvISYeyruaZsTZF3IdQy0qlKSE/mbDlF05N75YINUgs5ZNVHkeuQbKfxgamQiXbeE7++
OlpW9pEQ9dTj7Jdvh+Z3uwu5holsgd90MKmXB9Lo+PvwlcWkt32yjG5RajsFoFCosQ9/a3EnnyOR
ZxT9otZYLLLfvJ5FnoC8hTVZFSMXB+/OyQBuumkk5dcsGA7s9M6Ck4MXo3tOsKAVgTbZAe6StGFB
pwlXJ2N5Na38dhRLAwCmXjDUK85Bz/TWk844x7jSsJLlzRwf0dcdYo3SBoQfmuLsVgjYTa3x1nHW
VzQ3T6ebJs+roGVU/7jsvD/DHHKXHR5yekquBLbLiLBGLggiexyOfRlpt84DroQJpMt7FX1yD5VO
20psSi3KlkXzmMir3uO0i/gZOdSnbXp2WZZjyD6tGjtfEuuwQewaE0HhujfaHM4RSPX62ouwk09Z
FyZoqWUmd/p4h8Dx9iH1rwi9HQ/74peLOeNLUx5ygzuAROZvK1tqYfEiy/XSn+oIc/MikLuuBeoo
dY7khmYieB985iAUaP79qNWRyp1fVRJvSmLdzmBurUBQ5U6c6i2mLLKmG5JfmjrgOWU9xv6Nmwa6
KVVyD6ketWw6gVo2pTyl50vH58yNeOh4leklBlDrZgnlqFIDm+LC1hL3JElxevnpyz8cQq6bze2X
cGlEk4VufaROzrMXItWCIVN651Kcr8KHa32Wxzoz7imj9Wr9AS8VyxL0QeMxE/G6BSuS7b8iwLJ1
5F6eOKSVCvYVVywJjngyPmS78urq6HRXGhkDX7huZsQrishYEi9HzF988EpEZDVWiV08xv40z9GL
XRV2GxyQyb08oayej1e/EhWSn6fOQPujctWycCyXfm55HWCDju9nsFym+TN4bHnq6PzaeovDyl00
WxTPGsmuJ80HwUd8dU43QJHqVYf458KtrOPEO5RyypkYba5tWRWbvwYrqIOU1n59Jrc+S/JxpRvN
I3sdbfZ79sVbsdj1UbkanFnkPvhVEDJsb2HrW9eqsGSYJNRHfz97xwn/Oxva19KqrOOXvRcuo2uU
azPk4vxUUIOL/Q/BWmLiV60hBmeQpPwIqmmcWoLWsJsALSV1A3SkMEeqlrzVipf+2EPZ6EghV4ol
bXmTO4RvvRp2BsTkG5UB+ob4pr+4Xy6sH5Cen1fucy0YmSKhTNSLB9f4y8tFXUvGXBBKPpc/IlMq
VnA8CFm3M+JJ8z38k6Iixvz18RJQ7b8JAmndNbPqetjMhSdW4ZuO5h+egjVXPhvtEWZkmjJ5a6qZ
G2A9THu5oNQhaiN9kmCbcfNVPyKgisPjSfy3hIHT42ta71SyaClOdn+dCuHUNcpM0LwbzodK0AJU
JER/RC5sRIFSu9MyxK7Pj28gbgfzU95uMFCQ4WbZt7QmH4bI9Tld2Nrw4VJA6q00nrYaJkc4Tffx
phwyfPFRPjAOa4MaMn9eWV+tPO8C/CjIiJP2DQ3dNcOKYuThS58KU4SGqzQkOEatLqYecV3/oY42
DlgcvZzHlE6qSt+XAOmAxTK2k4D1dnhC1vTyprj8dExj4JQpclixQg7tKzsveqN9ISi3dNHyslh5
/Pqh4oCGJFzfIHdF+HkPdKothXk9xEuhqvV3rTuTot+bDC9LDT19n1gShxS+m+rXId36O7cSTtZi
n2o9sy+GdGZeTcX2f0oULhUehUGDSw5rPctp/KUkfz+aXcIEJyVxu1Kj5Kb/KZ0/9eCLrwVvUXNp
GBlB5TY85h/Ot8CZtxbPg/1y1D/MRAHIV8DmKzRrLekBnyOHh8zfGfLk2zHNx2vXWI5Kt7f8xSS3
GDegch4YY+rTaS1sWY2jg+srMRAUZegwqW1M0gKFJElBnZmE1V7KitFll0KynlfPjRKYBLe0yFMP
YGbkX0U38zCfMvjI1pKDsBcJ7hTkGpjpQTCvTJ8QzJ4Qs2Dv0HuxxW3uwWeAml/PrP/VbAnvGKYS
N/sWOSlDbEJZ3hb7hud0w8U9Vzfld+x+JBZENQ2fpesheuloIiceC5Zj8Mh2uhZiSzouCkjp3aPO
xFN9V3qkGIQKSx1lmiXhbM/bX++twI5SOssU/aXDe4gu8pPUZxmSkp6L+e9GiYKRbW9VM0rtDeNh
bfNtMcYEiukWZmBwP388EGHZXkcAbJ1uZEkvNZjGaw4HuvpK3I9Sz7xpFOy28o74QWIKCcqa5oGK
A35zf838kvb6cIevFn3dK+jE0s+ZHBfXyY+ygSTReFtHMOD4kQB4WAxoMg6FNnFZDxGEG0Q41urH
qA1TKivQL9sWNVsBRnJujc86U1eNGBhKCUDFeHZCJVQdZb+Yx5ZqRCNP8gJMekF4Wo5NfcguiEJz
EIc5zJUZF4bI/uUQxXSJw6ji6tcXpWAaJldmYsHOdq8yBYiumzsLCg84GORdQcxLRRToM05fGQQM
Fh7wvIvwDpm3aHx2hbAFEOzWPe6l0G6+i/skFkGDSgwA9jEatuDn97wDri0eLOF6HsDjtdD9O0rU
USsEfDhYuUj2hYvf7QCFZ2WB2DN3XhvRCcv+lIY3hUOjmqI3GAICPBvdoBeIjRopiNTp8sa2PAfn
r+uTCxOZZ49IZ0T2hQSeQBf60Fkp+88CThG7EFIpAVYL08J7Fa2m0oGWndzCDoD+WcFaxG/Oi5Fm
zaPSJVoBqqwEwNmAtu5lPwbv+wxkE1wVh9YzaLn4eLAJp/Jb0tGJcH2nAKBLkSSZ5FpL1HbdkBvD
H+SpDtCvjpKsDjO5dhGKdTcoDYKd2kOt3MFjUJckeI/x13z/XB4tYWyrfsyVPwrpPWoBZXHzSWMH
RahPX6s1kblClzQO+cTvYfxw5h1jE+kM9L4K8Kp3sbe/CSGNFJvCXI8MHA/O6+7uOAwTO9UQ700O
vtpVifn5PZ+2ZKM0BQ1s67DvbsV7uLJrtMgHGkkTfHhDBbgMh2nx3l3fMynR6yLojiOUEAocWs9J
/ir2UJVcUrMUOIT426fWsbF73d3s6zQ8nyc0aQXdmMkTImGo8DX9dN68qUn0fBMF8LApnl+lFTOv
Xp4Fzcd90mOb0Pet9+9BbXxjTW9CxMesHZ3Irl2WPOaZYmAuw0iEF4F99MVIsqm62b292wg3RDqn
fCIpOmRmJhzOkVZEVftohsFt3HgsPsJOEmll6VxZNAEf23pUjW5upXCYkph2CUJ/Ks3PnrkkkL2v
qhJHdRywclaktTbGNa/tapKE0PJ8IZhZLwi3HjCJIgiS+KoCvAyRpzv1Fe9Mb5pPwJUnM0rFMP6s
p02LFWn4BiFCH3zf6eMgcd94PUWgzXqk2YzTOyt4A9S36rbru6JJr4sNkQKiOfmenovaPkqEuN+k
iVB/7ekoNajfC8e9G62viXcu+5POZdrV+UXczf0utkb3QR9J6NMsevVkfffqKk1AAfTqzH4Bh4n6
qvmCnbNYDIztJz93ZKGg0jpGYo2M9wabsZxobDFjd5Y1hIJLy26f6iaTCIULklc0T0qnfpePQzsp
Hjz/WrwepqsPxxqQOPnRAy0EMrBsnPcivr4PGpi302iOQiNO1KI1iYGz09oNMQDe4qhoizO7Yvvu
20HDZHSgI9perrNg3TaT6eTr1VRTY4uas6azM3gq5bG3KJRe0XlFkwdKVbX7D+S4vnjocLQElywJ
Tz7l4QWYQPY65WCka17/Rc8gFYdPjTP2DKKaBqiOS0j3hVpmIqdLohv96ZTBx1TgV68BJw/nvF5p
NZwdIS5iYeScZX1nLTn9WQ9pN5LCMNw0kGJY5Xft6VC1/3N299/ZSXfKTbahpOJPs6gqF+z1A7Gu
Z4YC55mv+087xOdFIkZa93NJ/VTuFlCNff88THaHbkc/njDZrEPSQwO3bbrekeb+1xzK5Oh+SfI6
SkWRucSeIn0rxxUrOOPm0L43aVf05c0qthNoHvUIAUCUxbXY0/qPYVWUjuCan33vyISLsyUbJMag
QUTRB3rhjR4pT63WZ+SB2GlEfw8JWOKecIzGeKrFo/GnR+XSFCbrzVkXI3qmYg9vEDdKWZPmgFT3
I4CkyFxaE3Kui9Do81EEwovwI1VW26LseZmWvG+DZimuyMJ5/XW6a2Lr7zuhgSTWAduv2+EMyMlz
7zjP+JPbMbFEiIceGEwkHNGN/+3ETfehhC9o7ymwaz0HL78iwRvkE8Kz68P1pFVDPeobS7ann5Ck
V9lD1l25hWvlzjCKSMX8PQ5PwvXQnZYm+zFZl2tHY5HrOGnlzfiSH3A+nzvuFG0B6+K5Qh06geZh
rjWqxOra9RsqOUcPzdlveOxca/S3GjLDntI6iM8Etr2MRmcYAPXsQAcni3tYR1PUPiWy4pTBqgQj
uj1nlGYkUdaMCJmSjKD8YI84zIvpuOW6LjAAz7+WBSlHn0r0yDvLdf/C2UEaWKNcQnxDi7IL14dR
jyc1rSZKVfuDrNksRe/8y25aiIyL0L8bxCQA5oKc5p9qroEmoF72TLXwrmL6f/7eBu0GbVw3P1TB
0gQrBkzBxsN38o/m5k7VQIANh+MGWI+CRAB6+O4/y1SrcVcdrJ+MF7V3XkDs3jhqpyhmya6N4LuR
XGnlxfqp9xz69BQChuixlpmR9WEyvQ4g+ThItEjH7rN7kWhbcoYxkD5BbU6R8zo/nK2YdWDTXoox
6oFPk1ohRaNFMn9FdJTkSVWczvbPC+dDlZOpXL/uEl29AZCb0spTHTZnm26C/IBsmqvEFtrJoGuV
GSYsfHDlDkBNC2444m9tIR8Iia5hhWg2VMkXYgFcMcE/yM0rS40YUCRsP6byeYt157p0FHlsdVJJ
nIusxzKdiiVDbF3rDIQ3Z2UDIfMFPI+sIeoWjojNedfWUxJ/Vj4Y54BrEzDDJcB6TBdxkdj5wwzt
kRQN40CV9uKKzT+rNQli6wh1jhx5kLWYW2pNmpGqn90tGPZhKFF/eI7G7lrqkPLRXHrR97DDZNq4
7agARc0Cj9mAji4VjyHyhqhu852nCSpXffkYHOZYIYkNw9Qnp74qJ2ZVPw8ean7vdlINB0/Bulsy
5pOv1w+28W8efkI7+yLc4BNHEDAvN/n44CYdPG5p6y/mQvoAz2sQV297qzVdhiVpe2a23/JUWMnB
AsmMnk2HIfTIxyn4AQIZcMK/EYoS3BFT0oVdWouOb6HHd10p5a95CXzbq/CcErI09slyBh5wrgXR
3Pck8U6lsdwaAI+mfsxCzXqklx20jJUwQ0jKYHQkCCycpgDXTt57yNb0D81maNwokQtn0DCsY7B/
r0ZhhEiYNIautNh6SLYZ/h50UX+8aEh740DHZcINNBtgrfbL/cQTAToUIPgdLQljYhcVTihxatPq
tvJXAWIJQU9Fpuhi145d9tigT+0vkPlPt0PuqsSkW9ZkrrKXuVHHnxKzt62LC+QmTKCnwF69+8mb
DIaCzebM07MAwax6+/FPZNVkn/o2ojw7Ce6iVgGQE/mD9j6GSW0JxrndDzb82/TcR9HCCMLZaPOI
Dh1ZXcE9NJJmL9/37Cej6wg6L91Gf3CxUcGdOU9Sj2en3f9R9SIGkSdlLW1BTMY89ZSKfQK2nTR3
Y+CpH3xPYs5QXz/HOl+aRbquvzI/uoYefvxRld6AKKZEbV1qS2HbcIFzm50iXdTLGJMo/iiESCQS
zKkFcp+/3cY5jpDguradzznGKTB4uitUo3ugREKQHkXfVwyEqSq78s6C7VpcUlVOZ7TUyqvKM6Es
DVUeMI0CCDYWh81wMIEl/stAfFfddi+swp9ZGW8uQFMfU+7z6duIDxoGgmihOLf/XRChF3wqgwzV
RxQRTtUJscR6Oke67blVgEY/VfqV1DrJ5ELHczjf+AXUIVAJw9nz4K7DxV8xDhynHVoqPGujzOQ/
f8+pfgnQASsQiojJM6cUo0j76x2N2t8FmpvTQs6oaFxpm4X6Kk7JiXeOa7doipzTbpYGOLX9zYQb
D5Fz5DinNULIoxce7Mx8ei1SXSSgUzuoSxSS2IoSL0EWc1HG5RnAWhB/Xq9KzUKUrEhzn1Rv7Qaa
/VWxBwnenr5OI4DVOgloLqJjSKajftLcNjwhmYfTFzdWMEF2k+rxg01IqQA/uJkNt66hmolwhUs6
j005KjmyiYjGfTh8U1jvX4TUn2s6ZdyEAZ23nidzDHdxtDL4VYaqoyCSMczOjfvtOgnlMsyWA/NJ
K+xU8L2zOcqY+RRcNH+G2WVfbrvWooHc/wGjZB9hexoOgkdt8U+KfGoCruMzrCqVUTjJRMLnKbU6
oG/AsodbxvJWgBXkU9Wt2GQ/VPHKUivWDyOCKC4jFGTw09w69TZcQOAPtgjnYeU5ak1ojce2jHZf
f5Ad8aYFQMCb7Ed8ae0sOyURhNzjaMonnQv22J2gyASQHcpSnquLfxJbO/xecBxcvKFGCwrby1sh
F/9q6y5IKMbdT/LAWJ56Ue3xW50GlNV5tjorrdJWXcbgZ5vU9hzJL1OpBuGqwewn76YPY9YVKX6t
FJyqcIGLJ06D1BeGvdn/DekMNqJ/JlkMz7jpSARchXwyhqKhjO3BY1DxdO5DkTF89njUK/mlCH9e
5IBrRVcvNy++4kAQ8vIk5NJO2sxRcLmGze943sSIrigVti7MHp92wZ+AZAk63K0poQUBURRp9JDy
gHbdiROcfnHuxBTUvc4iDss0sJL6ykY5z5UfCQFx8PCsAi+R1M/1eTKO2HUGDyv7Fq24lcrmMqSO
Wsoffxpl0T0mlhf7un32e43xSCCt2X5x4qEFHMcAw2oRBj0dN53b0aDIrPhijNkBcbsfPWpctUHC
XgrKohAOLzUbJVdGd92sMfX+mMNeGEXgG3MlfaN6l+PEksY+OViTf5vy3G3WLVI/QrkirivfbTDO
BGebiVhrL26mDdjTgci85BBqsUjorzxuKvdoiBSufxAotR+vqipol5BOkyqzsDR+K7/N/si0TBs6
L+EMfOseo7W3xs3NJPMGQ9LUafGbhJdqRlbxpWVm1v2+VZd9oaAKuAHWFhlJfGo6+WGJPCWpGDfi
fT3Jp49b2JK27CpA35ozzrLvSedgyHvbVoEKAGdmfvUHPv79TFgMKxnbi3LeDYg6zmaWkoyLDk7U
eWU9oBRjxioCRpCjcpx9qAOoR+iBFaBSMjgRJeoD8O+tCbyyZ7aZfOQqM9rSoX2jEe3udKzwVH0S
tGJD5CUEUvBUh0v6BbLmC3FJClRTyPoAUoVNzx87U5EH9jOZstwlCPpNDiWsO1h+2LoRsMyzgdYk
Gvzfg1ms9dYIC6UVzbdjPyAb/SdohBdErkNbj0fwr94bFXiHj6spREMbxOMo8QFzhaHZAgN9i1Sv
nGX/bzDam5Fngz8ZmhR1HtfYN+71zXhw+xaiwxp9NEoC8qMctNCW3ndZ8xV229r4bFE+YdFS/Ldz
UPmN2yOhA0qJSq2IRKUhZFillCW+d+LwV0UzpvqeDyCCwehOGafGwLiuvWSVt4an9EplLn0tkOEx
6hWg8mQU0u+J8CI1QzEnoyWhIPULo0kFffIp289Z88N+gzmYIffSj1KscsDNyzM0We+VkVZQuIlK
DiltvOFIFz84jzxoOEBUIMM1CytYXWjS0uy5i9Lus2QjudmEGNkQlybdjgpFdcF2ykQl2fY5bIPJ
SFwuuBRzelxn2w0nG47p5eZwxaQRFb/r81Ftjq/BEj8p9AgDOLmEc473Ke2m4b8rrdKgYmRQaon0
HmbdWB4YU3nKI66XoOg0z/QiIHZRXhbKKYdlLJewuXYytRZ6xM2pVkKxrOEO8iZmW0/Vi4kEYvGB
QanCEPntgGFuKDjZF0sXa9LjPIof4WFCADARK98D1DgG6P6ychJPtj7xDxwqXsr9o4nxkWTSBKW3
dezcilNUgdCx1zrrVhGZEjlQAtb6grR1XwYlKIGLdiR2azCbpQtmSjCBOdTQcpBJfQqVx7rKiR5+
y0/R2QutF+bybPsXw9187qtizV6hd0O3fk4o3TbEdga7pusjs19OYdUMStYjRh+PR/QPaMRU/uTf
Y5tvai73ELoQyjjg7H0/EfJHjUkdWoyoYBz0bTPiQm2P5I8xSiJy0Sen5VqalYwCwPcir+6w9pJ+
xp75zLS9x4JlcjayP7T1vUbShDWncgk10fqhfjCyCErLe5bHvmF16lOx5MvkdjUdn5CRasnKypI3
vvz3xe4tzOQBoX5qyPhq6dYRZFheZf8iAeTfPe76ryXiIwXOgqzVBFYkxJlof60WkyGIPM3BtQ+f
GWP1Jk00COZ3ajLw23ddTikqC10fnAn7TWNF8uCpFn7BLNM33BOWYtiN8LR6C8dlk39pvfjihKtf
YvZYYEoOy73iolYZpZSSJ+xfkEOgvOq+6LL+qRa7Jc/hbzmTWhMtsGWdhFIlXT9D6e8G/BiX7Fcf
W1ZROAc1ST+d+MTZBjAuXDZLAHlQ32Tc0j7hUttuAknVVpzn6CXVyKtrWb28t2264rDzKmQv6XP/
gw8VsT7ZhNjS39sL4ctsof9C7bNVnQ8x8+Q2CtvuEuynX5yhLayKVDcmrj2M9tO38uAvKsSS9W7t
+7CNgjjX9/AyxDkyVrobIqYI1IE1CxRAGn8D4DlU8K8ZjfJ4U4DgItuuCOy0rWxfG0PM3XjNWyPk
yM+k1O6Wg69ySeEPuIXcHWUqdeuVSdDSpX9lydWPqqUL7HhQ2D0U12cLHGydPcEzjVPhJVo5W7QY
sOhdxMU8J9uvfthYkpCSEgRh7l78DQ2G5tced0gw/fmxwaNerpzYqdNmOphwN7ewo0sngh4bwFss
Cg0j5i6V5LOCVd7AxWBBdg2XTeCxnldWObesIy6sb8mOjMvgckmMNFXHTtMUv8goNASo/AoDuwTU
vWgTmBi7NcdUhe/dJoI27AZzzdq6F/ljdLWWb+wgUHwHGG/OpVLljSCXbjkNfRKQFE5LLIZHgMbv
jkgJtZpoic3hQrJZi9c/5lx6GLIK+B615ijZ9Ep6zs7QciubAkITxz4PP7f8B1fzTfhS7/XNhZ9+
AtwVjLBOJ5KF04887IJsw2rfTqU6okN9kecnsc2YARWxemGKA5e6T+e+RLFiacUkJPEN8zzKVXdp
dsnz9USbnCanLJVv40CNqeuU/GZqDhjl7Ajx/FNBrWTdzWQvlSoENrMWgKnVVS68Qb9XOxAWMSRs
hSOTUqZs8mWoGQwVe3xToFaYd8hm3uwH8ct6DOGPsZWRnA5Fzz3G5ofL4zeoI5CwbjMkq2Ifbxlr
jMyC3V3auv40+8JLpVYvH/xNH/L5e+OdGahn2VJH/6cuiWu9i4snF6BlL1AP84iB0G8vJafDN318
gyYD+LeM4HMe2BO5Mhlp/baJwx15HDKXA7AlshE3B/ZbeR+O36yuu37RYdmNLrjdWboGsVNxu4A9
k12nlqj2wwRrHTgpqSqmbu85KA36nKMYJ3RYzCrWo3ITNR/dbW/+rilMFFsGO4Zq8XBMkOT5tZF6
AKxWIjQ3DORD0KAcCQjF3L/ujxtFKFDIe6v58ddgwc8UIwfK9hcyuzsauFdXZvCWkf0/dnFLi6C7
8S8SrHMwRnHECJ6kwjYu747xlVK/i5fk6+91fbgzuBhkWuaPNUKTQ8IgcqftZkBVf6SC9s/699KJ
JWnxLnBoZ57MtOm0E+8dLLAsvzrgECBO8c55KnRGrFWnylPuc0DKSwgx6Gu+UH/BZlH1exxfWfIV
oWVla7XqD9eCsR0iMeSG1F09VNf1bu8M+fgLd7qf+lK/mX4GvIYS7Xkl2wY+63qQNR/h1Nn40fBU
2PWgQgD4+7mlqmqjcyH0hoeaXMD/PRmYPfTYjbQEQrKLP2RhNrIqkkfX8kLUjXw2ccrlXqQMuP5a
U4lf/DkOBPlxMHO33dfqu5VERgbdHis2ngHxxTJW8mIzFaC0X8O4thsoy1malmUUmRZB2LYgsMEP
x661nFUY/zSszVyt3Qny46UiQ3w80fSMJ6O6MUhYnGWraamCtUXUWpMWZj8U/1e8I2iISR4dRcc8
AeliggPm8cEQaSiSiUUS2Win3aR3wDTtGLGt+AsrJHrPOskpW7oYZQrDnaccYEGgDloF6tTBeKyW
jHHAPmBf2v0L9UbTo3AHwjB4tZXhNaK0ZD+WXGIYorE7BhqmGFzSVRTS9YJAyoUs5mY+6m8nDcZl
OCr+vGYfjYFtsqaDHcQMwDpDxIcGuzToqNPfRzW3zcoFsNey5C4yn0B3J3r/TR1/KnJewZZRkkUJ
ONNUaX3IRcS+iH90kyGrMryfKJCI5PkKu5lXdNMPfJ7PexTwJFeAkmdwpOzj/awrX96Xto1M3DKh
PzvCugD0LXzNfsesJs9yt3g3pr+nY1qdFfSdWIK0meuq88F3qct2LlwezyX6jwrSRnPic925dxQK
734WoLjosJxjnh8LIF6RCbTCkjYEyfGvcngpUYqLhrh98EhVqZTESFEnrylyfisWKcTMmkSszp4m
5ssFCiMT3drOXeRAzuCC2+AV6JlO8gRZOVqBDAF25PVhmevlWDwOvgCWBq9jo9hCo8KDpb6LfncF
pd+r7ncqPpTMAkDDT9M6m4UCeJj9uEBqLCkVRqiVZTKrIfcK8fvIHUJOBbctc4jX8/slFnDJSOts
iT+g5/TKngMoWE4Gog0xQycGop3q17t7P86xQb8Nt4/7IcZNY+jOBUEQZB0jboEtdjWjsZG8elw2
s9/Tjidk6NUBrU2ho4qIUkXy9axggxTCL+pU7c4cA5V+Q28ktvCq5nzN05BU2O6E+YAlodrDRSr6
8pvH/10B1CtdvZkpvHMkg6C7NLUEna1NTX/BxGz1pj7tFuXs+D6ECImRSeAQjPR8XwejUuzSTqIc
HQLfRsA7n9f1D1WaNW+ynRR8M8EHhF1I3qjUNC7iSaurs+KVKZ4EZ6VxUumITFhwPhieIHKfFNa3
ZFdiGENexI+QgQGAlwYuOd2oubau3/d/9y6CbB4K69eaXinfIfnoLpQAg8HX613ktd9Evjoa35lF
W3EwCVLqZK9GIjo2NsNgB8Wf8CHy/stwiATwNQ1/yihD7RyS0n/MscnnWQN/aHPOa/Rk/tqnIK8m
/KqhEDY56eQ25GdNHA81nIkUhNtB22iqYLu6EG4q/Q9PzKs1fTUrZnttDjDVF2K0DAwiEHq+tFYV
qHfHtk/DSBldBTxJpyeY1xZFe0k4FHV5R6KCvzLOP5lUTAJk9CSxmQdfK+jRYehPv0Gy/NZMzF2o
XcFEE9XAaCIvn7wVmubD+on+McjfN82rxdxv4glXsmxMLgajXxxnwiEde3aSJt3dedAaCL1rUcZI
0zX/Gaz3I9P9QrYC74W9b0AU7vOOaxgtIbD4zDLvdHS2fvhvV+uSl/2pHWALuLSJv8PMS7TbcZ8Y
7jbHhsa645JamoyBLObXEuc3Kt8FQ4CCV1zPMzxezsRUJJbAslDburECjei2YwkWKFyBGdZ8m3J4
7HU1hslu8omwU8Y/tOX6BMCCLrMtvn7HgKsbMWxMvdHJbvfCyqO6vgvso+D0QV50x4NLvQ1+Q2BF
oDzlM/NwO8jkp6+wuRXUDYDR2LBMGNK50FNrNwcfVjZaZ37lf/k4PlNCEyp3lHrAoQ1nFl9zw/Xc
PKNUEypbjaU7r7LrfjoJCgzMcDmtKpsP7rJy7weciEx53iVM7geqyQKJptVBrz057TsvkWK9MkPf
NCmp4ihJoNNzMERfHiz75JQ2oE3uSzycwDCaSj6gXt205aVkMvoBcqKNwylwc5OUoSFZTEAJCGmX
h5o5INAuRgntLp1pQJTk4u8S+AX04dZlGX2UQ0l0yYP+J3Dv+20uveZkJ4Av+3O5sC5TFkBZWvoF
aRg6IK5IQSoBS9BafAMfwvB8a4CndBsJgJkL0dEDDmEjFUYdAOM30Pc0JR4UNEC/R7WFdUepS+IN
Kk0dTIpiJI65eMuG/J8uCG7XvNfHWzAeL7jlsJHIOQuIg5ZUr3X80ftgFqcLQuTlaYRyofvD2/K1
e20YlJlACG2yqKupH8bitjFfYZTs4xK9lIxJw+bknGE1EW2UpPJtnzsHfMayfgwQlrmoJLKrflZ8
Nn33jOTNzkzXYXids+x+96+4eCRRTltxvQmDPIsyt4iPbeaEWTpMzIMr6JitcWvcWPm2tI62MnE3
/lJvY5O2inctzzJw/AsAwgEKI644VEzUnL7Bnxb3L+d63b9hhyA+tDaaYb1OrMQhZ5jcjPhlcEe9
yz2gHvj9dNIUfpytsm62bKTqi7CgwlCOXvxjV2SiSZaKk2ulx1QLObhnShCMhfhAxEJEgcwNsIf6
G1nUnnmBhRVHEu11T7oGq4+/rPSGkjMq3UWhlarIekr8JoBVjIG0CrO/dqwXqNmaGXalOQZRUY4E
+HYi7GW6zCXiNpSsTgI3doiUL/FgwGe/422SHj0rm17yoCLTxBCA0jTrm4WsMUY9pDjKzTaSKnrN
6PpUy9bUdggggBFhW5s6w4SszI2RR0IHZWQTkr77UBCd4vV1JVB87M/IvvztML7doZAZTFNgFpyo
neTv9/Ol9rOznjXMJ5nk9yZ/BFJWfCXVtKArmm93NOrYFf0NlxZEZjTZqIP9gyJZDxqCWkR8zmnl
/MRoAgcA/IBn1JV2qCOsPABVQGw1lFuv6mRTuKUSk1i/Vk1MZHZMCnrdKi0a6dZ3lUhKfEmjnjqF
rCMqMkN2uDEAfB3Gw+kOGYBwTj/BS2XNXKOHBCD48FuLWE7IZLr/qrqQdASP3+yKjv4C+RogFOHw
lUaaXSTysp8XoYPOkAO+laYWJpABeloZOo4atv8eNnUJKTPqMBy4VfO2tAs/A0nJ2bdneq+7347w
MNJeJ8t9D/sk4d2GWnqPjdHw8sYOm3WXjBPPbro+lfq3KDs5EHilfgjEzy3rOOkufdc7+IaB9QK8
+avdWS3bw4l0uP1zrK/Ur1327vqKi1AAxIcjfLY2sAzyFViefRJBNRi//PdR/yor+91FIoQOOrFA
A2oJFaTh3hbL6TRLYJ3UGRhvmTd4ICpn3oD0km7GDXTX7IqJ+3/OluKZMF4108Djs461bRqp+GJ7
lg5ZbEWt5cBckM5O7GjkE9dcjxtyJ0Duoja30KC0kdPp6aloLD9i5RiYrxsTdyubIGk73rf3Owa4
hnN/LcCpTAKVpxVrFEsmuHon2q5aqb4XRv5mAjDQPBzED/9YdLr23UmhJj5TRmDg/qTiRSMGKof0
QLe9bUGsPNmze/a44nzpYeGsMuDetBiSJSaAT//90/y7IOMqvF5haxn85DWs057wTdX+VfD8Y9QU
wxjT5FHEpzD+L/zvCNuiseE/3A0PzyD1gq5a6XStFlqHO6uFF2Neg+8drsDOV4tiImyXrapcTgL8
C68chEzoSEKol1DvAsr7xS7ynJ2/KTSTrms1nYRQVkvcEfr/uoqIXPtbqTEmGWTLlIor88ETb+af
o7CyELYhcu5dmDrMkQremu8D3Pm1T/QwEsfYrPeVjFtLQ46TpP9bV4y43HgHKwSQ2e+Y9eOqHLxA
u8C9r7CwxmbL0Bm3buyBktlCi9gZkBigzlf1r9YnK0P2M+jc8WDdJ8M4MCZpeKeWILkJ3XEVzBal
bhWD7uisO66s7nSsL3yxz69zA3/TqIWE4WMIx7OjiEhKrnDOMzFH35ZYQz5gZMCHWOO2Pr6jo5g0
ddioHN6Sc8IyQhiCG+ytcffl5SnS+4DbF6b3SEclQGk3BxUxlYAFoRvB/yyaeZIqCT8kXn2t95oi
JKXEJJHDkcNklK81dDSMq3qE7f0NQQgVY/kgT73QXvESyHMOwerYfcpMsPDXBFaxHSEjo/h7zoOC
yEroJxUnavOpiHFM4j0NrUTTDrItq+xsjuaK66WXLlm7CZopMxJw4UkKxgjBCUmBR2Koo5y5zIP3
Ng6RtYqvzdvKJkVX+mCNYMJlqajkln69LfbEXPBjXQ4QCWAUN5Y8o8NDZml1Dzic0Db5GdEqlbcN
uhJlFw4jur8ODxUklwDVT8tOYRNrLqmnuifn6Px9EZ8z1yYUtagLdQxVoMkShnb75L5zWHX+CrVr
bPRUkSUYBTUkrJPCe4XqZSBqSx07OiIz/sGVtDRvdQ1/HE1/bjz8w3sTgE0d1zUxaEJJYttTYhC+
B7sez15rqnu28fF/IrJPPEC05R4YhaWCdTfwJVoG16suG5j5kMEKgu5UX2Kj07cIHpkEGHfERY1P
CSIMussGwB+jGgYAFBm5l3Y+omC4pZXh82BQe/lzWkKcbEmlkV0CP3jp6xoLWLyJ2OvOY4+W74ep
ytvWzNMFaTVz2uQttNtMx4lggl1abCox3s2vCoeIWN99mM7iyEBjWgLEHutnxVKweb/U4acDg0hG
kIJrQxQtjlXa1kAS9mlNnchFa7wKC+Xr1pRMzHcUM+tKNfOPge5HShowohYy/AP4mmYQ7Dz5Pm6R
b5lEVIjPR8Fz67m8chobJEzPyjCIWzvD84hku/cCjfYIOEwnnzqNvt/Zd7N2oEiDbUpVmJ7Sk9rq
l+rO6W1adThn9lJRxKmVhaSTaojlLxmhhBc71y0oyeResjw2CpQ12sC8IJKXvo6olu0WGVjsSA87
yyWB7GOtKeJUA21VIQDjGvkPVP71ITHsy+RbTHBfRe7poxP/yD9ONLpiNX2bjJS1mQ3PXbU78+EF
U5Do8GM5n5VYUejnwqauLBiwI9w5uqsdP2FOShsImibWydQwuzXGhU380BwM0vCU73ttkzcp9XTx
ZItEzaOhYcMbHZikUKOuiRmosokG7INrp4AT9DrML/4EudLu4TdcFleD15pkY/WpGOWBr9NyAxVU
vMWk2yKANGxwVAJa4r3gskF2p8X+L69FTlAO2Ai+k/ji04k/ZBSoRxl6JojOGf1LXbxJbAvdqdLO
DmJmOQbdq89TH+FitB9xwCRN8jSwLjZb4Ja5W5deJFUQXyq8qmYpgReBQtUzrwYLjzl7OBq8Spjl
o5j4of1ObR1B+WU402IpVefFb5TV2WBj1Uc/+aF5Bo7pvMwV1COf01h1gAysZHMvx4Nx/WhzK4HQ
7o9EQetAdGEXwUnZ+OEasZzQZLUgU6ggH9TJqcat1/95sAP1Vevg/3OjjfQVPaFJLjPR7920ya7F
OlLm+quxh96qM9NzdzsaAoG3Lddctc3I1MxenhiipmoUEejMyeTnxAa3yZoeWrmRc5rude6CwCkI
ZiK95RcNdtFpsnmy30CJF7LfftCuQ/Maf/qkuiUNdgqIc9NAJ9hyvAaS71O9XnV6EEi/b39CTxi/
QwOt2SypmbjH1X2f3gMGddq5bDfgSfg1ebG1SlISOVznTOgSf1g4WSGJIVU2lMyQ0yW6okK36Zll
SJRGO4Ex79aeFhZcBReehr46MqVrfo8z+LPUob8tv2uEI2hNXFXaLND3lerid9yrOhIg6OGcIAsk
lac7W402MKfEuYknRfte3fEgLFdt+4EUAmpPLMysemXxJDCJMl2Cyvjjau1hPNXbToxPpyJtZ4bx
KMCFNzyImGKX5R/EFWvqzeaQjjSL6/Xw2F8Sd5GGwdiNVV3LbhWBNFNxC8lc3acW6PN0P9L+Yqoh
wyxXM7hvWl5/yeUJOP4RQNats5ICw3vq2nOfHh72u/WcLpqVlICKFHroERKQgLsJosmvY9pzeFO3
03sXDRNCv83SPpukMZR1lFea5ykkwGGy2YiEOHk7GkeXSD7/5TV5u9pOsdcc7PyVJkj8rW/s9pHu
DQ9vNQ5wywztEO1UYM/ZcChvUzpSR1krMtd0PXye/ltSLQTpcyOGR5Zh1ZqmP9LGMNHHcsfU9HMz
IYaA/n891DKyzgl2Qm6mqUw5xXl39RHwbvO9PzvGTLGGmjw85TKazhbZA7JAnYvkcHwhXPQeRIkD
FQ9IXiZoFJvk72Y40olHaTWrSTDmPE7afhCPi7LrPTzcpyXF06PYwWRLv9igQYIzy69UIrdjovgs
kcPHXleKO856U5vcZxh8mZCOi17mQhsBsAM1svcDMD54uQWj0NPFSNdkPlcPk3IJpT4auVXk2auO
zO6x5YvAcKQLLd6k074nwdL91Uq6TY+qf9Ttl0d1qxrPQOjMUZjGgzbtiHLTb2knPi20TyMF4gDj
p2Dwd9lioxnFzF6OGrn07D6oebXjLqEIZBPlin6so1YHn5tY/8ZNimt8dv5VVTP+EhcksIrkOWvr
0B1wHIdbpQz6pvkILXM/ZsiNDJ4jzJ+85wATkVDfio/uHV6OrcMAMiThaGezoBCLxETKiywv/KOF
hbinskocSjDURf1BLx14axISBgzl7B0zWB7VXwd/TZBlyDdzDMEppdw34CSPilvw2atxT9Tff2bG
lAcg9KwyLn6TrBrIN56UZMFp7mCYMRchftcy26ihJXlI5sWQDZ+F/sm6lb+8GQDkokJHCFV9T30w
LA5WTwduGn2AmlAIbfKG3Ly9TaedH5xWS/0oItPeDMjHQlHFZwyKki+15v0/iu3bpK5uGdcoKfIq
z/yPwg2V4OE1strAQltQ3XB5bWTCbCS8ogXK4l0N4HFltTwtAtscOYaIy7clZLf2WwaXZcCBpyiz
vGXfnHgVo4P/1rD/DFl0Jzm2fxVJa5MxvYSsZIR3vJHWQlXDywxZaX6ptgjQq2sN5Bldtnh7Xp2z
yTPvflo1U6qClIMlKsOlgodgr6kJ54od5a+IRbEd9DeDuNG/olg9ikKxPDOdgdJ410E7DSFdXekV
I2UiJhwN/p0w1rMNVcjYLlF6d1Pn6zt9S7iM+thq1z5PcRe4nKQoErUzRha+evQApFSDMRe7olLE
LM9xmMI3djEqFckLJrzTMjTV4MBo2es8a4oA17u1P5oZOzJ+PTJ7dzqd1FNTWx5lM3WuMfbcRux/
VNy2RF8sT+Re4za7PoQ/oEil9ZEoZTM/Rc1OHoBMDX3rN03xprQif8lFEY96b4ujpG+jToZTeksT
BOZ9qpJlN2j5Fk+HaSPV91kzogbl2Lx9ryinDblpjDvA4/CRxMSZ1ogwJDnccqgTYstOMjpyPHmZ
Lt75apcTD1CVtGr13oj5/33q1qGhC3Hyr427WOzsrMuN9HokJAgXl47udma5AbHlNr+gi3fOyVnN
lx8wr2V8xDgR8SG9gKz/aF0DPWdeSQkLPr3QIsw9kIKvmmiS3x79Ln2jTDz56s035fGob7lDWjW3
1AlcXIpWROglV+s8vDnIP+RhJvHA9A96vG7lOxo31J554dl1JRcH05J8aItmyTT4M0kwlg8+ETrq
suOA8uJh+wMC9oUURTIUsuOOOHZ8uUKAlhtTAokTa6XVk6qVVWy4vDbeo37PaCSNDFOp2Oer206P
N8V5NfnKKF6h1n0UR4IhqMNv+73BOc9JiBvBN+YiAQH0FmUKGe/ctLC9E5uIVXysIhWABQ2qKGuz
gUBLO7eff+gFHiSahACEtW8H5EERrSaimuwZV7XaGyLosMTxClRERIPfPTG7e7WdOKjlFKa4TzBa
88e0F4ESSdI2scWkVtHSaU2d0RBAweRxldGXNwWA1wiq6wjz9k9yAuCap/N8EEYu2YDv2dUF81Oj
YQjsJTluQamWjGP31mUVn06Zx8iyS/JVwUjEOrdnaIqkCNtJwjpIQ6n7ABnP82C2gN1u2bp0DlEd
RkDThUcxVDmzZ+h7eATXzqjMYnR3s5KC2FAqNut0e8g7BAqKiDk8fpG+trQ00wP8Nvicqtk6tS1U
R6N0V23ZP54TCl7OGDqY+JubouWzg+Axk6LYqWQkD7iX+CnoZARAJLq9/rmHn4CWzhd4asqbLl4y
OHn9wuB/6uRmZ4F79UnuIYNXA8ar1hfmMwyLDkW/61R5AcFK1C9LUmZTcVB3fUx/Zzyi7CMaTZzP
hrQBCFhc0QAS0B39boWKnAFnTMQB260ZFDKlR7xNmEppJPsefSbgdk42Cya7+DIpdOBvBFaWJyFr
3TGbQNw+TpUEUOAgGY+lCcABefs5hsnz0Vw94LT4FNE+zb4XKjFeTdjSY+ooVWtMgwSWqDfyTv3j
XnQn4I6df1nNhA67PC8beHIT4dAmufq+VOCv7TraWZL+ReU7Sr8Bm88GQIvf11i3aMFgn702J9tT
g5SAJzc5UJTQVbZQcsI9S3qrT02lbdNeYtKnhaRisL8aPETbR45N6KNRk3M0PBER5G+smO+dI4Q/
j3BzsGdOwtSuROOscu/DfupucNQyx2HTZfWnHsvCWZj0BgkU8jXNuMgFSztbR+CRZ88H8gL6ZsEw
qLDSXNQQh/cOdOuSGZ5AACRJdZv/O5qKJx4xdfBrN4cGgXx8mBqniMpvFn6UBD7FPX0S+vd3glWz
5pnsOq+1CIzyo0EhOShHTfsybXGcvrwnanjjw8xYxf5Xcvn+bm+F35SXczTR1UkmOt7oIfNZRok6
c3ZoTDPsjwhedIAPho9qOD7LntQzJ1utWZrb2XU2d+t2TjULbEp7C4AoIuq8KIrbtsXQu+YdUM4e
r4qI+B0L2SMVBnW1ZnxzHpxK8O9t5SgwkTuEtLembg9yuH52iEt4cEVdCCTJxp8aoQzt4fcaUwwA
w2cRKZtBys69RBovg2Ye1tOKUKQl8MaVdBqcaw0zKiuyV8TtowxT4aEtTAuwaekeYKHBatQFEq3L
XtaCjFCa0e9ZUaNDcY19DeDwtLlHXV6jix+uHGNulpyA8syCED9Of15346KRLLV0SFzCtusIWhuc
Ze7mdKCcF+lWddBj5tv32/MbsDKvB0RlHgyAR0KKDA5FhLFaEHO3rQLq+jeX/Qk5wZm1rYqLuEOp
yvP4bYv2nQHuV4449OGJvHldcW3m0CgIPDWP6jAdXQB5vmwSHG5MJJJGOEk6AVy4we9RF8nQaFMH
IFzH2/LZGwNGPkHP1D9ms2duj5zyuvknpTpu7SrfTjGkkaKYEXSMYv5W1dxOAPKocAC/DWLOTTXr
EDBEYBWJin+aFbPihrCjQteJ0EDkFdKMPli1kdASLBDxJXa9F+Go0Rr7nqd4M7HfPhQJmwwNC4S9
0BXSRVrGCAY7/PsvguS32uhA6vDJh5pE6TYE4TLvMEE8JSCc/l8xv5qb/mcC9tSrfvtOB5w4FUrd
0+5VWkQLjW27C+ohGhMF/z6jz+CqTEEGEJmxVk1bXbfdN16fY3oMQ9/NnxpZ9onfs/bqJRzsh4iZ
JhnXP0TXjP6ljcrWbkPACK5eYHpcQRqZmwS0ltz54ITHb1P/wl5SwnlBUwvuEwye4nD1fzgSMk7p
W1SX5vEgRFji9Gm8oKVVMCsG6a16sE2X43h7GdmTuIfbbQwZkulOfE+ct9OuMbIUdo7wls2GWcuC
aN2cgelUKsOi+0/1DcnSh7kDg0b5bc9VKiHtl2hoeiczsuUo11qxp66oqXX3Q10OssTZ4g9IE/PZ
io9nuunJ1la2tjHN1sdNacEW53VWgnTaFWSNrb9lNkDuhwy0Y9oWitp5u5QTAKvYqCy6I6gNhRaf
mGu3NfdZ6IWBVxBQbRnowmmkdlqObVNz7uGfsal/397gyFgvw3wFEisKr5ZXFBCWk4e9xja2K2ip
rBvH7Wco9K3ToDDITTCA5JsCo8ADfR0d8yO4x65s85ZICU6c6rNu91gnz4WjDTTRp0Uznkw+jRTC
irzfmmOAmuchkyqcT03zy/aG9jrwA2I7j7eGXwBVrzF4YdjifWHRX7S5x9xpTLZGGi5iqZx5CY2H
ZElNYcwZLb7melzqGKUdi6cmrRSNzHfk/Y+cjl7rAxZUPgY9z33Z4oHZz5cSHWuHjb80Hvie2lM0
m9qLpuVcaW7DLAev+TIFqtPlo1WirT3ciHwkfELnVIzAe2UnKtdbzXz2qLmIPwbf7/mmvRTqM0yV
ZGgE7/VCtfPsXDTEfR2Ws2LX0u4ybxeXn+3UVXWKcpQbAM1BvsFpR2jv7lNOJy4HSsUjP4gwHM4g
O42dWxgwjzxYUe/QSJvaO2/53dnGCaT13htQi4YVtTdRcU4ZAIAqPyTIG+01q+nbxJQ5pTVmBwTn
Ox6/XcokVAG6zC9YbW+APpwTViImMz+UEXkCzojloHyoDHKlrnEvXtwX9WNXSaQ7RRfzYvkJ2UQ8
EExd2bR9IeHdVYG1NGFYgiTopC4Sx7ybzBRSDOvCVo0IU6mMRsI5Kt1w/XgbRthNsux+o5L1Me6d
ieinPx47f3ha9BuZ01GeZtyqaScNM3eAEn3Ir1aX1qmPUm2KLCAFNZ7kCAOEYSg/cdYSMgxDlzij
xhVRPxWJoox6E46vumgexrD+pcqPueXKvu33pfbzCy2VlNOUEhJcsC5VkNz8KQGcErJMzd85DWZW
7q1Gkju/HeWxAGcSArXhRhiFAjpNu2TQuBqevMCrfdWEA5mBWEkWVs0E38/wBum/341eAwEEuCfj
Nh0bIl/ayo6ICy9E6H+THOH63tFlDKmIbrB1B99mB+GHRbhUefgfeszK2U0t7KCMBsy/YdjtfWM5
4lS5WJNVBZ6MDBwGV6SF1/j6XpesdrDow4TrZSQktux5HWsvZu3FcW0ykPziQpG14AFyWFvdUz0t
wH0CWj7ykSkhH9/5iJbiklHL7xoxJfh13LJzdahZCqnotMF/PUyOD1nZSA3WCIwjT9HsOkgNW8l6
eEqjIJ3rqD+ZfZCMKDLabZPvT03igXZptqR88w0pzLKkb0aoQ+i+eIhMVq0N7IOPGkY2dRIl7onB
kbhbh0QxIxhgdn0HoPtjL3TDO3n4qZFo0zVprYQHZi+XCskOf0ERy7pDcWZFsB3DrrUDpF0iDtl+
r5QI5tlh6S+mO30ZwCxKrJOcsr3YhnKXrTiQ9Vv+3aPK5Ir0Nf4kSlbk0XJ2d/iHJtaj5H2iceH4
hkxnHPGNVoplnjYN5ejbflDGm9xTlawhnE16kSqt3E5KjqpBvfARZxcz15f0+T6RvRnp2ZIhR0eD
d5Tnc2gQ5EzqfMP0R36szHWjWk65jL7B+frlSc7DcIkvt0Mpb93Qdt6UoHpF8LI82RhdxLptsXW3
D7vz95ViCXpv7IIsNMx30YKYuOOHW7JaPPhphtendiEUytnZQ/BmTq/03vsuXxCcu7JnIYoDQwS0
2Tro/7UoZnmRWuz7moSRC8D14xSGsxCAMJr+4BoFRF7bo3aaldmjeYBwgB5yyo1QxDj2GPN39CAr
md/i6yI0KkT/8bz/3UUJuqdDvQXXcRFM2Z4RXA/wnk1BuR3wyh4fDpu6KVgRVVDm/21GkZ4v/xQT
4mXFeIDxsW/luWhh3ehkPW9+6Crxu0VYfF7/+U8p2uYbJk9Hr252rAo50K+3henLkIAnBEY1d6uL
bq2dOIAdzl2a8d5uamZbnUs+4dtBABxEbRjvyuoOI2umi24VPOTG2BMOuP2xDdovWD5+IYe83tqY
K4e/hP803C5oeMaPmz3yBGTSfYvx5VpVUrKLQkW8KGsH9q6501Myp8wXroekFcTxVDvxcXUx0A1w
qZZUxcCrYR9QpHVzvuTKXLrTO7K0HBlrev6JBOIgQBrr02+Pa9hk9mLUAPiH+i9+8fAseSGG1py5
DWjbWC4RyBcdNE0NS5MWGd4RNVph2RjHdp5wABZ4lHJaHbiZUdADdLYYZObS/qNW0dZ2rnESVqQO
X+37JIMKW6z0pVIL1LnMA1Ul6C6oqyM1EXeVNRRz4jr95snWiz9Jb/Ux+rrELNx2XRnneWgu8ngp
P1n/0/tBY7tQAGf+otufS/EAxMdF6TF+k+pyYzD8dTWWGAg2A4QWdmi2Li8+VMjTPLj1/Gz1Rwas
q76IVWofE8pRCaWNtpVuOd58XZSfoQHId0VLH+fBYhFnTEJ3OP6xa2psJw99BKuvrY333u9c9yRc
7CxHL/b6Dn+T8uXpofD2RH4ISW4+vBjbrSKHtCIIg8PADY1MBhZxZFmc89U19l32FkaalJkOUG8R
kJUvR+Ls7B7SRkl+RGtksOBOTKVW/0PkB/wxtRCyhtuvF6U4QqWSvyDznMLTGHHHJcuEPtcGzl8O
v+EKK5E3ubtoPbanRicRg4Z+MKds2TQQG+Bn24xzrzIEUCRYuB/G+B+TWS4JmchJJB83vxOx8gDY
Y48cfHfPEn4vJCo7zzNkuptw519i+JTx3Z17SBjuVTtLIrRTMCl/zjheWsFacLSg30ZPlErEYqgQ
ZYIk27L5f9cc2gRkqGUXDozaCIvllCh1PjZ6x6QeAqn+IpUL90i0JdrAC/ZoRIm8t8fhyIVxl7eW
hmvqSdvisWzvP7yiW0hmvYrpbWFvog8taAHn4AWbp+H8AdPOjulLUO5r6HOF/u+GH3Tzgu1/qWVi
e3ylxWPz5065fEtZrm8D84h+Y8aUmF9cxO+kMcY+3BF8XFKjGbV4FCM4sKmaac9PkpES8j1DiYhX
8/yeGVrx55SpuMKTNAxGqdtaMNVDb5v8wXuqM5zTLn1JRyxcUs0rDuNcMcI6GiAM/oBDJ4du12rD
MUjrYpnTpyuhVuKz4cOJIvw+EtPLVebnpPFFQlkduQjX2OWLuH4PN1fQLADncFr2y3jip7Is8Pbs
E6XWYophx1mIhyv+6Z9ZsibV63HnH81NLzqWuQ46Eb1SNfxEwok8DuHO7RUnkvWSw+ghM1q8JSPt
9s/fOdGAuO9CVbt37Hxl80idyIV3uzENWBaaQt+K5neHDMQFCGgEV/b3QfwlDLy9t6ahr/YHoAIW
t6XWvYwawxm0sNNECZf2eHnboMWhUNXx1y4Ts7ICVKmxNgSapBavuKplN9B8ZzJ2P3fOjGwqv05d
1Qqa7QOo28fCCwnjh4msFKXMt42tvShzVITASO937Wj1KnoNkybmdi3VzYc6F8HGQkFQTC4QlF/u
WauMclS+K/vhguqDojn3yy+HRTiK/dEChrjMN28hRaFKMApbbBvtPGxWgvZmkSbU/nn7zwC/mSUX
L1RauV37ft//TPZ/nUoGZzZkbz3up6UwesbOI4T8uxjc9lb9AaIbaf/hpRb+WoUW0qMzinJTHuFM
nqWtpg3zO6SV5jkuSC74V7+8+Nlrsskw2Cu6e4Jw3ii2pJCC0hCCEBJur6a6voiNcTMVmgx4w8IP
sRHNbm5Z7eu3TzQYa4UxxyWEh0QNyqPKxdMYrM2WAK9spdNhv9GNr5mgD92l4X/FZpjSWjoqeVL5
p7AiqXGkxWoO9PgwkIrhzq3q3oUT3lhz3raRkJnGY102GVwYf9v0p8wK8EpcmLYKT3vyhpApyjgf
nDJB+1vOF+7sD4V3LJoZ1BdeW86yfzncxjEDfR74yZPXbCIkw7E3bUOFE2dkyEGhKdRTXYVZxwEa
p2/mtCtZFXY0iWcwTi5EY6U4KaD4JLTm6PcoqZs5cMNSqXjdbAC7pv6GKQoIBTtF3e+wDGlmPAqe
ltPRzt4tEezldtYRXFC0D4VGfZ1pdYRfUy1JBBb5qL/XBPJcA/q3fFNeG51QylLohzOYf9EoJ16y
Yy9AZv9zxB+uJmbE9VnT7YGpF2YLarrIg8wcy3tznvM65E6RbjRJRi6GOpwRqQIPNXG8uS2T60Fn
nlx0XwIgVgMHJodBU1KxOWN4Gj3pYfLBspdXXFUkxp+AiZExXEbFQRaBnNleeweiV/T8Np8INSY5
7l/vbbgEzIBSo1LkoR/U2yfnsCV1Hrt5QeWmGG0oTeN+OGU9/2ZO9ZTuoBvhJEIlhDcHvN0L+v0B
pa5ANSDjSzZDnnEhu2KhQdi6KI4S9BYPnp7Pmoq2U2Pz3ra/hZAMyyTYE0kxpe4Q63BIcbP/8l86
/lNbQLqB28Db2jcjp3CbMWKw8poVBggjwRlE2Ts6lYjFerzLpVzEq2yZV70LbVWqmWOyhAaTvjOS
XCiXPoKJlMg9py8y1bY03EsbnugWzJh5YIs8GYK6lcxd+eleTX/NtWFu3mZjhPP8IM8CSxlXBXcr
GvlBjrHZZsGv1AFZWzaML1RumEL0gDIpIKjA8P0DpyDFMqIWr6+XTWJwi9wtbD22RsUa5r28sATb
X0VWxABzldMyVZA0uWKuxyJxSIPOOb4UaD3q9dQeBrdCxdfDeqXYFvAwSYuC5y0EAi39It6LeXgF
izVYoC/kjiF3QRDO4bTorQb6QPrP2EP9V9jdFa8swhbga+zgfGBgqgqQVi6vUHVdIKM6B5WG5DH+
BUAzN0DIpjDxaWKN2qjYAj2ajV04fABU4lMTY4nT3wBqNkxjEaoSHdrrlyoSCIH7HssSaXxT0opB
ABjdTsgKed/BjyzuwFSbiM9LXGsGyoEcdF6F5XodZTSCopIsvQwG3DFNErI4bYcku3vxYsxtxZxd
9bUMn5LF8tyjWsyKutKcG+rD2HFyuVX4a/0dz2iOVXfK+efIzAD3Rx/8n8Ulsd0Xk0gSYjTXJtso
RcVb9T2MaxPklgPqfZNzz80CNx0OsfZ9Vu05Bi5h7KBelYunyK7EohxQnowY7g715kzyJzQamlMd
DNlJsaf1nbnyv4loC21xJcztBTajlOmrw5wuQcSfGRCuGCd97K+fxBfEtm2aYx/E2K/40rGstOLK
poEXiD4+5hQtAh6kkPxLKKhifFa8jF+MSjdr1MVxGyHxxHxcNzc2a71ZGGUp3oK7SnzLzZsAclEG
o+rX8e7YHefidb/DKo5XxMTS7vU/xeCIQ307bPPvS1b+EdY+DzD+VwL01jmmR0E8xxd2FxYJqrz9
JSNlGyFFOsos1XAjZS3VLIRAg87WAzpsomJw74NRP2NkeGKKggFrG/kGhFb33aCxJGmy85/+PN9f
n7y1Clmm3gO+B5imteAwwcp30Zi0L6QMAjCre8s3y10a3/VuAjqEweerOjadS80aDfKpiUoRI2MM
rArIPlIUTjQMSv6VFv3SHyzApx6xMHbhgv99aYHydM7MDlFmtfTZBn1uoXYDEXI9yLvbTLTojsSn
YSfsQwwXTC8hj7j93AnaXEMbBJmzXM6PSY7aVrfDV25HLiudZgI68CoVt9YgDrIfSMhcU9merFzj
UyzamwxqrwTR8shn0A3RvX19a9GavssrfkGsRnQtAeILKfM2n2DhlcrWu6o9V/2VsDysm2Rma3O8
x6O4kCp3+nmCCccnW+6xb/8NSmRYRMzVonQ9Y0/1vTiuJtwJvYEq5eKdPSEeNIHHK231VFUE5Q6E
mKaYkz9E6R8lEB75OILflGG7t7WkyV/mFdzqoAKTye3MZkbJ6o8/5QVrjuaHAbLoYnRJblyIflst
5dpJf5rROqkGuVSJNcygbOmXs8XuT/DOhax1kVrYvWBPo/SZl9w64HlMAWyQr8cC6CNiwLyU5eY/
0WMXb3Ft+cuL+dTYIW/KJf4zHWUs2KVjWF9FgzE1n5CvSif5PFj/2itwPL9Zp1j2BaMbsySNOdkX
xGVWr3jN7IBH6dBWmRIiDEoR+s4mMi/FdltyVDK4yu7gwfTMZHuzFN0POZQfyP3apNf4u21w0uYH
36PYVKR45nmuddNpxiF7B3eK+AryOajnVDhQs3LGlf0u10QUNxwyy0Eh5fGeQMrrShpAMvVU7mzS
d//KcRsqsypCPyAsai/domfviFoWtlTKc1UZd4o07rlJwgubPzjIxrHsLkW0pa91/Q0iWD8uWCWV
YPmNMBRrStvXCduYIXVboimS7uaBFq7bRwb377raSCdNGfUeGWZQ+u+Ze7yLfA+w2EosAWDVvkk+
LLjwKUohbvi1HYQywfxm0GczYr5iamGPixe9SfOG/3stSCFLnLizPD4OwuN4pUFAjnt3jbTURgIR
d8e0zVS0GLCzXetv7Vy2SJTB2pMQoTIFnKbgZKRq74JGyBQvqRP+v5Uy4Kl9pftS+3Sii17N9s1U
f3Joez6xGE7cC28SYVKAT+U10AkJf7VNOrlHTbddQYi4lyXgu/7Bjc6PDrOzUi1td7oQyqjzig7n
Ofpn6WvBCWtDsrbT25OeIJ5/V7uMQesmdOkxMhKnUJDKfEJEk5/yFipJw9E9RjJDHzzXrjXCO66g
4WRHAyfUQqalGvmIr2uBHs5ZUfFsUaiFEsE6L+RcP0L0MXdabMfLOOg82dmJbrGNWbIZrReOBCbR
QbApGNt6mxEe39zx1jEDT/kWTv9IttDc/kTstBPjo2fGl7LRTpTVn6TVQoG+vOvWldiZpabXmKnx
3n0co6VZ6WOwGaWFkdZMcmNiI6okqGXXS9ymQRo5VbXqI3rhWRZs8hY0GJkei4R8AUsjBZaQH/0q
QBXwSa4CHAXm587KX1sauJJS89nhJwNAuuq0rSe1eaPsNNfkjTzZMtc6BrBKhsAK/OgeES9mLPVU
QAXvxpLUs+/FZnVpI4D1NfmHsFYxk8Ofufm2zMvGn7jLLx3+usk8DnjN1kig1UhsQJ5V9HuAAKgn
MtIvZl0HVHAgQuYSMh/B/OcB0aDmLJLOSJTXfzpyiosBrbKxxEYw/y4HEya6CtLjrA+zZT9JuXhN
AfgLUj8WzcJJzi7J9180Aj5DEKXu/xFJ7ERgeMBI27Krb95pNryONOFLHMjUEhEFvx6MqcK3r+rK
FSFG/yg2rwabr+sSVg3EGwQH46v/AfadWFVQeDC1M5Ia5L7CnDoqHyLQsWOwqq7foAwPLIOw3hYY
BxxG/bF9mKFXZUuZJsNDZq1vh/cFQD43miWbqSq537bJCRc7zLRkvaU+4dbuLl5NKVrtglljILK7
F+2uSkAsQBbC2TORjUfm6/BIHhQFsniid9Y9Ht/m8kiXWrO4hYXxmMcvlbrJgebjt4BOw7GoKLRh
UUjEZz+qitNALqQL6SJ+FZGuQfyY7Je6NzmLIB76yrl0gqbXixZ3iz9jnSwbfOxW98etMIgv43sQ
pkJcxXHjlHUd9piA6aUsSnQjK5LXvKYjBMBoUWIvdZmsH2DIU/q8W0JSPobTb8vQA2dlW8WXl200
NFWSaf/cpXTZ0V8NOlEb9l/z11YZwqAPV2k3t4vushHAxnbUx3FtpU/7VtmL3yw1yRbWO+GJMiAD
Tud6M4TNroHRCtnvOZ5hhgqwN3xgVbBCInAsRNnKatricQN2UsZC1kTbb9CHpEBfqy+B0/xsJQSD
iHw+OXgJlqQwboSpTn2rg5Mb9cvhrHPZFRH/YJNsENtjt50ORQk25RUhrhwxdBYiGE7CecQmb86v
+PSCOiEk5zugm145oIM6tdCr78uo+c8Ay+Lrf8XBRt/4xdzKbTo87eClRR56+kaVrtdedSMSm8z/
pfiPPJD9ErBlefLk6IKfI4LrYLKANDZoOLtVfYb9wN7MAN2hjZRGXCkHvVMYrgrA10XLD9WKdKeS
varKVLqrsp1Mu1weiauH8LFX0zP/1pQ86WfFvsX/dDRBja6UA+ijZPY2Be9uQ6weDwqdSSkxNw7Q
xlRcAVnOfDACXrm1U85147jx/zQ7DWd531hrm5miSN3Uf9o1keFpPro8atGIEjuiP0wz0OLjyEyS
Dn8vxfwee7qeA9a+Y8OrQm2zUt/U2GIVgxQUvMw1O0dVA/hKUYvzdMcwiraMGTQn2R/q5HxXVfZC
+ZEUaUUlIQRTwK+iQv4q1npeoO0YPkKUL+jZpQvovPpWxJ+BfpXjO650Cr8RvHP1mYijPcD4Y74Z
V5TSYfCPFtXYY4n3Vxk29qoiTTmUWDsSLTSa+OwcBXdND4jo8JUmGGCH9XdV6oz8mbi6dj+cwDtd
sTbxBVR/Ro1M4zxN09kDznN6xTC9ws2HXusBZxJSCHltPdwHcI9z/e1awyxAs+3ONFdjpvUbnhmL
B/6qDyJCWrjno3q86MOmAZ/5JV2EidHq2nBDPm0Flr6lXjBHq/g9j6B6ialRuRq1aQo3msqOxsAO
YmG4/b2F3Nc9S6QS7mRodHrM7NAU3gM2G/RFUMEszswYYThfcGE7Bgs6zeNinoxcWjpnkb5N98ku
FKOZ9QoF6A7fiBt9O8okv0qwnvmhugpzH4kmjxGyjfcymihF4wYXRvgEkHFG7Z4GAvoPOskNhl0b
MVIS/Ef5zONqTWUl/zuzKwPL60DTvx11rmDWyU6nhWcGSsDScR5rjk2eCUr8jSlCU8Ie8jYbgqAI
jtsj0r3/thmGzONLf4CctTwHHOE4knhEATcH3JdYwNapBwYtwxDkVhF5zs9wbBgJQJspLZrRZKAa
bvlJmjh2GIOWwMtvMy7ZIr1m42NaM1XRfJmlNfq+2vAF/T3ESmEdD0Qy4wMncn91bBDlt32xA/SS
Zv/PuRkd0lZzsiWWJ8lXy3DQndegTh+6fjdeqtsLIPQGvI8eK+uL4j6qwlSo8L81fqP7hY26AEN0
uzJ30AlfXaUC+kTCwlFNGj4tjEzr5dCCP4nxqHwkFklLxE2QWEbD6CwSgTO6uYHyn80NYWSGMHF9
xr2QLfDeHS7/wnoP3q83o6yfP7sVXBxuWfL3vsz1bVLJkUTbQLZZ9Qtp7vT51nDVrxCP4I6irilC
1TfBo7OW6p8c6YCxkabTrR3SutXuq4Xmu4Nxzr9V/oJCzj2/9sXHdnDXVZK7MQ3uKu3h6iDDvxR/
0KtKc7GzptRqaJvLYqnOSGAgu/GM7SvzKNkCVf82KQpDfYr9SRA+MPruJAdPU++P3I74LJqSGTsE
jHgS6NrQ6FWuyjdKfS00YoJCs3LsaIqQF157zNa2dPWuM0xu0FUSEgSFdUucHrUSOCyEDXj6qg5Q
xiCygjXZcygFnT7wgVUvklhSzkgVMALl87bC6x0JAcd7o2MX7vo0cajRM8lr/SZ3PELBBL90MCDm
d7X5Bjp4+uthYu7YEmDxoAUFUz7hW6IN4u8xV3hjN3GDlu5tyxGWug9Bc4jRnVYEa/TGTAFh9g5t
iXP90ikD//zrie5469SAHjdfYARZhppjQvfAaj/eqM8HheL3cRp+Hpm1aHS/V/TN7VSR4JV3Bt+f
oWe2eva4iOq5mhLaDErN5fFivMLn8+Mseb0TcWf9wNsA4s7j3To+3LKt8I6cKiL6AFBXveN/uYdz
tRl0dVErPbKEQUIHIfIWK+8z55bYZ+latKMi9wV61d07KCYWbpOoc1SzhqchD0ELC8uiy1AR9ltc
fBDDFLe9X/B4/EEwQlmbvWwfaLNGIdmqnZ/uPaZ60K7/xPexpwquMzmTNqY9r7yjLNsfJzufAhWp
YjjXNvQscjIRCZYi1yMcH8JFw0TXhNyyFE/nnIDZ7ZcOw2L4G8fo8j+P7Hjd88grAisnLU1OtDqZ
WKw1XSgglBjz1xqRXd4ZvrpBNQcP2CeVldVp9cB0y+L66UMK+96D3+HlZKUoAFzeGgIM46tuH0fH
5fj4m5LyKsc6kp70kWpZFmnhwyEt2sWgFcdLLKkzx+6ENpAEiWxqfAJlrgJLCEq90Grw7nRKMeUX
17XWn+g3jxh2haIGCmqMAL8YOxDCCHln8phQ2151KVoZOry6RXrReasAXxGiPjk6ZsFL715Y6mkW
t26tH7USdluiGUWyPDgSCTXBgbLgpfC4BeGIw6zPUd2kwrQofAdl+XH6Z3EM7Dvv3GXko2ti529T
74tMRXSjRuCJYyIMRyih6FTCXqyPLZ56BMgAqxj42axlaoKsIhHoLnByuvAJvBTYRsaE73HOlQkV
E7iP3S9TZfFMM0RmS/RTOyMVziu3i9nY7Rt+H1pJAlDdnnKP/62gKiuAePGj/uHSVm6k7BrnNzq7
4XdYjHpcpkoDOhFbaCZG2WL9VVrqWs2eIUlfekxLMjSUV1SLMrkAx16Bh5GdaDdwYg+6ODfHP2Xo
N176stPf2d3LfR36fgeh8E+tjCbKJuzwZZR2C/yxNsrYivjj+FogryjVimxUEXetR2DF7NeFVBk1
VQNxkf22IouVUmI6QIWWTImwmAVZ6YixjSt+Bz5JNm50TXeYRTHD/OBFxelkRh2YEOlAoXepBXQl
zlkdGxmlrHclZcalb8fmtLbIe4z6ve6zTCphgt97kA28jQH6MepzyL325UzCfpGe4+e+azWn59YE
VH7yP/FmEbSB8q+Q13SIsV48qwvVoDKojJkrbNhFM8vtO2VLUEJZKMw/fPvW8bu/qTxGz+UJINf3
4aJiv4L0awqv/lgLDhNszGHI8kKC32fugQXxtwXWMScCIZaCmD86O78j+GBGHhH94PdJYetFRm0B
SVCah4FIe5/0TvGvn6PJcByZe9ofzNj/Qg+sFbokdDqaA7Q56GBxAQcYnwPIwGn87PSfU30qVw60
HP7H71ciLOKdktAwJo19mFfBbdyNTlH9gxxpVyecgyzjYvm5YFNkjMe7gJQBEXANaAsnR9rE2yp0
TUNeCu3H31pBLpXLL+aeShsslrOiYjLSMP2Qp4+rPAGGo2YD3xLVe9k0QDOnOxv5sVFdevL/t7Em
FqppmUuQNTeIuE9HH8+eBwKBaWUWdFeDBR/yyA0K0dxfngwSO5ATjqK31mGIQz4okRhDq8ENCbCU
VzReBbtwUAn8Mb1i3ajjWU3Nqjyh5DikwIfDYspzQ58q7RMOHP/KSDH20PmNYk3R70kEYLEW0Ov7
nHWJZ41MEFRbCS0T91aGHkyDT6FcYD/Zuo6BbJzFFIQqeBD9uEvnsNDUDEuzYJtJ07k9AzCombCx
JF+V+HKwcA8yvffLc4CfpFlWDmIYI5pbWJN3uV9SLt3yIA1/5WXuiRAmwJVhr4gQ4E4BcQf5Vz8M
lkDUGhrD1PGgm3jLZun9Cn65K/0JZEX1hk9C/PrUmklTN/z4ARId2/OtGSRshUwB/X7ErpIt/03t
A1+Sn0YmgLVb/jnZ0fQ7dZZ38QnSHt8avoOk7129tSbuFjoqntZQN2pKwqoydOyRk63oYdPkMbCh
4UDAJ4FBGyAjtOgKMM0CjtVrvqfyo57OozLHyK+qvRFhTaKJ4c9bJ6Dw/bxks2h63ugktm/itKNO
TVfa2/9Dx1/ROZbLbiYXMSJc5BzrxOTKXFFfllZED6no9D4t2ADgQm6HMumaDeH08OEV4FaQbwXE
IfLthvyQh1UYSMWvd8E2PaE8sii1RIpOBFv6g/C4CqRb4qbThoNnmKa3zK38IGnUJZYSlARNIOCS
qt3wc7RzZdOS+Fca/KammDNi1hdeVTTDZUC0wVUo/km8w+9+XIj9BcAatqj1V+Cv/lQyiFmX7J/6
vrEr1XWWmZ2eC0HK4Df42vkdEDaeKyd49vVKPQyNCwo3c81K+To9G/R+IuM8MuDEjPZ7UFNz3IMY
CXKtw42GGraLwyxvp3b1H3f4Ec/3HdcyjQOSLUALPiUkG4i86oV7ORcB9e3Zj/SHRvgUk5aC1W8k
dMMC2v3j+BffIMyGXUSeq9p/hPAcZihNVrAVDeQzAMtBOCQkvcQ/U7+b5mlSqlLHkgc4yWSbX7Sm
vPqxgbZ1392V9fQRkg531cSApOCIEhVJGaUCw+z0CdN4if0dmOET2HJ9/y//WcLuT8drgpAzarcT
fRaql7VeekIhdkce9BceOOkGDu/d0OJns61012+BengWKUs7n+1SQ8+EiRvIc+x+IS8YxXf/Ynth
GKCIeXfmuZRITtZHly2GfyzICwvHrd+9ia7X5MMQTtm24QtruZTl/E9rFkN/5idV1/RmLH7x/9dD
GqZfGKGHrUaQCy7VXibFXYE0RdZbyLIdrPd+43k0M1ukOLXlWShySufHX0WGjIOs78nJpDLgiMsh
U7umN9kHYdIPnqh9glK+tGUh/3bJ4+6aG5Q58p+GLvIWd8sJndAE3wEnv5bM/44HrFALGf1st4w8
8RXQbfJ8osZNLs7Bpq2QeObQeVtS10MBJX+k6SkMwLQvpULIRwmzhPKCfq0UWplliLt/fYFtaEGU
zTdJRA41QcARfIr2qayFK0J8q0MyfWrJjABACGUuLIiOARifUvZmcWAaR1JpY3isbAaY19BOZpKk
dx3HrIzPq37P4c8MmXmjS4GQq0JHcS9rDJmI8LQK3TOoXliETanOyw88schmRp4utwLNbDiduStK
BsoPvc3fMqzGYGf9/poXok7kIlccOYcOTk4jvIzQ+7UuMWg0a+UrfeeC5DgVLzEtHvPn3B8g3LqM
oK19f3PAvq1+cxw12NUEEKEqoJFAIrKq8LuX71SWX3v9st/N8tiulPc4xvMhecuFZWvUJ8eGhnp6
atd1WAVWdW1XcbtwM8XKKmPpM3ja+KnL3FrSC+WkiRQf4SKQcZXTnbbpmQc8VlhV/XBeeHpAZ9IY
vBXo4N8e4mkGBVN53AQEyVulpwpUb/b1et0AnDmwq22aP3ETsM/sZuI/AlGD24P0VF08TxUl42d0
ulTF8jdc5jL6mr8Fyvt/eqbGltU+P7Xel7EDKwBTMEXqLSfkFZ4OBb2l96PuT++b9QdYCCDqmpBx
U8XAiZdl0AFHRzZfTZ43+PzlIk93YVhY6QFbBKS2LXqPg1uZUs4ZQX6qICVlY6bcN2MWvblZpsqe
Aq913gTulOyTG1vL9iZpVrtaHIyryHT6ieM661FXXtPlxk1WCJ/gQ2Alm2UyYaYfBlTjL+3KERxT
Uo11+1TQyW1a6oKhqp1dw0V8c9ArcoIoV3+sOIDrI1j7ndN5xDY4/+RIKJzjPhHyacZc9TR+PwKt
YNnGCh3Z8BS5djd6YslexBoUfspmAzBbJPZidlas5eitJkxnJBk2wsW6r12ngqRRNEVHaUnAxbm2
L38QPr78kQOvImeR9/I7n0TCWjcLF4G7y3jxRpA2kFTv9flj/aoGi6GqIaf4a1RySNVFF1oRqdRK
F/mzvxKIzrwPYFTxyguRpPvuBmjCMaUTPeRfVDmOt3zDhJhj5hdNXJoLAQNdUaDFp0HUXrT2hyZU
qqwBmGYrotKGV0g8frkNM3wtwao3mPR+krDgR+JmLlryegTzn+do59BUooZ1XDE4B+XRE6qZROUk
OX7arvT7voQL6yQG72abtQi/byZJ/qwdEaM8pFnkeEV2Pv1pZZOMBlJRnK61fBRP670hLnsyzZ4R
1YI/5dGNin3NlW+HZqFu2F+wpaQ39/hQiYOqQvUZA9s2Aikb8EEpPocLSt4gs7DiC/9kjrJYy0x4
y0Y3bjUoLDoDq8TzWv/5QxviEO1x8U4FDVJRXdsZF+S2WEydt/f1spBcNQEdR9ruREsNYkPreNz1
xihfNrNivDOXj4sg7k7bCGNmAGA470C/PuWasqhpxASAy/Rpb0FTPyFM7MtP08drilYzbusp6ZKv
7+FTLw4rpzyqtXMMTBRWl+nbcrouWrmaHK1rKxxMTtpeOVKzA6u5+32kiBXSwOfQ9ZFA39xLvfL1
qhvIxT+hWquLvPzWCFiPs6TmFHqxF/JjBk682837uvuztSYtqnQIXyL2oiNo+WtTSYQNxcSsSGlA
QIv9ZjccOYBgvM/gYw++e5XaWAyeB6gjS5UJpEky+ivBL0c4129I/j+5gLDqVw8wKhIvCQj7vnhI
m90CEpLfk2BkklH9JIUtiKmHXlc2c8C0gahuFfsczi00mjzNBrcXrvgz8JjceaHnTD+2rpEb5TxF
NtAcbIm7zEi/95fuyW9wnBuSCa+fIhzjpdt1O+JfnJXVVakhwSoPBR1wsyoQS9AiSD/aePp0aqcl
Jlyfx49rgTfNRZxHSGs+COOmW0nISOfL99WBSm81gRdycHybxlE8fVjvHOMsITVuz4RcSOKvfuWM
Sxoej5Q887G1rJ1oRJrTXzr4SMsLAWEDQy0V+viAU0AFRwuaoKOeHPMN2rfG6N+ShXVEtfcpKvaw
OpWuWIJ294Cus3fJSh75SPsgwepHURuJgnf7QktgVIIQLEGMoK0qJTCwNmThInSb/DQbcjDLpJU1
tYbmRGCn8vmY6GtBPows6ESTyvoqLgn/BkhCHd2ebAam+S1JPIcAmX371V8cGyRFhB3lgZZQl7LM
BQlSE14gZayLEKGkGIK99316MAdmpDz9GXN0OdJLISVtM5ETE/70ImG4qTZak4epI/b76ZGm4bZ4
yi5GBJx0SmmJC6otmM/tFN6iGrXGq0e+r3IS5Y87g9XCMJdyKAJJtvBd/ERz8/8t+k5OL1p5LDiN
SfH8XgDYuNiP7GPPji52r2jzy69iHIoJMV2m4gby6YzkHQBv1QwIwEfjc5dCddM5DLXxU43BC1Gv
nZmEmcr5Zl14VMYcLI2ChDeAeBe6DnAT7AXhSppHSuk2NMA4Y7kxHEKCc4Uc49kmkrH+pUiXpuhF
0BQyEgfQXKbXLtqy4ENVSqs3jVw4qZvstht0828GhsVZ4YWKH7j3y5gKUHTvLYMjQnpHm8TzzXqj
lbSlrAK6j9nGEbyI0GxhmOY4/8mQ5T6WApEG0f//MZKP0BUuNt4ecNZnV9U7A2BcBSeu2/EAUTn+
r5tI0XUyEkOcQK4LkfMCHhH6k6OCoowbgSRyUkfnEioeonfmajt0k/GtdNhzeRi9HNfPureEP5ok
fWtcPBQvhAfB6cbK6rD1zPBnB6q3YCtH2Hh2kbgc9QECtkWXGaU0hTbhNSI23HG+J+XAdeuLJrmI
bgp/q+j84Zylp9JGk8zZOOB252IMa/VE94bFpTRXSG8QROFVcQJq2YAWA6ImpF1YLzOx7t+EpMJF
besouDvtyZMo0sZPQRRxW04KZsWQRkApMO5FQs9zPG2ILOsQyX8CtPbAEWjo99zUxuYA1qSrxFba
8dgmndqHjFfhzTp7tP+7izSglhWFv7ClAgydnprWqb0gACIZx9Hy3IzWhPVzDuSs4seXYPkh9NUD
H7gT9OfSOt8p23mHvcuFEe2SI4PS4lFxaOVDhkpUtdw8IwC3uqBXc54uXEz0g3nyagiy4iwLQx0d
COJdDEHKwv8IfYmyGpa0LQ07mEVd34dsTTjsWbPJTWfO4lfRoj+3de6p8OOSvNkx9NxsgxLFww7n
5R2glHiUj4/5HTg8CQLpo+LmIbe6+BDN18s1E1+O5esBXSruOHkfQDYIcdRixOyCtk6hF6mQcUdU
cmZR6DNWL6m1Z5siIg03TTS5lp5jFp8Xtwp5pudEllKeTact73U/0FsJhSjZWxl6yTIUw5bMOnpV
oUpatcOMSvK5VnlenPpMmbjiWdMc1s29OdLp40NgpF1hN9z312NNBQ8XR5MIJorm+/j4e/Z7Xyxl
j0fBJgl84yTOlVTE+Fs63REkti/7g5pQVAkPaZ6hPr4JKTE+IWDMAH5+fz28t2xIyqHl8iRncXyZ
Z6NJM/6Kshl27sxEj+f0yIko+Up8HI6Z3bixct1RlKjTLq/iZXrbJMF9cDDJYm2l5LsbFEZQgUV7
qNkOu/3Rt1JQzq6A6CJ7NnI+6WKhwIsS5FPDlA/+OO0PXSwPkNytO+iPgwuHbg9Bz+lcOdCwNbQ3
pNgcYm1lcrmvz6F7JTMkOfEIOptLqG4YsI9hBsz51ZNPcpuyZSsmAB9NARRgz4FzJ6+RUJChnIJ1
tKvC1bz30AsWzPDhS3SQFe8BYfp6YBcQt0yiiL1BVN3RASBIUtms/GDB0WVPfHnxRhLoYTxyjZ5Z
ILXVm0lDAWazKdzp4IQaKSLBbOA+RCijSAJcHfqyguH2X7xLbS32PpCrSCMs2EgwXP8ADHI/Vopg
cxRfAuqvijYALRMFKi5iGp0wVSaQjF1VDVeW+TG6LvfmZTNnMQd8lkP7uP3MpSXiG+J+VY870HYG
i1cngAyR3ixAiNvGBvJrbtyhf4q54ar5pK90JtzWFj1EmWCgkxnVe4bkbyHr+xjl5VLTNudyM+Fc
ecQVsuKcKTTEqucYAnGP8RAtJn1mSJBR1Vz6t5vGOqfRvleh84pC97DdYp2CXhOV97KqgOl2ZbHM
K5Em3M0GZqV/EkLWUwtjjqUwXNLMZUi4dzlQsfSxPHUpXsaCLs4904N6+/QXWllsBUDYltcTJevD
ABJDpnWy4+BJYwgMujZ61Kn/C64zfqJDm3OYoePjk9XdubVvD3mqvYSEzeupVR9lOERFoqDqL/0f
S7jpHRsRvcW3MktRvBl2hmDjKxtAZfnlcXWhYmB0WQRYwwUiNnCdGZoCVIE4eLw1ZRDowCO11PUe
qHGwNCr5znjvN75m+lxjOlxl2kUmlwJTws1Of7K9X6D5fr7OYV+qIyN/DgHydgGb1EWhSAuAwHBs
B3Ec2J3cnoo1AfdxZE6dahbP3oZ/tUyBQwWwOASN7ioXOC0DregZrKakUXikbmAA5s0zUErtiD1t
J/1Tf3yoIxwt50cNcv4aMZIG+4CbJdBepAgni7Mu3EmtLIqL7ZhDggf3YJqpPLP9ovybH3gL2UDw
sOrSz5yW95D4rsWGe606lNipelbjNpbinZ081rz3R73pTscmHx7ZSUpH28UjvIoR6wIj2+ScNs+Y
xvTFpMN19Ehwtw2knjAI16vd772oXFbvoHdW7QS2hDB2uXOTJfl2dbgEmxaAV0XNc+hBaOTfBCqv
1krVUQ4VA1RKSJcJfmCi0aNpFkz1jET/RbTtBhD3fweIXB6kosXcI4i4ox5dmXWI63H7cXzXOIqU
NkcbraKF6dkS+0mvKaC5ga7De1fl8Qx/q2OCQkoXZRFyfDYU4ERF/IZ5hHCzghzMiWv0B2w7pfCB
q6lg48b+tvjd6xLHMOmvY48jGcZX93As9ef+X28lb6AwdBtxS7rXmF97wW79LdFlqHBeQOycjYDN
kt1wJvdQwWPQeW1+6RNHQO4ONioyH1g4NCp75qeguDFFtpmcgsIjc9Xvb5icZp1qAvE90ZP5jp8+
iLSSaqvxRT20q06RWaB3LkxliuHqzEYr0PnygA8ipoqcatpf98a/llBJoubNHWEUpwa3JaleMjmk
GvHVJQl0gI0oi8URAM9ZBeZELsY76pEZ6boQUyepQW14n05A0IlAml2YHbEz5SoZmvlVagABk+wF
6E0CFSC91yFrFBuTu7AzPpBcCuftkA7k/adcDN+J0ox/ZI/BWSBSi4CTSW5yWA2OmaQqnPqg3bAo
zgTI7TOPkk+d3/wmfJZPN8KdJp+CQaQoV9VW81Cv8FZI3Z8OI+C/PNJeJGRmb/+EVjT7q+Rd5NWJ
vZzlpCMnppl6m+5AKjOMdGHSpgK616wXxN5TZzcTWFs+SvQFTE+LxDUEU5f5oBQA4FkslnwffT0y
OvydOLP1O9BUlh9rZE3QeJIiJf+Dx8iax81YMvt1JrKNvCCx7GSgImNQqxVJS2A52DIFvsSUXQ1w
sFFAKJMfqndNO6p5ubaHlNb1gdP+zGvIwL/re+hZDHxNGtGrkQIZXd/IrtgVaoY+gqJCgfWQlOCB
ZVl7x6YB7Ki9dVDLj83Rr4jUOFlG2wlGESZWBAwli56ydjaLZ87KxwHwXdOFT73nYFXgkNHdZfXN
tck5kFNVZuhlG0fOHj3qgwk1ptXikYzvZwG+XAxs5hTG+pAGp7RNpxluGZcuP3s2VqkY34GzYe83
H2wpQH7tOHHEOJ26Y11nBHnV4UZNHOlJUtRFKurojOE4M//TvRtlJ/OowUIbP6Pci/CUCrIONkH9
N+rhOngib7eS0stP2ULN16bl7M0CQBthZSAPdOvO4wuQ80y6COa43TIkUze1kq/X85rAEWmsMY0k
PGQw+vGZL0f2DwzB/fSSkBSbVG+psxrNTjwRJzzKgafWwEQMz93VGmjvRN/4A6xJrwBgtCqmv7Bj
r7ZXomZJ2dncgYHzoaYUmh8/SyXY9OQGQwKAH9C/HqTrFMW7E7lv5rAjDD7Q+1+46NaN4CM8UjYW
FWdbw+K3OEgJ6vkQdORRmzX2+49PXc/yUHS1JCA6BUWKF/H7cAhW/5hpiue+GJtZtA8EXiZi3+18
LOiDcwM1UmjNh/ysTeqAdTggcwUlBJmQiJ6Lw805u/DJRUL7TyKrhN+KGWYfWN2XoMx9cFjpnnW7
nKyBa6LJHIfHyhGRqbjmStnlhPt+Db3W7bR1pTCYerBT0wcqThh3/IFxEt3O3Fd35kDksfOgmezQ
6SOJP7iV1HTr/ja4OpNJGDgu4LnQsf4+vn/7Zy4J2fuhrBrW3cYcPNNBT/SOJnn8Uq0i7pT/czOT
R5/BIqfu7NGzJnlcWGE2mbdUkp6nLrifc18yh+FqrnPBezBO5ARCJ5IP0Fp2dDMPM8fc31tkeJ09
Ajy66nqZzomyCaoX3SgH9ROpCBzpH5lKCUYaZEURSjQ0piRjb0seuzNza13zBNy2O4Zf+7TmCDhu
E1hw1sFk5F5/VIl8AEH4bn8vjklt4zAosdVELTfsPRnpk2Gb7sVkA9C/Mx64HtqlLGQhXMY4Jq8W
Vs5UCPnQTquUK/ODK/9wfW4OoSkU4KlAyqJEdTA8+0ajdSWROjCVSONvHUm1VivVKGbO2mQfnYGR
XTzCoOudMKXFGSMH/AC3qa0o3zuiZ+Lj7226l2z/uKqLxgnG+BEIoRZI7jzfSDUGpk+9FOHIZRaI
k3L0yJfIVdvKkNdhev2Bs1D1BD4TTKZ8RvT55jXVod0+YYuUCv+DRBuZh6TYxpsTKBk8YlJIrQQC
q0bKT4/pJMvAXORhUOzDtqoU59gFNXwPbYJVOpgFxS9+pgrq1YOQFcT0xXQM/Ep3VeqLQh32SMIh
OapKg3viDrk645/6wOPCoy6ibomRceRRMFBWkjvJb9Jow3ZpUgAEWpvaKtFALomWYTj6pad41CYs
g77KXxs2GSD/HUlRNkzqGc0SdAHndpqmEZ38s1e5i0YczvPiU/rrV2xUmRSKBmjR5ms1I1m7+0kf
IFq09FMDf6y+W5zAbuHN6ihKum0eNi+2P6f32AxiL2gx2zsjRSwoqhokoYGjAi4oFoVIt8gxKCyr
3hUo2rMMAsoz0Yto+MdvB2gs+a0V8+ipVUwdZIVkysWBfouMKu/FMUFaehxRy77+gw5QDm7xJ2dA
rMTvoWjzfGD6tn40MyrDcSUvoeqVaWCMpf1jbE7E6ieFHvflXJONWLzwS65wdLulKJl3WE6hOY1u
W3hGZD0Z6oRmq7teAaAaYaakkbAfLhGICD3mFndNfUQopRKPWEbiTvNNgOlvSQWQ9de2HeQEtmxe
xMCHiKXsXrobBLcPgk1lOVQQ2Ktbf49K0JxuRJceVsCLmWXt1RkOsauGIPUDyj7VDs4T8UOLFwEi
DC8lxnmbWImo1X3MuurX3iEfJPnS7RAGDtgDoj2OgrDNLWero2ri+oRgH62zgxDjylgCV5W5LAa3
w0l3c0RqDKvNQgIOwqExJC8ULGWDuzxGMWbbRorlu27Zc5+XaHsTh7hLqaMLqAwQ4pMveKkwHMR5
5CWqCTN7ciVRd/ZYnFvWncFaNA74G8uIPGS8aC3M5L7/tkz6NZMv9pYPrkvHczvUEG+mD8DsjDKf
cRryWNPzPTb0mY+ewaHRuRoeh1rnGZGGImgcu5VUT9uV5b9IYCCZfl+squ9h6Tjo5Hpygu9Xp5YR
wlb/ip6krGLF3RBfVOdqXBCwPJOeFuGUb6z9ihiBtlKJV5jBrBngp5AxW5wuuZiv5FUU5M2DGYi4
f9On0ByT9RtJujdvcWNWEm8uCOYKwyy4Ykf4cCgTFf8bTeVJAlr0ql83dAUjtBiSbV/LlYg0awSz
ocleGS5vXfcZdKG+TAlrQ+epaHG8EaSdRXFYMti+j2kmoDJi4wftUIgmqTitsueXWiltR34mkAEt
6Lg+RoQMvA+A/pDaIvWaMDxNbGKxd1Ftqi8XglYMIKNxbdgf3H99DKxtUvJWjNKE+//Z8ehAK5bo
rZzgB640RNuKJxyXNgpLQYm4EsdrWu9by3QDTYbc9fYigl7sXIMnZRm/azn6jaLN9R78WWC0Rc1B
5mVlsEEWqlRnQfqIBm8BXo4TBdvtelN2bKYPrHuvIAKfpa1eQCyZGQMfjx0nZUWiTo0CALg4azV8
oJmM5MicSo+ih39RW8ju/i5pT69Y/boMigrmQ7bMlHD8HhcoDFbb1KZgCZfnyjqGp2UojAMCqYoT
OVsyb1mPmad6xJd3E0jRDC9pwOBtgbhDd1tjJCWjgoayTMG0W8zV6B1AIksuVk8tk51HbkxzDCR9
iT5KaKxYihvUSt1+iNC4MNOqrOgccvHeyZK3yXnhLZmkYAZxH7ffGgTHFM8+er5HnJ60+VJPc8HV
aIPIR0cpzDZqM6IWu2nYGNXrL8gZgOlmrDQJkt20XEup69P/bHPABVOfs10FjO8jfwg66vmsay0q
kA8i/cHDn+MBwqKFOxGyXpAyEQSGsCPjDjLYfSEduzPRxQtN0q6I0geab5PFa53Rx0jbm8rqRmwe
iU5UaAdosNUwTN/L0kSpY69SW7BlTbkVNvKBhyfhwvf4IxeELOjNWMIKibs13FHLXhm2dumP+rWq
+cWp45w7XMeqDsvJVWirhkv0yG4UZ4JwC6wx4dEDsSQOVfgu1XLKrGrRd/Onq8BjBwf2Gu4uKgtK
PxLiOvnbDXpWHupSZgRVedHqjctOi1BZwzbrFtCh3hec+y3o6mnRABX4ebJgIBQwEFYE02Gqy/kr
3xwBK+kn6mSo4PtVWVd+nONIvPkTkOdtB6ua1nj/tie3LggYtWGqltnJ31OQTFX0LoxwKJhiO69n
Y55RsN5inUBY3/k3EoZGECcYeC6vlsT3iPVWU7MmDROxbfWL6Y819qssZgQkCXAdetMxvJQcOHAE
F99nhnTLNDp79wwGoPeI2S2YB8pTmUU4G2bV279isojVSRhy1VEg8L5Nm4/ZKGIGLGK9wuJUvX1c
X1v04SZ58QaAIAZK0/MLC9NqQWoAKYktdcvlkaPz7pIdcbtVwrr20L8Q22VwUegYydbHfpSxt92p
PjdffbZXcQwicz5NjyvbItb5cD9ZhRC5TQ3ROMNvXUdkR1hPB+j9my2n8523X5l86XazvQSow2OW
aP9oYEwOoLhFjTI61FeifFvQ7RXHpFHL9OoAM008WNc9h4wsxbXX6jsJ8OUZYmBItqnBuJT4RsZg
BicLE8Pva4m4AV9Q3KUw5tvTMJs4cZlIEZ2LMii1veIV5HLWxgyRC+AFXSth3WCzc0zadeaN0alM
vE8oRNlgNjZpKv78Nz5u9PpOhBkQFtJp2okI0JwBpFz/VGIg/SefNcJmu2eWYGd0Z5T7gPGaoBTE
dE437LWc07CT8wa46vzctS2EAPRZhNIeK1RFOE1ShTFASIxyKG48nOaB9+jXi4mHwmXfu+O32TKk
qvB3hvtFjQo6muaKPRRRtlIzH2pPbGaXn9UWEf8O98UT6oKuuo5N2Z+NIGMe2OpwM0oKMSEOs9vv
rfctPSBCX/mNgYOM0hFfP10Fc880a+neWraUeWC4S6Nq6R0ACfhPgQPwlJTHbhd2i8PFvUOrQ8nH
AjMAEVojVii+zmrh4b6joThECuC3UsMeQOcatF02l5sf1Skqx/8XOwTRGPiI/WSoCpMmVZXyhuNz
yaAqiTfTlqrgonFnsaCQck4i7CXwX1XrLnLNMBLg1FprrmkugeOMmOejSq/GymPJtI6YRWITVkfu
hESPxAnfYQyKVTQA+hUWD4ADNIlnDoti68ttdcEcSE1dUY9Yk8Cc10h0TvrIAZcpc59xv6lnB/9u
9mdAvJ0AUrLS8iQoRMXP3FLII5Np9o+TGP88YbwZNzbEWWEN95TtTNBVSXKICdB6us+epicI8cDE
NRpQKG3jQwjfnlMB7km5IwC2GaawN6WkXSfDOIx3kRq63aFfgmFw5dMJjS6V2YyojqqiuGzTUKpo
YRgT3TPnwlW3e+9TnXT5Fxaa36NeZpMSRuARgkuOif/4hkCWZN2UHK0EVc1yCxqJbKNuzjB3pjRF
W/xQZDoTPny5L9wqxVOMWVs6FVsANX7ww7VBDBHLVOpTMETK5sbtcCyii+LK27j0qXRlOi2qKLrT
5xkNVbtLdRsWHdIqpHou3/PhOKhNZMGw8g4vwgf+Tnt+vGy5izLXO+k0UuOUeKScojx5zPjdNseg
1Mb4QY54/wDNZibpPbZV75hVOFEvLDNpyThTsKX4IFa832GFEbfaKi0OAVocrIyS5PrSpErHlkGo
NoadnVXXEHgd6glV44ZTkZZoX8wPpN+w0T9FBO8w8zqqmmsaRAhGQTx/1G2i+2Dbd0BSYNS1pGsa
rr9MyZdF3YDSbhNmHvZw0NA5b8Hrnc/1EjMx6BjzKstyePcVgK48NlMIu1306JzGxe5wib447Wjg
QcMKLPdvewxnbRGyOKzLP03EM9HkGfRVDDwEDtBmykpB8bV0P2C7WfWLahH8ynxftIapksLLrmo1
gP3VWJGZbAvBf9U50yfg85c8VsY1ZqACofoAyHpvBmZAp5vLPjKgon5JwCplbVUhCEgyXLT7IfGK
ftpfEqL4Kqr7AvdggI9ijQjyqh3EB74L/Fj0xmEWl6jcdLAQaNH40j5T7bt45NAz54NTU79VHYb5
mP+v29d9yV0CFtZXZoRCU+syG+wxsjC2Ffq1Bdo8p43c1h8wv7Qqi+8uPoNy+n43zNncz+EDVU07
aSiPBNwJPDL/EbBi70ANaxE4C/+D8JGuZRrHGCI5qZ+DH77TCAmTz9F9/UDWhaX5pBeyRlvcNIPa
ob4OKTh2JFcv2PCCniL550pBb9LbNYLfD34hOEkt4lA/24hepXtHOWqNvLcKSRu9kFzltwaHKyuL
iEl/AAkU4CAmVWu+eyFNVdZa2mYo+DbtHfibyeGLI+R6NRhCxTKEs51KqjHR0oTHdHQxNkIrR8+k
AkovTb3O3zU0ZK8xA4FWNRdZ0CVtenS6iDGJ9mSmROrbm8hKAWlEl2RzqMSH2hYVP1DG7msnykRE
9VwzIYbZJD+2f1ewaa8BBwtRUTF9oOR3yOKZhqXPFJT01OUPSMo9lUEV8apFnkvKLut2yu5bzebF
HozvNaTFb4Du6DSwQ7xrF1MDFblxmkrrB7cbt5U7I2/dhMu5xSRrShPmo3DZO8Q31hJsxwFTRb4r
nw3YkoQmfw1RHTOPZuwOT4ud9PGTrMHZj/X0HdkzvfvnBn+/bMFcLK+fRf4xYDLWLLqPEJX3VHVU
vfEeNh+SJ79TaPyFCCXqdFqeJEXhk3Y1Fi4X/WYjXrwi+etOKnF+EDFyRcyKf+zl0cJm/MrmYElv
TUqjNixLPVcSTF1+fMySnI+hdH2D1kPGSSuRRu+BNOmA9HykgEKxfRaCokaoOlBpstwgujGk2YdN
fIDQr9li7QUR17+jRFvYlmaS2GqXCji92xZPv8uEPiM9R8nqBcfi4UZXeA3+tjiz25IApLR/LePz
MEfXOF7Mra2RkXC9fL/MUdbJPaA/ZsUByrSrXKbbe9EgUWvZf64+EdQ0wHOUiZTFfz0KPsUBY23w
uBQXN+cug8ggkbzfkdjm0ssoiSHg60E/HS5qsO1nAjs3vFz47ArmAS0l28GCKImtsNuS9NytoqYO
Hj3LDxWdfF2v7Fu5cHMcBI9jKhhbYPKYIoshZuvyl3CsFdyGTSgbM5KRVwqBy0PRNIurSUvw8wXF
XQu4++ZHA1P8f5k92hiIM8Ow73tXn7aF9XxH2IjmFbJ8QAOr/CFokTI/ixGdpgxNkX71wugWmsEZ
t1cidcptj/k9X20QGpopDyj/rkN7LCskPhokSL/4SZLrJTiO6LH+c9Ydh5Cs/XO7Ce9DIx5Hpmcz
NnrSQ7zrf/ODlQ9Lr4CxQFBhTX2nYOU4wtvZKa47IfO+9zwqXckLKoJV/XTmPZp1gwwN8sgo5yC4
AVD9n/6PTC2kLY5dwGuURrmYPnEVzJKrcOpVKtdAs9ecoierknpVEHU/HZ73aru8ufsn6Pz9PipF
foBaB+mssMusCUTZaekUa+92oaeLqXuTO2HLBbyMSPpVxnxhnU5xxOIV/2BtMbCxN01l8sGuk/sz
6lLJzmPQ7KTq/MC5tFr73auRopY48bntiq7hSgpVpfLlbjYfgqSth8ygK/EkPPL8vS4BjA+fmZnq
0FI8gpGnEzaNuqayy48Coa5cwbG53U4gPTIU9hx+J9WnYJ7NXr+/SAS2Ofo8rzbMWTgcxraevHAW
ZdjebiFIskwj2QJLyw+WxPELR3SJCM/EtlKN90VHXlspAWcedj4kzzjEKTDDEkJjFjXmhH8yN1q5
0Pbp2D0rqz0eRXvamynXbwJ6MaWX7+mIeUR//VGt0DFZ80s5hIxp7cLZzBxr5CpamPNLxv9UsF4S
CBkKOMNkFSLtm0kAxAPshcWZoH6gePqBEpHQONkF7kuZ0xrwia5/LPyLSDnTb51id4P4PrFx4pUu
LfAL5IgbDXlTiWy9BvgcjQ5QRJPmdwdqLUKpbYG8KNspu7UvR+DZWSD5M4xOTqe+zO+D/CqJi98R
hp2GMZ9u7WzHIYEnvpZr36v+ETcDg/wxsHCcDxxY+SNUQZV27eiSCx7yxzOdMsqNB8h4+aA7keKG
xtMpfp5KwVDO1OfNyN9Gqdc+CF0VLkTHFHLowaEKzzF0rUIvrxawTnO5dOglgM3kcpMUOxXOb0LJ
vcsiHoEO5qmYfPcDVBsMNStcfXgwuRTgU51NTjn4jktOV4AMuhvAujlVHrVxoP7Do29DflpGttwu
Vga9SDg/YJ6J1dWM75JYBcL42KObPvLm7TXj+NZkEMcKvwKeHHGRRkJCcyREt+/+1T+97EjM9h76
eIA/0Ht4VSVrUDolts1lpPfIoFWMwXESpFixNtTm0CIwRbDMeF5h1ddz7KVP6CHhZGvFf0ATqiL3
2zA3/8SERRZ3/I/8d+QoExaTtnZUChsNEA5IfstgoizEpxBOsQhUFxkzQvn5Yvucg4NM7WS7B1oU
UugYT6D4sYRp3okM8sS9caaIwx5tRoU4giwoVOX7IWjRLh7nCTprJ2/XJSbj+XcOeTCrDR3qdDIx
5iYp/dpX/CKg+jPTZY4bdl2K319uGdLTxhPSS/ddXseHFasafbkzM90PfglTL2aUPAqLrpKj8zQ8
7dXuX8cC34RO6vqj0589KdW5notEkjwTk1N89pmRyG5WAg9RPDW9r8B2IKcIvyPoCgOiweHKeCyb
jVLi3G/d6nXQjqbK2W/2w4uKwNVTe2wob9SjvSOeTBhWHFMtilGQNJZX11SCOooxY/K9CyB1eemx
8w3DK7aVzgGXNVk/VVx7wB2sr0tiZvnuoYDJDxOQSMbk33nJ6ZCDcKNb+T1AUOp6LEEtVxGyZ5Xu
7/S7YV6LfD+Y78spwQUta4Aqm9nyPo7m9sgyf/oXwBErlF18Rex9ygJew6EJLmWwJ0dcJalWa+mD
FdmhSmzzzqb3z2Qd37r0o88XzswkofOTBoT15UUw1dgBIr251UbRL5qmYvQw1POHkFnrtbEbAxqG
fDzRa+o36feVkD/xpGCZB9vXZ07/0vXC1DIn/hGs3GGHClJAayCB8mJ2p1kiShXfP5h7GxqGt1bH
s6S79dGtZwDldWvzzCxDowHuuKUsBcLMdzi03cNI/RjFGH/6z29dD6/txGI3DSjZmp+238Wy7+/I
6BeGs5zX/+/YTR0q5azUCQmYIoVLjoZwvGgDF94arcKovmlCJkFMceiBXmn5hRhuh/5YOqaF8s0/
izxAaZ/YIVFML7mBIaKjoIYOg1tUJi172JhYmZ1nJzZXp2AJLhqyCBLS41CdiNyn0UglN9DqYLPI
aBv1ZZixNYx3b8jxe7JgELuILXeEQhnIslaoarkxddTO7540AwZQRCsrHIM35Gl7nsojV2iKoqGk
wRjfSryk263WyZF7gBuWHu0a/KzKAn1hW4dIJJoDthtlq97bgBPG/j51KIBJzljvATHs4XiaR1cI
IBtdMGsXPJp+4f7IK/yk5PgXvHR+LY7v6RvLkWwcOte+jh36u78Q7FCOOukCuUz+HsQf6+NX/OR4
RftQsd5S9hGkNwncYYte9UU5Av3EvMnvKSCKOgVTMoTi5CXCpExEjPifpC1pz0MMbyg2CGsGURiZ
y+x9m3NX/MhcRikDVd8MTmCcZnkgYUFlF6sMj9cQdnxVc11m4XDyxXbDHNr+c6sq0fWLAggpAHlE
ZyHEPqpOLExwWocgEjzU90x0j01L5HVBI5hUCLlEeNfFevTG9LqHxYMUatVOdnBo8OnMuTtRYFs3
cNJZoBJohauK96wngqm0adv+HpuAs+lYFjg1u7hA0b/jm/6aMlQlfpef3dolgj8Z7eVp5VSd6Rem
IMzuZrZ2nia0PEtsWHUNAao92GUePYdvqCVvcjPT4y1hVCyrBNFLcX0s4YKnZP9HsIMpc/9Qn492
RGGGRfUz31eeQ8/EQEhlZV/5hGz9D2AZQOoMuZnuOD6twqH+WVBb0+g7GL6G8uw/F9bXefhSN/r3
II2k01qrqlxM8bXi7yrcXOJb9e+YxZEhe4jlUUQgtglA+EUSL+L6j//7zDl3C+WADZ4utVmA9D7f
TB5cvNbtfm7E+h24jybdqQ+usCkdOSaEDwwh+OrExn/4jL9vhan/lslF3E3VdUN3/sQFfS+vaK22
fY11kWhC99j87mC/hs7EfduO8W38VjyQla7DVw/N8t7iplljJ/Pyiq95/XuMlmLKm0lvPkhaRTvw
WuV1RXnojscaPHlO65yzpLaEh56y3ZiR/7fyWYzv/gOBrCcLz9F4uU2CSGmtgziVRPAPKOHSWdL0
4S6kctlLmLlo7PaLyu0ZRHjrE/4iOyThLmgiKucNU/f4dsNlUtJp0WGQujxOPH8yebtcif4h0Ot3
9TxS15CiamhBA5y0240+qQqjeUY5a4FG+k2Bb1royXwMha3HGO4JL6uwiZWUx5xwUK7Hb2aCDTmM
dRkJzbxpZseqbEtI8TBWLOOo+SHlnIA4rizk8EaAjyMgvQX1lFrCGRx480INK5rbh6FP053FLjQn
OeoPpi/YzPaKNffq3TUSrId+RF5pLolxrS+LjMx5+5XHQFRaz12FTkPISpFql2qv5Oy7q6hxGOZp
LhdJfN/5YiLC/XM7YrF8IBZ6Zy6/t8lWgm1C1I+dMV5kpzkFB8pqMVpaL5zvxoXvYW8vZnIM7AbV
sz9zZ6G9c0aJbVBLQKCahlxxvdE+jtgUxhp2IoJMsxfjNX8YDEhb9Mc+ItqBf1yhrKJLxC2G8Jdu
wa6eyjJUEeOOd5GfwbK9rnrzwW1Df7kw56Ub/2SPHxo3F/SXgp6HyqMVAjnu76YcxcFLQq15dGdW
XYZmCAuFLGbyQ+AwnXuGR2Jrz2qATIDcx5Q/fSo4pbK7m6JiQwMlti/U0mV+8bs/0Vkfy6f/JFOJ
NxUtfMiB98XL7gryyJU2Jo7I3gJAtlNxTj/udW1WnqVvpfkDgsnwkFGslmB1QFZt40ftaPMZTRt1
duqJceO/epajWolSBqpAgG9ku47Ech1g4hod+m/GucDpSpPua+I9dtYil1VjH/j1NCwoPNeDahoa
jfV1arqJ81IpwtMcDQUK0vWse2UrpyHBOMHNjeeLRISPZzuSOIfEczAZxOvF+oxBDkoX3h1e6ZOg
uXxjyUzoMrlkiHahM/GQbBsSTLbTLnGwoCb2NKVSnfrxpdmAEv2qQ1sTFEeWlOa0Kssp3nYLyZ0J
+WbbxQZ6a/m4T60So/jx/jx3vIYV7A7ROMOwL1wXiVCfDNFKBvyjNSdqGpQaVSCExRR8qh82iL+R
K/r1VORL7a2c4m8gFUlePXiWJaHmlgbRNL+0GDCZaB6R6uT0eoLjjFhEYApuJ5myzI/g893fMSin
DQ1cZVl1o3uQhcM3XtKww5MfwZOtv+pAjE1ElegMeYd/bDIeW31koC50QS0iiW68yN/xQD9sx0eR
P/LZSnxg/OgynTEYm8gLcb2LyoCDUUuS4YNEjamjYN9T/VEzEOBrX4QEs5XaOIYhk0BxNuD9+5wR
wR0XhXsQpec/ggUrsZpyuYsHv+4CmJFYxheuzyO8mIVaNyuk9rSgt9KrNl+G1rPJMFbxr1RxH68Y
sZ2ynzN6bFgUUPThcr8suxEiEftkSdoLB3Jm00MvA+s4ub3Rq+Hj7z+bHLUpSk9Lax0lfSranIXr
/VmJj7zB8HVrB5w9Bn4Vnppks0n7qvAlAYscSMco9Ubeg70VcEpYpf3tO0fZwa0j74756EHQQzxx
tDR0exykTwRGt9tPkqMN/5g4Zdg4I18RGJdYXM0K8b/mobNk7btd7P9kD1LiA7nbF/6sbGQ7Ba85
a0xc7W+HNPtZmTRBbNRQdl5spGkpj9JcNsma9yncBSZTE5hvpEabLEMzxfpNAtJKTXfJg6qomOSE
CyqPwGxN6UiNTqiYtZvB8ATEzaQag1Tj1quypUblr97R2Jnb02qaHO4VZQcRz/xPp6K54lblJSg7
4W4dLYPmyji+Sh0pGYpsKjXD8KSV1IVfzdF+UmX9Dde2ojKJqdM+jWuIXehH+s7asaHPLksvVxqw
pRVsP6+svbOdSCJ7275J8Am/oeLJIiA+/Q0PZcsJcF0XztDCPCWkxiRR5Imq6DhbEztle+aYgn49
YZuX80x0c+k6CUZpC5TQsyjSQqghPCXZSzi047Ac9VHH6aUezGI+VN4orlb9DXGRr6tIq0fvhG7v
ympEbtzLRxfT5E88Q5XwKyyuNLTawdZMLQYjZ0DRo7kFwmdIdFE1+VrB9pu1+AHeg5AsLAovp0fk
1x8QczkoaShR2UKUor0GugY4joUkD6wO1R4JVL7OuRV0DYg7QvbcVlIjTDpjYvJRx1hbbdIuUzIg
TA8hcJtUI9+jA8OvSmXOVTbG8w7Jk/nKEoimyWhv9hkH1sofMGt/O1Jbhx6S3JrY28hiccxCRkrn
8tojbqsBsNFB5sqt4YU8N7w7hbN4594nyIYNeqBCHur54FiBV8DtEQx/p2X6U1S+pLL8AMgWyFEC
xAdyJX5i2q5qDQtyeNkbyE6tIkp11eHwzOgze7fnIROFhieCIysgjttpuWTk3AnTj5xinSJWGMfF
znXdffhwIVzah1FYaFrJU+aNJ4lWe4DO8jVy1hZImThanu5ixqJ01VycglLtiLlMdnZJxgm30ed/
1P/4BB4o/ENIHNpTt1wJZ8aGOEaif+abfmmmdmK09MEKcrDN/RFJot3nJvj+hU8j2eLuXdvOs0mD
CXY5UkeH8+wGvYIspgh1Eg7qhK82uQ7opDR7rTDdMvvcsIxmVlLolp21a7v493VeY6TO3JZFVPNB
oAvgjEQ+ejYhxwaOeXDCGaKvaZ8Z1oBz//gjaRqI3fRkUGCkIvnJ/Rnpgkzp/tCpTnsDb5jXZPq9
MaL9W5u+Fb2O3GDg2rI+NurNpoVKVpMQ7SBUD0fSKMskc++vxydskAt+hOVWjgwblTdGj9xHdDsN
M9UygX/Gb6gl09idhxGydCRudqmuXOap2NpWqbw3o3eTF32AJg6GsG3H2BgMvyWCmv0RFv4/aj3r
TiUkldmXYp/NQZCExWVbomEiVwurtFNhDdiaFkqlX9fQpKRGFEMskfXbstR9JSt8fiADsZHFehjC
eO8U0Ie4Dlnp9qZN7Q3qLsyrYuEhzS7ELoluMS1O4sJSM6gSB0W/W3EcabJ8Aw8YuG3D3ggM4G2Z
1+1peyIEpgJt4hlJXKl1aGv5EmmA1IeLE/VLiZoub8rv1rrjfavgeWnSdwGui6mLIomRFwfDFDe0
z1fX086q6CMH2ziITHgjlmRovZEbeeb/N7SlR8ptxJrLT2eWvcnvAgOTyPeOqHEYgjO3ag3H1Gxw
d9mKRJqc8ypl4aJwTKt3zOJB5oy49GY7AkQ26Vpz3UR6featHX9n2pcbOC4Udhz4oB/BKylgQ0r0
DnD1yxxla94a3riiq/d1C2LW2yd+rvhGCEiHMBdWV/+0ieJbzZUQB7wkR2vzpAu6nfS/bWEwbQ+n
HhIHBNHHsQISMhlnsbDTPOL1iebUOBpl4mrxLcwtJftTqJRB25c/lWIbFGo84qlVR+Y+xu2r1Y5O
oZQxPEt8/VTCIssTciUfNXBVgmWgp/ixZ2yxJVF0KFe5D+Wsk8CYmgbaOpUc+By5LdEn+ubAcKlL
QlnSLViw5Fe2kxchpAYgM3F7GDkNlhV5rL00Nk5SjughU96ZNiriBBbxDdslDo7wTNAdujGeNYmc
BdC5FQOhgQdfUgwDeGVvJeQwXoKePorLHm49ZH7nlwUpWbqdHzJNk/KYGI4IMdauvXftnRTxVVCQ
H5w4aN77VL0Fj0NZ1HbJh9xHawZkrBfKZ9/guZasXNKaNb/aqGfGdgh+hp+edxX5vszQh0Uq9eDY
gJxguAiWSIe6WY7UNHP3kvvCOp5T64FgNG/MHtRVg11XTGy5VWdF+iuFU4G78p8blWYHpmrlUbYH
vbBKw01CYoZ5gjyNhHxpWMoqeM2GnehLM+M54UrXKFJQeA+S8kV9GMbr55/W/5fnYLe2wwc2pYsh
gCnAMz43BYTzY9it9bgV5mCbUpuV5yO27kadmxkvOT7KUXlsRdOsYTJN4wI7mGKMxvVu1jw6zFYJ
c8F+qKJw1pPj+h8E4Da++Z7ozaCwV9haTo+3XpTCx1ygxOTXJXuB38pLkL4dNPlB1Qnc39BiSZSK
QJtru1E2lJGgkpcEUD3iPYvDDKw6VEx80UVZPthcu3X81PANtxBblpIrvHvq+9iWZAszKq+sUv9/
P3M8PAntz5cAJK/h/4k7noOrSz+3RHqy9jzbEuwEplfP/Xns9TQdxj8Xbso4Ir8gQY2TdhUeto5S
bdj0TgYWFWThvTlpFIkSHm2IAXissLTwDZvVk66jo1Un9QGgxgnvLg5YGsRtsRcEgALz63Yhy4hq
2rRZ137/de1s7YvHnOa0Lv/PGShJ5zP8GzrvQ8n/c0QklPQlyQgX1vx3WAmWD3QrYO6rQgkHO0Kq
GOIMYZQIsJ3dqUFSSErts7BA5oETZe1m6OE3bBKRXA3NxGxyg8eyNMbWvM3ojRAMFDppZxCwVt2z
eE1ZoiZu+cPibmHdAK0evXnUpPLgDGZoUbimB8ZNAeksiygzAOpeezDduY8OrfUAkW+T5JTP5Oo3
H2A0WJRrfB6iVs24ahJKEIKO2QRVRmRvvmznf+2wdHbsahnPxK0GDbHDdPTqIz4foyhNgAwwV4vo
DKR3hq7axhgX3jTwWRDvqb+g+xPKNWPN3/BNkXlogGbAP2a0kzvgQJk5xdWoIhz/AjxpWMPo34sh
ZrHUJ+Dcen9/WkA2WbLX8fGxRwCa6548kpstuG9NAQPoybP/y+m9J1vG9PJvrGYOeLPArDL57kwT
2aOw/h8RABBSFXv8qsJm3rRsslAcWPerJB9emSdNQ1v16SZfUXc/L598jxo8FkPxGKWyd24BdEH/
k0oknhxTqv1N00Icy2v8irVRHijCGDsN758MNUVXMfMJE8xABgt0ZktpeTVCzcJdS0iM2OgOZhzq
W0w5Kdl4SnvonzxZKraz5f5ERkNwczF31YGI85y74KJ4r8D/KrVh1H9XaFFz9lgdQ6zN6XfQvf+H
0PzgB1PVZfUXsDL810dQJIUI/94EIB99vDabjwwcDZRt5ARdK0qUMVvpZJYYHZggMiu6iDNV1/Tc
gOSBQZLA1Cdp587ivlnLnmjmC92gl/xJOQjjriZehHMHayD6K3lZwiGImnFE0GAZFD1SDtEdQ+rF
WBkh1rq+DBDTKotTzcGDarAOcEa1vLhkg8z/dSdLusYSz1FVg/t7CgAJHxjJW8jZCS1P2KFIXPAl
nru10Id+cwu/3FWGlgpk2Dfghikr9gNZ6lVaYajcsxYWOfJxqtEAAAWKpxPx256XIi8mKrUpFTdq
GqBIGLqQDSb0QwzQfz1jkstSKldM12hEef5RM4OCjySPzK0BIrZugIWiM378yHykeUShgzQL7MJD
dH2+CtyRW57+wFXO0JxVjYXHRo7hp6EB//Hvi+nplTcoLzPJEiUvVWmaZqjBp93d4u7F7AAez/qC
swtc9olonAvhpjN2oQFTpE80OH1qEGjXgEm+EIf11xst5ksVVd3Ffw5unhnUKfjORLyTvzrx0J08
q4tXFEABGjpKKP1KAaHODqpYR6NuToMfD7fmWFJlxwh5xkLUQrsOsJDpWWnU9ZzL8b/mfCtyM5EY
UTpLqcQXOOmu0owdoiHbJUOug1ToBMEi4uIFXsxJoxOa8+BxUi9sLOhiolZk0iIATY+yJQLAL2n6
F0uPk+qWwtyLz45qDfu9xFo2kFfc1WbZoE/hQuviAeMgG6K6NYLYu7VdAujS3QQwZeUZKns9rF6d
H1D8xp9BINBlo1NWxn2E0ga7gv4YX7El+EOXLWFMFkxaOZTRFl7EkOTI3ubHgrVJ7ouge/rCMRzE
pjxJVHnVzy0jqAD8kcOgXcbSyQHHUsacoOkKeCBHYnJp46edAG8CjA9lpERCIjRxuxEQz0+3hxGD
0ammZxMUw/f5QP7dmnBh9PYbgC7URsfvr8nTa/FZ0YvlxF7PaGgtAYHR5moFipEZlaf04ymOdweT
rz2XND3rUbYLppoc4D2MKMswD+XugtCrYq+MYQ1KlKAFfxDvYuxOBVNe6AWIuxnvRpbJpszUrzTV
QLmf+9s9AJD2cq2M7x/eBY2ACvlmNPzcmvHxUmM04JBDvegELODD0945PgErpmCvtRVePysMsOPh
jYfMstj0mrSfExnda1Q9gaSYyBt0x9kFgpfgmZW1QbAd4YlPGgPryc//febgQuDl9BpY681pKYe8
/Qya0hK9NeeDhqZn0ghhegHfqOb6Hkk3c504zKKSOw1Q8sA0w8ixGxGz4JgHDX+RHUDdw5UenbAg
oqy6S+ikRfCMQ1CENBTzsMqkPhlUHjkBmfcHrOQhq0TNZ60XN5YZOavMqxeqTTepQosR4dVCQ8Oy
Yd65c0K3MWi68Jhwn5FREpjnGMVWRQ2krM8o0pfU4fS5qq4vii0wuPIqnDqjzSgD/BtzAHqIZAZa
tn4mbOnwCCZ1cRJen7KhycHlTBtHGg7NfoJgUMrklEoO2v/5smFwlfrPJYdoytLXhe/jGnOtQsp4
8oEu7FpZxC4/Ld2gnQT8o/nZm+x/sHLNgIWvewnfJOYovc4KahUSagPyPnPKzvvbLC50kKkPWXe0
z2PKGaYPf2qSWV9Y/8nw3oDcGvfu0q0AjI+FsYlFaZlTEfZHJ83nFtp9pd1R1G4aY4ISrsTdDAyY
qc8HiCb6gletOeUljhxzO1y7zl8NspMs2pwUrbIA2bhebO5ZYAa1D2jpQ7QfTasIn15g845jju2h
pUeXeFJSyntdIOnz7OWnxFc5+wBOR8NQ64CSBrVwRWMn3fuuoLjwiMC610bLuQyvsf9HpVhTv7Qe
AvY7M/cbQU5u7af6SzW7kFMp9kHUhvjm1ABq87c7Bqxu11ND5o80kvdgiHpRv7s8imjWfVTQLSon
90AnxsP9AwiyQv2L87gVG8PabRRcjDKwx0WF9Htd3QpDUuJOlwwZ0iXflI61Cg5XpULzHZImCOVB
y+yPMUV8l8/wCxPCs/4dPTNW/s4Q5mX6obo2W0l/zsqs/bX25TvR5hAaqkyrxuq4Fg8ymJZ0Ank4
/V19muAMh5YPD+OPTdvaA3Oj0JcLDgJ2jvx7ngnJn0kFVzkoBBA5bAGKzJTrV8IIz1oT5UEsssI1
lRT6MnhfUD7kdMP4aSwZx0r5Sj7OqpmILGSVex721RNK1mW2WYy99/myK+ztqEX+mwT4CvTyvzD9
fuTGR36Gnen1+mNYRSaGQlMob+cgIIpEBqVqAYP/I6UgZQ8YN9vxWcOcs/0bUSC4bXJThdbLYCDo
8Um2HCRUGQycwaD/XhEQwpGMQgdlCbRof7S+vn/f04H9OOq0T5qTF5MeEYMduE856ZK8VaI2/DU8
lsiWbCK/TlkyS5u6Dly2seYnz4ZM9uF3YTwW+XIqrV2UzHG1rBkcQ67jpl5qqGqmq774jvoyBs1Z
HmdYT0VbLk9j39EtPfCpn1Td5AnqXNd22qlO+cMm8qeh7jAOpeJQrgXd49xG1GTlr+uaBpPfXP42
X1tMuCxgtnQQzbOfVJsbcnOpWGyBtD4lyGqgu44IJ0LACZZlHINzBXp37sm1Y7gjyMKkd/BQrT13
lREGQvSgBJtPjkQhzdsVg8D/Izr5qMrW8Eens1K8TseixVEQ8D0QLI+mr064DeNP0dqRKmuh4QpV
1wvLdDtIgyVNq6a44cGOT5Ah0AHdGQkxw7DgUZVvNaPVk5wYLkKp1Ltg/gynh1onvYL+KefuulLr
3fDTOs7ma18fE4bCGn2z/MAuvX8opGNudf7Z8K6dRyCVq2oqhGeMKvRXjyAOA4BzYuVNwBpng9Pp
ko5GHEU+Ukfj0pSO0hbgwWE1OMaZUv5JvB2kI4sHYhb7r4oIgM3nLbwVfGk378N9XC5S1TEbwMWM
4ZugCGLIws11QkrS9leJPs/YUrPigdLe62hnSG2+JYt4cihTZSj7Ysn5A/IPY2413Jn2646iH4M3
pKEo+3JZdKGE3ZN+qXsjkC+1OYZfhZ6wZOURh6x2qKfNHoDOlylp1heMtbO6CLWyDOBRr/TVavnM
9IxIA7WL9Pjj3odiJMINTGta2B5u33Tp3Hvgok/Wg/Qi2ucbcfJkCnu9HK4wm4+zigpHUlU5ftb7
KMmE59rMarXucDyz6Ezl/szL52CyBo/5wku8HD7rH8HtgGXKxh+3RLgV77g7Dh9hQhGD47JW//60
cJjPZJTGZcGuCmLQnJs4WM+jTP67Bpml5j173s4iBGUF3rJ6WnECiV/l05s0R5Eu1cVN+lnOUP7p
L7sa9ZkaHHvzgmgMbNPvjwqIrTyAwH7XuGJJlCoLQe58CI6K3PEqswRHTOLJF31Pbp9cIV4UMJKu
ODbI6YfG7dyZbijI58RSVvqJOAPirMCDIute+HulRZLEjQOMSIbS7MxxQat7VqdTuj+0zSXGDdjQ
0ozEweaaVgAJn5g9U5LIKl7NAqKSsytE94b/ITpnn6VfQKkh98p20fEO4diuoCFR4orWL7V0eOvc
WEhot63ObUQ8kVZ01NWNGiKnUgUa2DYP1o6502rsgYLk3Ihc5slt+icWQw4fJkWxxld4eWfqbFXA
qwtmbXR+dwrBDtGlIhpsWNIf9E3ZdF20P1CXZL1UX1ABL1BPzLHQS+cGdO46ZSTNKzuwIQb/vO6m
VHlDj/7c5QfP9XhsYVII31aDrmFo4phRHecPs1IRsTkU/d2JsF2bUEc6lOiCnj+8aDz7/oogvX+Y
RFQeEGCb0GmOWlBuUEd0hV3vzuL/IyxABzeGb4EzM1z1ANQy28Pu/weDound3YmP2tmneKQrnhAz
YWQ+pKEM8lwdgB5/lnDzYOPYLmWRorfmxFfFyV0vrO5OQd89Xtny04L7ystIpk9qj3R4c3YxvgUw
uFGqi9gA98iI6WdsFb7tlDypUvCRXKEfY6lN6cvaqZwy5iLOHQHBfmAQalWJfjly4ko47lsjCQHW
qIxqXSMyNbDxZfnBfCKBKsU1Pi2DNhiYom45SN8NAZnqbcbVl8xxO+o3WIjzvAvsYmE7Hbh8NfoP
f8QJHGUTLnN2oLLW6H6zF97Um5yYrsuauwUMPeEMUHirOmVh7q6GGmcFajSFQpSyfssz9MaEnqA6
HL5HJrbuJ509rW5rtunWCssNlt5xb4IuS2tjLgqTANBuDrqlTD50XhdYr/8uzHsq6Dkt2jdMeNOk
qs4uWrwTZtdUZjFZH9QLWCOfbKnyLsf7rZWFkZyimcfhr0N9lnJp/BhFReibAYeI+sUL4YV7nVM/
E9zj2PvuWXFY6DUUSAbR8lPKFtm9EiF8UTdaWl+uSn7qPvY6ItvUBlWEMvuvHIHatQZyFCNpeb7t
1MWgfJ9Zb3Kjibjn+X5j91X0GeH8qUh7ZZR7FrbNeHGWO2cVeKHRfJqvhi1mobEH1x7MK8ijKb6v
jevWYXv0vWbpLsSPmNd0kQliQKluePyej3Ci3zqWhJ7YWbVmS8/PbfhteXEAf2ik/v53N8mTPxLs
G7/3k/qLS+ftx1QSOY4OxyHWvUVQtNV/vcvF/gDjemx1SjyP4ZHi3vDpj7rTbjT4cqk77hoyvv4/
2EnKNTZwS8k2h6K2KfMUjfUJgveXFgSnknrz4W8CQ4p5ic8nWxTqdCyDfVG48ki8MX1Ni4j3hKEh
l5Tq7jw0lLQDGdGIKTRgd1NlqSHn6gCLxb1PlC5XNRhauUKwIHhAElFJbW3A4RX1nqzgfBMmBl+A
81uMFgSFoJLymsTTfziCdicYvOw92Qo22mhVofD9p2OEB5jZb9uxhhPMJWF6pfbgCGxll0TBQyWN
z/Mpri5gfHfI+RGYSddM2ZWkIIECpr6ipk6v72EQit6smguziM17f8O+ps1qLgCXpNybo+CgwKRL
RT86W8p5RWh1Hn0/svt5tsq5QRbfuxFi5seCqW0/3ZdaX6NhPJbkvAgqsIfPgNbWyhUWSNQgiQKl
xYBwnx4J0roHSftIw/6rz3G0pQ6+Th1MFslGKGr7NbeBSiXLx+PmWsZIhGpRW7rgPihakykPVhVK
fDaYLDPoXB7d7HIyXfnkd8IzXWVoJeaBbzcnGYMmJG5wWVxbfK6bUAkXySK1DevuY9y1BQ0rbiFJ
YwRcny1v+ystEAqFd3uoFGKzqvuc5VDSBXoA4SzNzc/8dI1Fafjn7+b2dd6w1Esyx9x9zSY6+HIC
W3qYSDUXMfsfWf/MzkV+uCJ87eTyCw7tm/SOJd2FjnSufwnyYDR1fu8qz7E9fSf3PBaI5EU3fsTN
7wi9NHmEbpiGBj9Hy+dp7krNIb4ItooCqPW3D+qWJbAYvYaq9dhbUkb49g++B7HfMOT4A+0RnFGP
kgGQma4erDbrm6OS7Hv2LCy+zRXM6Vu+0q3bVS5Yxdjv/q+oiObikTGU//sSlqOi38NmfT/0Nd3v
GtT5rEno9qm8eD7a/WMlzwbZMV8tbMktkhMuM89PcjcpuxlxaHUNLSbil410+p0NSbhsGEgIb2pl
WtI5NfIsETfbXTxt74VIzufU0jZYp9ZI4vmzc6u34PLmpHxiB2X3BO/W1Ym7jMJOkSEjdi92gQSQ
dQ08niLM0YHPZaGT/WsxN5rdMhZKfBV4UcktfSLKl7Xh2CrgavXWKg1rKHez9LENTqPXGOPpbOZ9
JczkjFbBwISOGgCfKr+6sG10g1qSDjrD5/qePhbEAf+ICpu24DvBQILxs39AEG/AA6LnIID/8PAo
54F+M/pp5ui18sSPsJii27v3yQk+G+VA6C/r7aHVqhHWBQQ/8s8Bx1E6tWH4Ii2r9/BkwMaWP7O0
A3y/Y1WrRfXykv78KJ7jnaQEw4rZByBCTgtV/SbVPdaXFf5UAjAf07gap4CsREas5DpZzq92L81a
b5wM4GXVxU4PmSyQnrauNrcaJo5D+CE8Di5cDIOFZ7Y+RSiypEfl/d9bIOED9SfFvJzM3QKjiJ9o
kOb3fjUqg5OYxMaTiPE3rztExbE+ietjiUEjdC2nNwyYg8Jwf83gFTTXH8LuudqIVkvgdb3x/cSe
tfb0r9oWA5Q3GzNuiSSJqt5z4vmqtzOVQipUZTfWHGCtTANEYoZOvzIZ6xlgvE2o3Q8A2GHXq4Uu
yYfO+U7SpByH8A5Wvu0Le+9VT3roMWu63qtPLpf68LzY0xPB+lVT6U+HMyuGDw8E66QvnDSldbxd
3yIJvBZJsqWFvKuvZ25sSEygj9I7Nrt2i7tOPkTLsUYcdf8Gr8bx0U/Kjxf21XGIyobZqeaEjX4U
usz5xocM4ZMSWR6FJ5zRpu0YWGReNDXG1EGtcMo1eo4q3ZIOGMaU77bNGGaJypJLsP30fADttqT9
RrR4YmWAPFhlL6sCPZ2qIDdMHf2IJRIjD6EgIqOgL0IT22URTshtx0m0UBL1QopKzj32J/XHxPX1
Kr4/HrlcqDUyhI8pnna/3U9aPZG5+SU3X0Q7EzzG5cv3PEMgZvsW9XPFfQEp83U4LSNH0ZO3b3w9
pNsBuz7m/mg3rV+sPvFSEvCwSkUuzcogorcS86ZkHWDTwJcGRtY2w5XlRTGNVy3vVf+FRXLjxz92
ZvLLaTHypu/aEtVNS9Pf9hVdh7vcLmp1n92iJrr1L4VIqdr9/QAbsbY4ADNL/DTMO39TV9LRkWxD
LqjrqM2a/5OOs40MCFeI0sdw+lC8U3UHng4mEU6xWkSYxOWcj/MEkgr4/aDTg+W1tfUp9dMjdwLF
mNFcU+kcu/wHme9HomT+IOE4WG+BxI4ax7nJnmLa9cIMtS3oYn6gLBGd7wR8fPTIj/hW7T/bIhhW
iu5zQtVvyBbvM4Tp3Vid+EAx6Co+pC88UGTXX7b1bNQY35Ee3Gsige5O8Q4EdlVuNXHXUAd7hy0T
V2h8X/FzWZTBq9J6odd6B7z/QnYBxlC3wHcBxCicpVtufx6BRJz988CMHSwdTueNOVSbP+QyhV1f
slVovTXES/EooLkoI8640H1ZHtRaweCiXlXgMcdCorW6aTKP2sGHAvJcG1gZ6/ewDjSDGtg8UT8V
kkXcGtoGoryXPfJxuEjxjtowIro/iqOANPEeWWVrrm0Az3C9fCoTGWt4UoT+faisDry/omTW09QE
3Cf6EkPvOl514hRwr3GWauz0nFjmiI3XEctwCKtFckyIRqG4uM+ujeKO4Ox4aREG9uRp7FCOvQ1S
g3r4f0WTzEiIXTO/FzEUfv7DWq/6ITIGACsstB5YcapxnfdVMWUxdTQjfcsoHiRboN28r9Q4LUzE
kzhHHOwJAfm2/VZ56aoLae4Flvd0mSfighryMalBiPqOPeHcnpgM3CtH9ZyFs47YqJn7EUXF0mRD
hNAtuJ4wjeFMsv1uvxFUwPbckcr80ZvIpTCfaiQkRr/frZ1sEF4LW9NP4VIjVehFJ2gnJi1l0wx1
NXbO/eSjsIJU6T8pGi5kJuf2m0KvKQK6INk935C3MQ1ra5W0tuIXeK+OcTIFA3nz7DoTFSyuKrZj
ZYNO7188rfaetkXj6IRSHjSvt2DzJn21NPf7JUoIBfi1l+iOScNBPwLoSRcXB7gkrjkLkHQofYc/
Q7tRmHe/ElcyJ+E/NGLIgfabQ8+NeVA6c6XcbC+wcOcW35kap/HcWwf1Eg2kujXzUmIRKvXxtGT3
TaVQu9Oa+O364aXUKD5rO8gJZ7xzOqUy7syCknEnsbE5DMSE6C+p1+UGb8TjV1nZm12iMZBwVLy7
IzhJ+t6WQolNFlAdMLywoAlojKXw68B1+ad2/nix/uLMr53N8uBdRTZ45nad1E6lbWmz27W5jb8l
+AzBS7ODfExogJEHfXrOCNbp0wHcDViwggxQ1G6/wT4LRjvuKQg7UNsKaUn6RDXqJcaL935DfzQt
Wivz7tubTe8JCcl0q9AJFWBRu5bjwgCgLf3fpWvBns/nSolL188QL+n0hxrtspE1ntDOpgDqc1qC
MbDwN4Y8F/M3D6zvHI3BzIamhkpeWDwM9lKONhlUp40a01fQjZD5QKvy4zSze1pSjvhnxIHyP3pt
PJmNtTdAvgylsF3JqLsQ6OWnGkyn8UXzOdablFTTy42jfhBjhLTIzvVQLFp57/O1gX0brjt4E2yY
ebHoxqZaXhXzK81ZaW0RdJzW5k31VleNhc7X1QnvDNOyq23M9lEFSXIz4i3gR+lv4Yy0elj/2tMm
a3QzKsHitZRyfTuer8LfXA+J9cZo88GlJKiemVWdqkvcZWNj7SL9JXS6RxPDmRi3Q0rGreqAOWBs
nNMv0tuXJWTrif3QtXB0c7i2xJnVW2YukbpCqyXBXCehuZ5cdAhPdTmbt1eih8Fn+00jBPGJyuTE
s02GqujsD8DDgHhrZgvczsWMoV2KQMH/H1xsUJSphCrTX9qtGJ4CnXGkYraLm1qdXznHCiIRkDjU
EMugxCCK+iDBZhSCPbYpwfN1yME4J4wua0WsXrBbjUwYQi0+akhEWZ1QVIBZGKd/qtahSeNSCej5
Hi3DPGZscrYL9+uAH8QJg0CdjovJKhpjlK8l281mQWNivq7J3S7ZczLILlcHDj4Ef/0Hg21ccBdE
PxugbMKcuQmFxfzhd236KSDDiJQlqFHfTOOjX7L/9NM45bHI/p8AvKPQqL6AutIXOYljh//iN47v
dy8l/YcpDW2djlUZhU8guwNtM+YEuAj+550J0fncnCvHqyoYnp3WuZwwm+BDKodnrNWwrbfWd/3h
Ei/eezn7BN/izbvaxKGjCMot37jfYg4mfnnlDniKtGLk06aLpSV6F8SujQFFiHWl2kL8U4X23z9l
x35grZ5fDvaVZ4kW3beiO7Kdnr2x957gz1I2fa6Pn4p9NnwRYh2/Ps+TtGMXSDbq7kxusCxTgbPC
LFIEaOobywTcFOA4tF6zfd6TP7stflMfhLxhzTmp8Hc5aKzOHzhW2fWLG/h/1BOADroeevRq35vz
S3+zPAlgWa3NrmBP1MQ0nbuaiFkH7FSrc0n9xKSyGMZgSkHJoEfiFgzo3DzsyIxqbd/KOoABfsO1
bpM0itf4w1InGrKWQhvYAxgvdf4DJW4DP5Jxvzd5NZ6KwQiXFD4L3fyEt/Kb4E8p9yd4Sa8Srytq
GEmMZIIzPZjEPvSGGBD71n83te/jUmhibGmLC013aqvLpl9EjBwkrj0jSlVpQ5yaBGIuP5jqYup0
eqSkym0PZcVEaeuDUkVIP1XY0DylaVqnfTvP5YneW9qLXYe9Y6bM9oBj6dh8KUJWJn8bnnaw2Ccg
Dpl5Ed/oB7pEkydANYjdBjtzADKlgOoJydTo7wV42virWwmtk8qlHaPqLfkPpk3UCh6H2ck1IBLO
mKQYNwm+JtRYdvmyN40C8yBbiHER2kxmBx20arf/BgAI/mv30g1b9b7cya0cPBBWTe+lV/+rNd0+
4XENUzu2it0Q7QHmqjHcxUSjo99A0+V0FapGbowhWGCKzOiGBdM4AbiLJCKj8lBbof5OYL5rVGjs
qeSkwe/d0TMBpPKT5KCw7QC3gwhvoSD4ShKXi+6HTRg4IXcc82dzRk6mk/puTMZeau2ezNRV8vec
2i1w5XFIID+cR1F0rDyAGynQcCrp+dgjZZroMX5GFp3ERp66X5drslom5GtBEGwj0wgVCAl12lzo
eu+A8tJfLCoNQRoi5RqW9BnEFhOghRsVxGZ85foUCTMxtIrFHfVPtsWIDeLCR8lBCECz6+th7a4u
Nwv8lMUlf2CQ3kjyJ0L6XY3NURDKjW6UPThdC8n1iwSO31yXdlcayWmZo8hoS0GOAORkaiLC+4XE
UgUr/txnZn1TRGpR1jYab8iO1kVrNy0KWwXscf5htXHR0YcsTO2BwEkOajqaT2OC3kyyOfunmRRN
kYxpSa9ymzjbuEV8J+5vVr1lzcBBRqzCSTug+YirxSiUQOMaoj9YExvXL/ujxjZ54hiKClCIWY6e
R9yZAmw0PZrg/gJJKYZhP+93bU5eCacp/w/8Uh2gwFGrkQpx/UKDgwfhYQSR4C+i3l4WRy+YkSAj
EYnuL+oQOMJKClh7GtLZS/pzv3Naiz8kDrkCrXJuS2U1ad2gJiev0x/+lqdNoMmnM4E9Og0Uq9c2
5IXkwJFKQCyiosBZfUdiI8BEzyK0bcu9FgRVlx1njtjOcXPRVkedTxP6JpCjdtVyqI0Zclk3hk6L
TgHrGjJHwGPpJTLtiUVbjHT/CZM1KQjuUNcUHDm619/ipGSVMbUZZvMQ7e0jJabFqpyGRfz4RyG+
9DLkteti8ZFY3aOZCMVSCiKw5myGd+BnyfypJ4JcFzAGTBR3GHmG5aIsmRFDiimeuJxNN0j518NF
t4xH2NMR+MT71QaMU6LVt8xwG7nmoO/BF0N6vGGSoOeOZWACLbgpsllQmGegc7y1uPyzbUfdkpZg
SKAVnYc9oblhjv9DORToIcQLJrl5u0UODiZrZX8ZTbujFlIkha591RrfNyuvscrq6bMdrQcA3xIt
nwuECQIYutypml1+pzs4v2yO3xmIs6Xg+XfuLQHgPLHauWfBODi5FMuEBDvao31ve6KvmSh36epP
yc/cHlXtC9PKEvY/fOuRMBGEIoJCVhVVrQjXxCIaGZbNBJLDV2mIiVcn34YUHNzJDq9Z4e3+OHwm
dul/yutGok20DEp00xjqgkDB/B8FYjP3/PBx9jNet0DJhrzSszgOjCRyw+feH51LyLL5poLb4npa
6nImhQwFNEcqJwpfamslkiU3t6GfjLUNsYlFcpgq42zsArekUWLIfYbnwCNZ+d4YBn7sNQ88YeXZ
ymVWoXIftiUI/Q+SgtqhUEnwkMfjFOM8Tx9vStouB0TFLZfx9lye4UG3ABunW8yIyN8u0AEnH8Gw
LgipaD7BihmInUBSh0PByaNe6iWwA1pd+a4dljp7gURo3/X1oadz3Gb734NAPvSlDJvV+xKNEq77
89F6+g/rdtU2rbo8yKZlph+JuSczDS0SReJiDwS6h2RBMqaoBYWRM8heHWxQU4nw6tkn24P+dOYi
V7iSJYvKCCqXZlYUOcK7G54jFaR0sxarxdQ7VMkqZx8FKqHtFvxkfaGSLh1YM23u/iOU7+erSTDD
ZtrvtgpYXRZOkyZDf7ertWHYvByxamAhJX/uLbIi6e4wdbiWWQ2qkbGTaaaa4wKlCuhjbbqhVcOM
LFkmY11d8zEP6Xw+svGIYG2Xweo/ovpF6EbPVOVxx9Mxpv+ItJbf0crkl1xgIcvlIFftnzOsWf7f
CN7qnnEhRgBCQh7Y8PER9uAHyTxMAlvZ7vQAopsQ6Y/rQFF8vhVjXeIzLCkabjaNf4LE11wOrKqm
wXDL1RpBfeihPROxM0jbiUQJ37Uu2Lw7Ncz08ZSGfSHOauwnwwvNzH8WpCHQvApEqjQoWSq71zf+
3RFJgYgB9nbQhcdFxX5jO9zR4E8FdLtVyEih6PxJmQOWFg2Zbrm0qjcnJHYTM+73VFlomI4Xu3V9
7S8Py/kzKgTq0Fa+5RHfHd7lfbwZULBzuC/QAeUaiWXFM3DvaTuoYL1u8U2EDxo/WLEEaWCZkltV
HyGNGgaK233q+KPE6Aa0IHJJnDrcNbyKYUmVVQtV/vQKoNIleOoAzN/FXPgbu9gUH3EaMufsNsaI
pLbAQ7zliyfklJBplpAQrbG6gYO8eO4vWHNsPXBEaJjBsGCwA3jHwh3Sdj6/m6tsB1+C/HlNVwBn
pNm7daMGW/7j+e7i1jLtPc+Nu6/J4ckU05L3+x922zP3Mw6csfjM/JnKiuApWCkV4Y27RigOjdGM
aHmHc6xqfr8euqsO2heYfWxRv67aW/dan/PkQQDUdaCBmFabdytrdlVNDMwA/BxGb00GxSdxHk+r
Ktr5xuPq+nSrbbQ/xiIPZHbkfBU3rH1xEwBH/Zw/5gdgUKljGFrNR6BQ/fhN9tD9lOJsHFc/KG7O
MNWiaJVJaCLBVpor5rVd9j/TdbZluejgdKuHz4Eicze5apZLkf0R/k2VaPPV5jEgOtYAiz0nW7Z7
H5tM9YOV9mh5CKLNMJgtwTVlUmNblNv/uWuBSXUzweFhvM4/yM+KgExMhmT35K/0LSSC0VLaoE6l
+//W+VRaxFhHWo5MMFiQgvmQtlbyuqp3M6PYT4fAEmQg12BfjvSwj+95PK5Zy1xG2y7SgmvxMdxS
pRpa71Bs0YyWopQTx4uKaxp9cPfw3tgc7ih6AsHtSNS35ehrdDM4C52X+5TxzwDeE9Y+0JrPbIeG
qIhsu81ZCKiG2XL/7tq6x4FPsnoSROFTI0vCpDecZ/HswZY8FzwmzTZfS3qeNcgKivkZISyHlPeH
rID82hAh7RU5XTuVvmlujsECdW1fP+0Fpi0kHTD+KMUsiYdvfnCSXMeScJs5GwhlV7VHY5rEgSqu
rCQPzRYeHpfhyqBy9LnSO6fnD/7Kmkd/6wVIy0nJqjM3fa5WpSmUP+u4DXWTGNxaw4rHXji2VIep
57pUi6GODCd6YxCu5t7NeJW6/sGtyqMwPixIfMIxiRTETexo1xEHAIUJrCT2+92ph4GFjuMAW8oZ
4/b1GqlMUnnw/XV4d0hfQgj8QBXk77GGgPchG4pa8zt83BGbFmUJ/U9vmgxkXgYRoO5zDpdL+WRr
AhaEC1sC7qDvbwwgZNkhcGXrgtpbIoemBAZulLtXEShgvu2azrTpCwLWgjDdvPbJCaE0RVVpMiEG
n3kP03Kj0tEZvKQI5oE1WKwrMz9enq8GTgJK70Wm0SBkXr+hS0pqo9279H9QtcpBJque8+vdjX/Z
iGymmkb1az7eLljpRmibqrJBvuWM2VzsSMKnvy/Oq9IIsqljbAw0Zs5XA7vnQ7lsGKM45K414KHe
Q2KzZ0R+W95mD5MIUnOkZh1S2FDj3bMzFKY9cXN7f9dtMP4ZWjxTIaaJVuYeaErkN10lDs/kov/H
Fr00QgxqvvGvNktyq0CK2LXPp58ZfI/zsR2l8meoIQCfEAN5e2EK8Nx0E+B9GztZPyklUqMv7FjF
JXsAMqWMtlBVpa731iW4X3p2JBb34Rr+3vNV8DaflyEuYCB16di53A6gRi6xYD74r1s0HLLR2bdB
7/IdPq98h7G/syegHp8O68EFM42FRQN6yL9IFxKSler1uG9y7tje6dvjvv0eN5jF5iVfs86ZsD0O
MSxVKdWlu/FuNtRYj10E9fvdFf1pIfOt+QpZGn/Wut+CAbKKqLjrx3MXWsA7LuT9Uv0CFb8uIGdr
H/e9L6cwxcWct3/TK+VvFj1cdN5Ssx3OCr+qpFcxzYGGgaSxBOkrRdyaItIcQ1jUjM2dQHQNWKzk
+iSSJBEHREv5Szyv7EOxkcmaq/oy7wgtD7lmx/mGkJvkJ+hhwlIFWVnkpCpTdA2qgJonsJv5VocW
p6qm2gPnYu5QGq+T+CyfV0KwI40VUC2hB0LSIUqB56S8FKlrhMuXbOvbMRIXDZ0HP/vUfxiSokvu
2BaLTD9l7RLqiiAB7cqXijOb2MANQMBoA7eY5PPBaI+NQaELQtthgtqdcuoaM+4L4lmHNPPukXCl
Uhw7VSDZ2R5DLBc+4Mia+po2EwXUJitzg1CPjqoWkF3eJRehjTzzXaNxc+RN9BmlcX0iqpl3BRhx
7zz5gncstfqcPUXEI5TZuIS6Na4WrsEtogHPzMKyGejODH+MryOonYOpyfPKbPiekYfMCpOCytI3
h3IpV52N3XGhpmVV3fILbF8qcoC+L6Zzn5H748RX2jP15l2fouCPMWMesYInePybqXJXIMRt9NhY
nKsvq2ahGzsVUcREbL1oCxs+xdSsdmz/BoU32IGxIbxVADVzg1twlb0RH6vRSIr06aEKqbV5uYjz
NityoeoMe10FeBLFZkqEllGO9FOOcQ2F7wwLDJmnera8EF4v475b/esTIxCU3M57o47jos5Y/VP3
aaRjZNdK5iD3Bad6Idf0k9mCCij9JxAp4bLI+0EMzrrYMz7cAypz5irge/M03yIvwFi4ajUrY6BL
CZgtA4YdRIIzCipI/1OdoKNK4VMjbHFxflGqjj6O5pUGQU7AlZHR6ZZU8d86tfsiwhdmsGZnRnSr
GX2pEXSLqoSHPgLycrNl5g7jkTv/Xa3e5Ilyx7VX+krfIdZ/zDAXisyiUMKJd9Zo+g4quYUpteXJ
vMEY0Sa0ZokJtHfQdFhfEzw2hgwmgMYykXkxWh8uPy0O0RMNPEnddjl+m1A90ohxj0jyLq+cNiR6
R+AiG26T8M7uDqzvPNkeMcrTCpJHlyqDbMlZG0LBOZ/lAAqu0ls/MMpY78Ni81JMsgemri0MYTRQ
9a2DTK0P1dtusgDAme6T0AnYwn9e2DBTuawOZAxduFeH8Z9A9LWz0Qi6ARofJZUicVDXu8oghbFE
yZq9vjCFTy46UcMqsbNJWErqzWBFpVXbXpfhOlywDT12yy90ShBO+wFXRFZUrWhYCakKp6GspZd2
eisW5K0iJrQjqR/d+mberhuRMeynxp7HIUWtRm93kaK8V6D7U1fUfm1TdFuCE9wRfnUHvmFAhOr1
Vrpwkp1jI83WViQ8ycBnDAa4ZcmoWQiZyX6p25/tBAzfyo2oq2vQNAGZ3S4mIkgoV1DklULziWah
nGoHY/xjk0qFurA6xvCZPFhxW/++QBCAPXfehyF9WVu7bzzQpgSd6qeQAEi8aQPK9qs0wqPKbXx0
EHoYvrGXRPynFxJY73APrDAx//PD/m9w6qrTWPCs97arb6chVnlDHFK9fDfCWy56AsOOItZckMUZ
Q/W/LP/zFvNuNlwpDZcjInU7/uA4ld92lDXrfYTWdglM9gWSY3Cq21TXs2qiH1n7/TiOF+jhH6Oj
ssbx72ML3Z3uvql0KM0W3asQYxbf85gshLEo9Aem1R1STHGHiH7fJLibDcoGugnzk7lxHm1HIjV7
lTYFRuMHLEXIFMB7eP0CRLYVEGOQd5BVMWLfpjCNx3Z92QX0382qQtUWJDNMaBc3lIc8XWpmOkOy
Eh0Y7bnf0YlCEVVlYqwN1cIT+qASJrCVfunsfLQ+xFmNL5hRCbjgEUej2BirQDS7R3zxeitbuCb1
9W46ooP3MSC7EKGy5uix/RZqoe1b325pxaEAfGsMwX9/GDg8l7lBnEuUV9NnZuHb8PG3Hw+pbkGc
HmdJNIFsKDDjFt3ZLv3J7fnkNnLUXkf7ptXc+Zz4OKF8QPagLxWa4a4LyBAFoKgAf02E8V8uAL9N
mK9SboTUiF2w1/UBVuAqW2ts6X6xWiiAxE7WFBU7MGfYP8becT+dEpuU2daUPSW/quA9uiEAwBEe
fmZeWewFYONq+WAjUbsbyQB6GylIeaRND8t8m83bLpPPetFbmkix73odpwe6XzyUMnPIYuzzve4E
ygzwfCgNoQitVMWLRM7ESaGOy61lvEw76LIgDpnCVYUehDvjjRGXgtWAuoTO1EqbkDyxzi0odgaV
G6kHniteQm3boT7MELbYStk/bU+Khubi+xTpkdDH0LDkz8WrKK0+N0Z/eWqr8hLePSdEaNnGZT9X
ItIzLTEtCdXrJ7M90K45Nf7EXgcb6evB/0/NrlPLzgSWcIgEOeJUhMpS3rAd7IrWHtxvqk2dmP4B
TfMw2lEz8J0MmlafsHtElVDsjs4oK9Rpx36X8Hd+wZe3oqZvRd2/+6e3Opto+Z5EF19U1sFuJRtn
vI+MRgWFjqtxFakCVTRO2XuhlQLjP9dQw4AQpKq1d+dBdpenhtuCQlA//rLEYtKqK2lxrOd8vqpn
zIX/EgrQKj9pE3DYMFuf8BrNwh1atEqmCEMFZf9zc8TpaXXaGmLvAEFh/MHeBvOGJyZ6dhs0Mz94
o0t136sZbutuB1V5A+hFKTmzh2ubPhEfWFnID4wV9hD5kzDaIhG/tHhuQayDeGPaEJLbaTUu5ukf
OOTRfWR0tYCoeJHpzGw+Rp3s+WElGxyLs/ogJKJvDAV9ZrTl0wNKrPPQ0L9PzQvEdpgLCNN8/vmC
NYKwUTEw8nfEFAjrEZCr3h/SffAy2h0+o9/mXLFOO+BAr+Nkzn7je7XjK6Yo7CI71gEVhrVCzmGd
fL8cznD1UvtfWGjxmnX2lUKF3HnpLLKUKJJsMC2YzwCXaeJHslPN2sQWl20p+IZpjozifDQBFgl+
O4PArLYxAMsUUfAYBjNxe0Ak96YkmSKjcRST3NvwF5HM+9DhG9OEIN90pOZJt973/yz8LkmOGpkm
td34IFZRec3sUXydfq9YT9zJu6YOWBtizs7Ytv8+7c9H5bpDgHXJC80TU92skHpfu4D0LcnqMyKP
GLbReVWVu7wKWYb5OoliAA3Loey/rk354R577EKQ3BJ+nyxgzaz8/ziXbfo9c0VI+IN9V663WeGH
66Nix4fLgxsCCCG1JVhGmOjm0x9YFc9/rIsvesl9i0J8I14Osxs6jQPV/ZonSd/w1fG1D4OAwAcl
L2TLO0lESvaxvLo2uzE6CWYCyG+n/ppqdRnPv8WFQ3/0OOO+ZvOpxXJdwU3zhqsycVC+SfisF6ZI
uWEVo6perXawfvZvnYnJ9rMtPTfsYp2L0lVtE3zScwmtgerV7Ht3faxpIFQQ59nJrlE9msvFXLcY
u/4ATuWw3NJ2EiRef8mQinYbsQYXyHertHGzX6AsiH/ys0GcjgIbW4+2ymk9PCcUSPk2VMAyUq9o
oxgX5tpglTWXm2cSh9EEr8fXqWMVz5wbNWLRjxpIefcyFNZ4f9tCQwLkISydqG6qMDCG0YAtiSwK
bZGcihEtN7QepFFPB+HndzRNh3FFw0PRkLexyGdV4yaPUWqlQ686KeYFLVjddCiczjVpumlye2+X
brvBhp0epNpEw7RLP1NEYOWUFlXbmAwPNcQBFPXWJlb3YwXhO5nWqD6uznMYQocOa7wxsQn2EqBI
u86R5fhU7a3Ybtu/wFHVNTKhj/uO2h0Ru0VZbnzF8nIka1i7wYgbSH19/FLfKGiVR5WuKQ+41VLS
O2l5gHXav2K6nQX9+p6TuGEkqfP01voNjSryoECcSbVIzYG0P3PKl3HJEu+pWXFBSmDQqu1tOFqy
CUaEFgdqPobgCRUQLnFhXG7SMqdnivZuwo9suR9YE0Oor7Fo3gwZmYeU2NE9C8bti+lgHhZKovt3
8I/r1knCD19eD+cC/CHH8f96uJKSV7NALKk8nFT0ltrBwBn7tyiY7I2m0ilfXkgrD0e31YOjydP3
4CjUfR5ZTK0kP6Y5IuEirkMXHZ5n4VWonNRFsbed6NoFNwSAwS30QL9JVoe3t7lG+85bOIu9f3+H
Pv6sx7YoIucKw6tSntjT/G16cAjzh3ObUTYkQDD5IBEHm5c0z7Q/m1ZvZIKfpPk4j+g/yN1aNJoq
6jenRbtQHwgN+mDK51UtsxPM+mBb3V+7/dcnp0ZxRe0l+h9JDzmnbUzrdGZMY3OV6jrsk8ah9Emt
LH0FhnVPxzO2Pze3ttW9eYrtI7/amcSlW5PZ/PHtHV78zgpKKiWAQWRcRWqtPC7KmCg9hq9fpEHx
flG8I/H1y1weAwjh7suVkdbkr/yGU2qgPpk7w79uvrg4VSNGasoI3kUasnJU8jlMmw/7wgGFIHzI
/A2Ib3eiVpQ/hjNtcbZxhc8/T3mSCvSNuHBWT3tavKFd11QQdN7GD8FCUGJILxV69fTh82Xrwn9X
abSDdzfW7Mwkk28U4en8SA5UuTkRNdZQf1PLp//pxCSvXjHJHYEiVGblPOg6iNh2FGrAUfJsJxyh
O/YF0T8xC7O+u4XkFCj6rNxWNvcuMdtaVC2WWWNf+XksyGzfTiDAipATM8uEnP6auza/JPscH93B
3AYOUhrOnS26dqJb32RAgRBGpa9dv4lcmmGl7ey2aXFmGBd2OjgXoABivTNjYO4qYTnAT/xusm7k
3+DF3o2Gh3q6u5TALc7KkrrP9BqGAXqAGEy1+3aVMBCZQd/GRfYSBkKkYtiZhhR1j+dV7xCI0CQ3
FsN0aXKSKMUTTsyddXfbRCum+7061Qo8cQS/MikxbpgqSdJQMDr65WwM3CJaBkKubtkKKHbPAm1Z
kyh9PO9eWZAGr8db8Vr/AK2f6Fe+a2BdaDDkmaaKAyx9e82pmS7/Ou+zLGVKreR3srxaQAwwqC+6
P3n3mlFxTuruCC2wC5LA9YVrhojyI74YKKMyOKPmRgbdi22EuOqG6SRNdpkdZvhlsucWZrLnPGbT
cmaWOqEnLdE0jABbfRtTfkBEw49w+SNAobtLVvHnSDsls/xfT07qBSXw0qROFBc0HhQZGa6lRJdO
8J3i3WntL4uJrpu6ZwdgfhFFgnsFXP3KyRgSxrU7ROeBDayyCiq4us0Xk73mWeWVRwYISECV80yl
uIfPfOuS95PHfu5VL/643Hq8jc0a1npau93iaOwGhep195Z1o4puZzrZA6KFkkAHauS2g4hF8EFG
B4tON4DlV8I7R8dOEapsUSiBink+sKb3wDIY+LlP1V42/Grac92SFDx3fP0jaQhnwh3O8dQe0bWS
Itqx6xMO2xlWqqgOe6wbxlUbPHjyNK7wGG7a/X4jXdAAx7CDwDMzV7dscKCQbh/EiW7ES4CPrKX+
otxDcQ0WfTP66pyJVJu941PQ63MClAqgo4M/bn1uFlRocAzRb3sf8C/y3/7ceMtarl8jGxCgE/oC
Oqg4BW22bffOljx8JKbZPGuQVRsSUQ3pbT0W4PK7CxFFLXIhK4Vbfm66dYX42dpXp05a8vK+YN5e
iW9ppaYQ+mezn0voGg1D1aFAFXiiL6xNp2k9/MjQ9x44dvAsujDNnnItVEE7X39CFR9d0bbHcLBI
g3DXN0k6DHLaVi65kwnwsSOJBVbx5Z2dg4b0QvVMHn79hySUM4CDFK+rGgBw6XRBCAaAFWPeG1F1
vX8cSFW7R5MOAsewROutvWL9xaAiBgafDKDoQ+nuulukdYnFA6UKxUUtCU8MvuWY+cSl5JwaSauv
QCngjE910KyCgXk8VVf862WTIw0l4gd5lRFfXZfh8HjvKZd2heuf729zXOAcXYNx/RMOTWNKpKFi
G6NBkQXoC5TCSwxp/UTQvkj4sm1zRUh4NvHkTTOOT+aBaNZOyn2/wHB79nBAqpxKJvmwaKgkPPU9
D8Ocsa9KPp8IHFFQkBMHTNQDY1Vtri6VLFLqJaG9e3a0Iv/rJzmmgKoUUXGbFh0GKiFMiO/NhWZK
k5QSEUsYr933jmdtwu14RKow7XAHTMYcDx7dc7dXoneGI2yUwHd1Oskpn6FDfpvfxrPyUlJVTUtN
1ZKk7PCEoG1YS41H62TS0i0HKyd1uIHxVJ2XRRZoS+DXEqeWGx9o4sxzhmfD2xDzfnUI3+iH9q3y
BxuS+tv44/8QBNFI7SuUkN1pnhrogj7JtGPlnsc7fNMzj8pM5zyL1bxVUva4IpSZe8TPanynWOU5
8GKysR65MbQOpvk7O6BaxPfaIzCZe1kSClmrIQNPAhW7rn5aT6uMeUJHeTo7hO/Lu7B0SNo6NhG5
zmNJAaVNdj7qkX/wsx9LznvVIf0S586jOFTt02kTnoBFcnORoZWiOlM/E2unynCt0TQE83fFX9uC
Yy91U0H8J0X3CuenX5f4d+bgnUu03Qk938TfPxHpY806nOUHR77biuCpbUKQKTLWrI0UZyMqdi6T
c1asjB9oWoiies0l9fxbZkjgMNGa26sgZ4eftSeIyO5/mfLYpPwN/T3TgU0rBEe0TK1ZfuGyD7IC
/S9WCKwjI8Zs9cKOuPRpFqgmQjoxl+AXxHhGXlwM4u4Xu80YXC5yPfABjt1ofykUuk7z4yA2snfb
Mz8/ni5VpGOKVr7hBUvRdvqIOmSmkIOcJAWoz4AUqSs5ltqX7+kNSX26GVFr3zoqmJkpPQzfS/Ow
+/m6qOjS/Ux8p7tv4Dln4Vr7H9cSPS7M1eCgogiLLgSj9MdXD0205TVEYKHkTidHcXZGKmS9AYCR
rhwsIAugra1ePWU1d4YRfHUfVT3mtmuAfv7kpJGS0bZjI89WyK/IkbXQLSD5/VbNfhjq0WV56OJt
ORuWZuuDbxJSKfex6tKeXaDChqmItYGCaTDbywBoJH1fgINmHfUP//yIih1CbOmVMdstf4TDEZbP
5FW/O91C69Oac6zMOZITSkF2E4W4vPQ9AfW/eg73fFHh06tLhM05aQD1QnsRCwvwEJMzIwo3H1/k
/nMFtFku+d73u3ukJT1I7xUKMuPdoxi7oWHwawOLKHd4u95M8d11VOCtGrOJuq30wtkFbkAzMOdj
YQFfJhqqNfvpI4RYIQsRTspShApmYXiu+HKP0bf8u0f5KPY/b5FIaLBcfffAGMKQHdkoGaSKr98S
nQZqpssaKboHWYcTYiyrkR1qEduMB1tgmkOmOb9c/dMIrqSJWP+1pReN/W3sP2C/dulqk5kSvpJh
gh4S9HwLgtbqkeQ2JcqczwPvlIKCPnlfsL1JJDlXirsKxixz+wXEd6ovl32K+5k5/VXTm5YyRldG
xtoAtQyMa++2bUjaiqm7nqhCdlMYeqbRNulm8Fj++npmUrlvbkUIKIwoeC25Miae7EXQMPep0Svc
yDUXdCWtRwkWNmr73UPHTVMwYfSTqG9PAoGw2y6ZcFrSY7N2ADQkqiWb0S7wEOCvmN7KwcGq1bL0
LRz4sQ3gKBAgpoaKA9j9L08PCOEelXo7mn+mH/QCJ2TMfFDKPc+b0N9jN9X7zc7MEtGTitYupzMu
gkHobSN81ORlD7gLP/Jvsa0UvGSCj/VwoDm5d7ESQ+HJdhOgAGTG15V3o4W+yfzVoJ0fm1PwPZtp
SkRhdFwRc+4dhljaX3zZcpz/MyDt9rqsmnRuFc1XhlFJWBzFSmsY6xIpEOy/yP40RDWtOhYYyiX8
GyNFfE2z4fkDIoX6+Sqg3IVLTrThmhjavVwZ/inUAyAc5cFByifzIDXCw9fHRQoqPMVM+Kww6r8h
EbwT/7L24xx6MzZ+fQgzUwESKO3en4tvdJGvXYMhpiMiwG315BPO08JSWypBUtDBoZPQA1QPq7Br
wB8dBeDTm8KdYdtGUxcyJToXhjkHWhIX0cU/8yTUEp2X0zxqQV0Ubbdj47I15IfoxzuOfMIOwx+7
annpYS9oYo9jml4AubdxrZREyR9Udw87TfzNWB10GUmygyV5ZTeYQ8O8PeZfJJQgZMwdvVE9fYgA
zi9uPoZ3+lRabuIM2/gvw0fedqy+kSCpYNtckB01x+9iV0BL2xWeBzoknPNPgZHEhdz/a9L6GkkK
ECOh1vBI3LZ3oII6FtIn0ayR0G1kHqHP7Sa1FeaGe75TY3STLNy15bJQECe6UxYLsHYAiJJa5e3X
EurrogbnG+MY7Seie7jWPfXfwrsJeMvPAFoZfQ5PNz0O89ZkrA+RLFeZE9EoFdKfENcyIbkdjf0B
IKm6GRDUGwJJ+E9luLP34qMICce45T2wnV5Tpi9e/7hW8sKVDi6jOBNFv2AoBRs0AtXvIIlBWYPT
5WqITZRgRajVFey9ufAZs/bQ7IMRDop0i6UHfa3aJVFvnoAxAniqsB2oP7tOlGD1S61dIyotUBo3
GrrGlYXFCd8sjiN1TdeQYX6w6CL1mSKsrw1zkQjxR7lPN1g/bYUYcC3suPy7t5/ol1f1VaZMyYtJ
FntHmQnW9YY96s43tc7RL43zvFbH3aXd8awE2dGkCbXHgo8ETN9DyS0IiEISoh7AcBkPpFd2AVGW
AOrm+jsOZl5rFLHLIw3rC3HLW6wRU+kEnjsF/wJwmP9I50oAV7h+4OiiVcEfyT9h8ppBM13LEOhg
hzZ52+YuolTBVeU7dBV4Auwjh8dZ9vuZhBw0qE9vwaZao35J2itNkvunBEuM6T3vgcp6BRu2NC9j
K69YNYncW0+LaFrq9ExkjlD21WZ8HwU0U5RUVqWjVkdMD1PviPyPyjmeONYj28C4W7y2YWWwis57
FYpjPKDvQVLz5QIj4JTN/LJDOpLj5kGhLPX6GWscXC40zGqQkPlivtb9cCpvLqYo9+zj+SqGBNtV
SM3qKh7IeaZEFtMXX94cBd0Bb+oQM7RU+3kEPHHFpRkJPoqewLxZY4+CMITYb1ev3E7jNvApiqJX
xAElR6JvmQdTD8V3+m7uNQBdcjiUk7z9EKctDSgY1Sh/tH8dG49uPH7yzIi0pW3ANlvkgkvkxCsV
tr//JIPxm+U77VkxmB8y6gabIJupXSkjG820aqnA9+d1upzKAo8ZH/QtkIse9tZ0Q7MWRsc+y4Q/
0h2nrLR5KYk9Iw1qkxfzpMtOkGnBMeeq7+zHjPEkbYPyGm6zd+h0kIBmOsWYGjus0AjAjH0zq08y
LhjByNbUtHciFCo8mRncmvNMVyzV3l5sL564WKtB4tgia93CXaY5m30UsCiAjSoEorJH4xOaOk7U
7IgnsFjbXoqpbz9QGurZV+YAAj4eTeufkFkUFNGuVqrWsNHEyjFz6FE5YbHDo1uPy0lSmlNb7hvW
4i624jpxSWL8I7rQFjDVSgiav2noPPZyb+ocTKTmBiu/g019XDuCs4uqZJ5w3sqiSPo9r7hYEZmE
CMMQIL6uN73WHChy3/ynkv1lRWcmGsJ7VUZDUM4EiKqr7u1mBxXM1F5ENbV/AuFa5ZCw7n/Wgc4h
zZLalc8oZHMSTIRKjyCbOGglunujdjzeqBEmnCgU+1ZjNZ+8yvJGDGlh9G1IBVQiy4HTNu5x2geF
iLbNSfRtTGyn3irU6s6USfkxWQbDH1H96nCIibuJR28XV3rOb7WPIhP4PTm7ZDF7Yx6HgnL4Byql
S2NoYS7Qqi7LUTp00kB/GiqIIIt9VwBw2m4lmi4f5/0EBBE/aWuhfHFj2CMPpQ2F7ZzqlGTnTMW1
J0jL3AV7sIlEeJnyo7g+ImPHx7xUV94zeSB11su1kluioP9EiatKraXoZSRkpeSV1exyJOQdxJYK
n60xw35AJ3ROIrNSPXQTixCk/bFIslmGTk5HHdA3O7+gL19ylIr1kbjr1ZKCxL8Bw5xYrAf+MEJs
n113cdJ3Mi7YRKLp43C4ba+eHpgmld61VxLgwisQUzxi9iCF+YtmcZDJ8O3zKH5dFSvqS2xurw8O
PSoy5JO6lS4CgGqNBsKMRXa4mfPLEoVB9NMH3Ths34IPhpDXebOUHA3oAUH7zt6j4KJCkmqGnXRD
Ya7oSteCO1sOsQZDOEmB9RJSjkZRj2t/O5WzTcZPgfOqMNvP967PEOlsyiXh2KCvd3nGmUODQfoI
h8vJ4S8vj2v1b/2TIy1jpYya71TXYmT7X+XwOAumzAH2A6MX77aBwvX1//y79huEIRT6k4kFm80U
xBkG0tu8Gyv5VzmJodPYgl06XqvWRf/j3kM9God5z1nYjTbTtRTU61x9B9Om9sbqdSTarhOPFkdM
XwC5qnqWz1xUxnt3Gwy97OpohlLNHBCHHRhkLmM65wXPgflW947pZfbBSU7pSroc5o7gaAhI14Hm
zjr8h8oAG4OxD9MIlxFXXXP5DBI8YJYh1MxghT24KOggh1okEPyydM4coSuLd+GaV9EGzQOTZwzv
yspO8kD+J1j6mu/aTsngxupluMSX8pzhOX1wTXTQ0z2oia2gQR5mHT563HY0TMOUX1oEdy5v6631
Nz+hQD8lN+mUowzVqG2q2QP71eFVwNfJY4mxajYhHEzjgZsCUcKMp5WzvJcx82tn2FxL/qBOqbIy
wdu1aMSN7Z/4+BcuWhptVt0rs9YQR4uhegBtDZ5r/UuKwhS1e4FzvrKT7UxoZKA2W1qc3xo/kyYu
0dtdYrkTyi2Ny+zjrkDvswlmKQu93rBXu7BTnIUFBiWKBFRqsEQNroKxPl7XXOs4QuTD2lqba9Eq
mfNPFh9l5NxJylpeMYvcjaCpf2TIWdT/pPacKucOJxEYbkOzpk8Kwb574uSrxJ0dzGX6sXxKVF+o
5WKeGX3sgaaQ1vqBTG3y94uOH3iUjd8fc5dljU9MjbuQz26LdhjCJRkt/OW+QJ1dp8WJSwZMydAl
vxqJnSwtvhLwj6556WQhFZxALs0gSFp32xdX8xFxjchbptycJgByfGQl7uKdGDez2nFg4nybV0r2
OoN9XExpCyI+46uKbBKkRaKVh3g1hZ0Tb7rjcdLlLZPrYVCCFy/31VKcZ5O4MjgOO7tg9ztia8We
HHeKK63Z4spuw9PdMYQcpapYkIkLdWR9lGLzP/BYcc7xeYWlNz2w36cLnd79Ieka1GYAS/QWP4Se
yenrOSW258hAB3SuHGs7vQVWeglZU1Vb6XypFxNCddQdwzPVbwGnabE9JhWXnxMEjJ9CXgrYJX35
EVWICm4kXRwQYZw6PsJfllZXbDuguWDP+ghpTLJbhXj5vWWH33hHJZADpO7kURzWT7hlt1BNm2Fq
Y7iVS0+0LqG7oHk8t79S1kC9oKYvykT26XdJgm7MfcC54xXKOuf+ecQ4I2Zz/5WwViGS5hwshHyL
u1dcnSoEFhS6GKoEV2lZkh0AMN80/nT/vzcAL7z6r5sBv1Dww3rzibhyDA3LWD1imEUTH1ug3nt+
/LhAy4IF/1QyCoL7OmkQZIuXwdCbXQzmjpj13wNTItFyGQwEfdS6htmD9E6C3q8x4yt0davNOd8t
nEN3FEFgjRUt/dn4eAizMhTA8Brzzv8q2FMvI00wPskyXZxJYWlgxs1FwRmNOJE2udlmN2zffN1x
wbEIMV+dKrIT+r0mqtS03FqK6g8AF7/PeME2rgrQ5CmDsjoHNAUuSi4XniWGc6W2fPvRSRwrUG/+
M3JYtNR/9iucYNZni7Q/XL6hAfMEtzWIIZ7L8xusvie56Ziv/HTQZEICPNmsS2MkCAG6ZnvbcMXB
RQorI7yf0MFdUxdF5rq8Lcr+SA45TVb9K9pQaNJyaY0T3uR+tEx3Xn/quAnLv9ZBG1uUM1M1lFbK
3OCd+pgwUolFz9kMJbG37WJvloz4sZn1KnPrOFRhIEXNodBQEYPXKSEQz2b94srbFDfCREMOfY3c
viHtTqdQHH2L+1JbgYNOdOQQIdhgJbU2wJ7YRhGjmfQOweOfqoKDd5WMjobiJ9K2Vbu1Zp+NuihI
e+gpg5ymPVD0uHEusXs1kUI95quCiQZlDqIoajM5FHMvrBsU4MmEUDZkqFmutWm0hAvUG5lfrcOW
9ldL1QPXpucZSOPf6vF7+FwrcSEE0o+GIDW1z4kCPXVswCOyIxgqyNQIUdnz2Cc6lKl3hpUjwQWy
jQfg62vhS8l8+dnafDjg4Fb5c+LeYjy2PyQRjW4xFHCH9P14i1aNGV9iGGTwnlBspTS6eHcL43Hp
BrD/XpXkQvsqIw0xtrjXdT16Ps7yfbWznt4lsMaHmuv426xxc0Y3eLUcijDDpQy1xla2I4V5vmaY
avClv2iPb2RaGjhIGGteS/SnkVN5R81a1bJgxfb32XGp6v/bYmd5gvHzdjhgotpZJOBR/18dXIZN
pnuFjwZCwOlm6a0PjgFXzXcxaDmWDe0+r3O37LBIO5Cv+RLHZn3C/vHnxOG7bolle374LVgF1aY9
vzUMjaqNp0YZChY+xe4W1nWF/oSsS4KsAW2jIvGrSdYV3qlH8Hwpn/YDFCHZ0G3J9aMgmrkCSZDI
4Njjk5ElIK/C4PCW3IbmfQPZO2dziZGEVTe6jh/So/G1Lsae8rIW3+De5seHYaQdV5LorgB+BPAp
w0YOyZHUTCOpV5FU1+vohNfUrNt+XIGrZm3wU2Zdb7Ie1eHbYjnj4Y/xL75qJcNe+G4kDGCNJlmT
rn/IaHRxXNg4wCm+9lMPnZb6dYMvKl9oQiSl2n1Sg/LBiWhjltHaanDpgcUUb/RP3IAYaQMR+dDS
ic0sm/rJvk5lucKTNEoOse0bh5D0CyKiP3zjzQiy+HuuMP8OveK55Y4WWxUJHanTHTDbnYoX8y9J
NXSEX1/PcLHUubEjuGRxuVGRppYGx0HLeWRTw8hBlDgHv2LW3UglAA4nc1swcYsdp2JUNkZY0Eh2
P6PM4Df+m3m4Pjf8vrbWdtqfNhlUCZ7m3PBNdVF0uVRr0b1FcO1c0TEkDtUR6Bpveb0/1KIa2LZO
ZuO2KyjDQry4EaJ5fnV1Th3XPSmh5U0bhNl7fi1rEeetM2eLBwAzN7CrEDrhHpsCDqFbEbzuUwdN
1J3UnpYlR99gBOnjhYJIgqydH9B0cPgCa87XYR4DaohpWhWUtIGq6iR2omSC/KSI9QVJzhPKxhUw
JZyFpZ609rgOI4ZzobDjFQtBzn4aBN42iagDQQyKH1hm2GFTrzyRej/5W9PbSCprHmURWn0Ny7Jb
KroPwramkOFMoe2GEx7ZF9gUMS1UC8IADbleoA18nmHjbBwzxJ12M1l6TiO/7jreKg2PzFK5GtBN
LSMckpvQ/saqtyTgSAatsREJsjfUKie/DCCYKuLQEcJpxLJjV40BgdQzjFk2oP49V2Zxzd1hktJw
yEbikFi+S6bx1MK0UBxaDF6Z+cxEXxumrhWhKa8opddlADArN5Gy59SjR7Bo88wTpffdWE69I/XS
kseWAT57LdAJBCdkAoK2vIC1HWTdiE9ecRB9s8GQIZ+VgPdT5dcY+z7wXiDXACK0bKeLPMwHyRzE
DLLa8QEbaRVbObebMRdojPcJ2/Yr1BI09GGZgs2XcA+eKL6OsNjm7uTILm0pCwfB2+jZ+5+0OA8O
2UKGHPvi0sWmu34ooJWCvrBsdNpNMxN62OOLchC5zKLMFbdfSS1iFxV3WhmXOIlNNvrpQIYkMUeq
WnvdKbxoFIiXOqvenGV2TEL7+6GdIAVSQd40pQOIHyU1WfrfkC/23Z7EwUH7As7m2rUNVmYlvzvE
NiyKwePlO/yW6iPOIXZBpZNDbDG4CjhNHuy9Zp49iQJ7BL+lXSejfhRYQ+uwFPnF/OZVaOPag1o/
tes8mmuhDkOqDW+Whw9DXHFa1fC82rgkYk1EctkhryLtvE6Qa/Z94vYH7oYFXHSfA+onzX/4Jaz+
SSh3xen5qimBimHFcSJ7sjzM7j17YRsWm+4lI01VbNCiIP/fmGCSdBZdqZtkTMcxJ4ZRllBIEtXZ
n8wBkdIUTqdBvQgWz5zhLggcjDc70uE2kMkMRuHQWwlklk9m8q1/n0uFv2hWK6CaReqGvRR5nfLe
zfMWDyemS2SItN02a1Hvm2xPpigVpmjX2XIWI22/7QN6xufC/WqyG1gCDiXZZYYCXanWBX+hmHoJ
DNHZuG9OZkqPMBGBUa+2lXiDzG30ZL7yReaFWSjSHcJt5NCtCJH911ZejxPkakHNdjn4kHZBIWA/
f8ujSv7vVbRbeeeeis9K6PNjGkFcuIdUyyUTpd5Aur3OzJAhSH8ev0YZBh4kfvbiiH6G0Ls6Lc5Z
7GiyasEmVVwBC42ZB6Nft33a0KDwcQX3x3puk8ZkYyS1DLsbgIwuudcjfpP40g1YJ12yn9wRu6bh
TlpJBf+6pkukMxv19+u32LulNSEI13Ls94Kthr8l0wov4+oJuS14z555SHV6MpMdklYZ+1elP5BV
5QE8xbysRUTGuN22Yxw7DAEprYuURpmTvdItYEz4UR7ofHmfqQAwRm49kBXCvb4m9Y7k3M7lleSw
Xp0oHIqXYR9i10NqhPCYKnJnmVugcjmyN+7XRUqtGseLpTfO5xXNU8tNiYXOvvMzV1ZDlwzWshQF
sUaY+RXC9faUodlU9nviwiQKlkaSshvHMRP758Xo8OoyjJ0/TS3NYLsOVkEPiYRgDZWXGIMsvxy4
DNdAHL5FL1d9nDWLzmylhkmFn7HAROAjCnBF4fIDL9L4iAe/3rsTpB9DH4PcN1VPBmR1Rc3Mib6a
rx9W5+afct6VkJi/KYK/wiuvaYV19V525PTK6/rXjTuknxWjkNG7U2Gorhfnihd50bSihx1JEilf
L43zKd0hl+ZtHFKynGzM/ZigRVXIXEIML7cYKSNW6qtUXTapmRW1oLOgDOwW9wqtGPkNmdgYyEIp
PBGslDE8UFpV1fzr9nzi4hX9HsoaIx3BwOl/Lwsjk2DoBl99Rc2hWlwFIlmr2q+3HmS4/c29wUXP
laYBqH+IvG547xPw4acesflfHp9Mh+mc/orJPWLhcuwEhrEBgQREzSuO1RTQLnl21qw/klm6OcDK
bl/joFVsjkJcL5+IGXcxoKatM2fIP+OgZXxq3DG2llB9nwyHk54UUoFAkTmhBqZmAnC9N1+anKpp
WEloDbLxGhy/Of9mvxGp5DMGFGKz7UtbK7jNr4pL6pqYocx+c6wyGtzv9slWIUZSzG5QDSH7W90M
z2CTY+FIJzo4fiUllyPkSklEOOV/SEO7smLtq5J/pNtLTXrNX5pSOL3faUbnUoKTXsCUYal8lKTy
FSZDOphVQNN+seGaF8D3LbsUhWcNwG2pXNiq55/TWbLjxDwuUIzH7Q1lhXPuFeh9wRIb8fTOoUWR
mPSg8/Ej5ojC8a003dDWM+XRWozaAPZjQMZQ4cViWzdVdvgplVV7M7bojk+He68gVKH/5vjkrZew
6OiM3W6vrkHxsKtx17VIQjBUzBRNPLySvJ/FASerHUeXHDMHCZOPT5g76GRdJ7vfoUh4UYKH9S7j
3AYUwyCFhrmVUeSE2irIQ1A2NNc+3+GP6LrqjmRmXZkdeI3OQqGLgQ5/54WxG/9p6C6/ujPz79wD
fNpmjUDUyo+kVCCGHHkmVQMkL6st8x5Tp83zyvVZzsvI53bxXJOX6AWwJVCf0OQ+42fJN6MWmKjW
JpXjKOCJ+yc8OJ3hb1dqpCq4ziJxb91eGhQHlpeXp2MYXr0KLf/ObVWva5WwuZPjY9l+6654MX1V
ETSQsvz3CUcSCFeLtiseXLAv+tFPfUTS/ySux/eHIvSCuz0r7zW5zbksjGJDh1LvtMKCsLOZVWBq
Ehakg5gXXp632yrH79vn9OC5Lw6+fUKhCAA714L5upZq26bEAh16MOWyxTCl3uibyohGHCovCMU6
tT79rg5ZeI/LcNaZzpioelDpdlfErnVAlWXLh49bqdByVBIlqfBXWHwmYrLQAWu5uYr/TQ2mwDmS
Wla7rsPp1XUCOzNP5PnzJnFC+tywojob2sxGuYe2xQo2tOfOIhWrOFAucD374V8riw/nM7XONWRP
80dHZvvP22lcbN45UVE+unNW6teXMgE15u5Iba/ZiRwrLQ3M+S+BuhkdFlqiUReGa1qVldGIQIw1
5TCVOUugsFo5wrNmUkt1RLffsYlxYg+ifu17ZAcsXGdv6qokXFrt5jY1S9TfMLNcsM5vbr+4etJx
rDIsZ+PIXFTyEXey6Ei5Ffeo+v1zHScIxub73qfHvQPvtRzh5U/Ei5lKfk/mppKCwtzFc/lbxtGz
YMBOwyxrCwZRBHsYkW3osLQkjS9JDOQGAG5qVhpj0wc/19BJnAye3GOyQecbNdGRPdRmtqHXWhQs
qbJLQml0TDSDA8utbsrRFnOhLixIoXp1nuEF2w3CHKfbT9rYtjwTRBHkI20qO+YteMrTir+E8kL+
FQkIpJxS8/Ep/Z4TaKGCPewjjfln4IQ0d3DPIZhfIDSnqyBisfptuaKcT7CMfCIBoiXY+MUb/tz2
Dm/NJbjbvwy8I/pamKYkWriwVbYnYe6HSKFbbWKhd02RU+MN0nbv2Imo0fILyfMO0tda85ZGJ2vf
y6/WM7AtdXQVn5iTP+5SBwjyfPCLhgzvDuZ64ZlGm7zs5dtn3BQBUxrl5B+HhG/0CXTKB2eVOv60
TAxYzP5IXiVHitOE6blBaPdjrScd7PeTALydbQ4SSLs9wttbxAsWT0NNx/oRDGJV3h9t+aMjgInC
gYRykSHX1CimMaLycIWLeZQIoan2ETBihsOggqdyQDYCtgsmhuImKDJUyrEHK0RdtjXkrViPCdOF
0J6dcp3yhuvQh90e3Ygsmt2of5dH9elvAtDuiKdoEEmQU5y+tldbX/6epoYMZKEOLQyuld7JnJjd
hfF/QwmutlA+BGKHhgiUW/yebMAB+owrr9VyzguU19RiZLIu3WuveFiAucAVtyf7ynTf0oHEu8JR
kJr9CTdtcWX4AkK68EldQOnEw1//c+ggY9i+YMuERn2P7MjJueNzR3YmFu84hu7LOHz17bRakHz3
e7/IZi6jqVkrllm5J/X4xNZ73ttgU85XYZaCbKS7vfHffYOXSFBtKEF85P4FaglYf+lJj6plsEV0
XPy3DWkxSyhzTLw6owx9qA0rzCPRx+hUwCPEbjkka7D3Pqil9WXThF+g5MP9F+zx9YAPSY+ms8Nt
tTBhQ7yxWyV1Ral5Yi6axoqHx9gCne2pALiaz55mmvONFMPw80T4YZfUpckcQSrwfCnoFIZXNkJA
cOa7cL1ZSL9jLS3eRGj0pIaW99xxVyKDUtObvkqKS26Dgq6sH9IXGOMJuyVD4gOgiJF2FG6O5YY4
MFYTZolBqJli0CZruo9ZuE5RxmzKUvu2zDk8MpZGmLC7C+YPvfumY3aeWsofRU/GwBstPrFMnnFj
LnV4ihaN/LGYFkaWvFclqE8/Kff3Vwl33zIYGWN9dZ4mDMeyPaPBI8T7Fdlqnh8yrOSL3cXpwXLg
vqAYnaOPDip2YQAHt8CJMbcJf0DRs2vjlZPhMKQ+i/e6BqGdyriSLorJlMn0zXtxxOieDUsj+oIA
KZVUADtONHNGvPwSvM1nW+m3s/w4TwHzc00Ye6tg1vB5zBLqOlrj/gQJYL4TQFvevfdIsdInE6fv
JPmsSpQBiX5IaI7xvQiYhLp+VceIVANN+ACtmj2aN+0pt1nov8I0fTOaOyv8YIrWvPDKYsQpcDBa
rWXkx4LKYChjSfOTxeFjcf3XfhJi+FfkR3If0XV053oQNMFOjiz6Hkn8MXXT0pj+9fjLv654X2QT
Nr/ynRZs7RaT1Pn4BdAmn+LBI6HsR29/gGmnXgxPyLP/62xQXVjgp25jrf77O1EO/iug9Ru0DPDJ
Yjl7zxsAEWFAbr/pT8T2wfjys+72eycdnEMsiysyqVvmPO2+8wL8MTEZjtkzmatMLfVUVYWLlhYU
K/5B3zgw0fKDOTn0bDFPEPtAQnPa8tRQJaQlGDqiz/aCRlUeZAOPMqEXWsrZbxZtg85M0YtISS9C
PTaXW+sfJt2ftufcGkwyBDYfvgJ53YLetrhXWE4gpJzOeDbgozopbI5jIx4oUKu/Y8W5894qCkC6
W/O+QuJP/5x7RcLwDUKPS4tUUlOAdBYRRc4ROO/OJEMkPEPVB/7Oyydbf9aNwA1sGDzRk0oU/l0L
sknIDAiNBEmPivY2GHDWbNZNUNH1GlpcQKFzbk3LxxT+diRHX8y4hB7/6FVyLoH08yhChwZXUCLg
f00JzEET6M9v7UwL3hot/SWn8fTV7fW77w8wpZVYBl+MMtYc6+QWZnW6TYLncLhQWFyyaaXssern
sqBsRCQm9+PvRPk4LJeNOiNTlsbNd6KUT3JrilveS/6pcCUOdVp6Ytafggmud/WjsO7kJNA56bGj
6wrecpySPray99hOJCQZZJwA/VGIJwh522WIYpRtbKUVC720L6oFMmg7dqMqS7aBsxP8/GENuPCh
anup/+R3A3QPZDnwTcBSdNO8g+wPDY9SvVmSEnJ3j9Vn3uYp9423kGvMlWoVl1ViGhqpYn2HbfcG
4Z1VV1NjiTQnzGpALB1juTEkR47/RdGDeGmyxePZ/iqEdlBnLnnPVkvfuMX23ElluJ6NACDGWms6
R+L+xwliM8eRm1sZb28z6qh5wv4lPUhEXXH4YJXQxeJqW/Msr0WdlS5jbwhzNMzBTtFCJ8bDdqKO
TX78RWcIavoWDMtPtpd/6GA2Qh3G098tKPdxuUNbMnYlUXtMSkjxmQFkPj7BI983f+/kX/tyvI/J
+t4t4Hj+Ns1/D1w5SOVY1PfPbt66cTxz7qcJEvuKbaSQJ5iUhL5b6mDEaFCJE99M7Ss+SVYiqEZH
jbvA1FpFnjgb65zfdKPJ55u9Zlq1kpmEyA7166qDx2pN8exm8WlDfeHDZNXF0jdz9oCWDfHAJ1Yv
4e+34mBiJWG/9p3WSiCVSfQoiPcw1b763YIJUgj5ZkqmnwjY6TX6OYPyigAEW6R7lBY+3n1J3jkv
fU9SUlPNy1FEehgC1C6G9UJGHMNbTGFB+w90jbX3A2DBGd6VY6KfdsuGhW9e1Fj4LzepXTG/EcTQ
S5ujUICmNnDarW/aAVTAGCqcqLSz8rPHcVahW8E1lrAzSVQdEcePiJCyNLbpGi3yCngGNe7xsaZI
ZYQuoA/8jCCcN9GBfGeDrEZlHxJALn4cterxrN3kfS0nRc0L38pakS6SConS3X6duz34Znxx8W2/
h0M6xbowfxb4MkpHoi2NEmB3xivqxaIIXfLqCXczxOraL4VpcYCLfaUWbPWCSpejm1HS1hEfrp/0
njuUi9Ck//8NfO0SOF5DSQeYqaNrq7c2tgV2R6FpIZoTGxoiXD0RH670cEf4QD2tXctf+z9j3dwT
da2BvekVsMLN77a1XydHPHwluUqH4ZKzTaDv0pT8ZH8dRx1IMxNCFSNsNHwW7+NJNjg/eSX5afkO
l6fBQ87zOBWG5WwfHIK3oBhjMJjLuEPbe8LeOY42ZJgDFyxPaViEsgie7AqG6SJGRgfZ9QFUaSvA
km2951/Ti53GkNvDhWedtA2HsSJVNUS3JUp1GZ3fvgEPj0ozccu0MBTcwVrC5sb41Xirbel2M3ro
vbcAOlWumC/SP2yHnApVfkfWs8+1xNjFU9Le51M4gHs4dbVj16YMxV0aizyPRG1LJUhQDXPkE+3A
ipgjQpFrUGcFQ/2EWqYqP0EbEI9VZ0cUpXEKYj/mEh5z8Fmi58WQcsmYuHKO/HhgyjBIso5i9DOJ
8+qwCtIC+KA+XuzF6+KISV5hvOKIO4vgX4+AqzlTKZiD7mWpShTvnwEdzrVn+K69WeUR3rkEny/7
L0GrSqf2aHR1n4ifuk5RGPp2cC6UyFF5hPKr1MqEZ0aP0OTGlw1HpaPcgFR0lMrFWHtvi/bGUIWJ
a3T3bZWVSfhI280r/YduG2gsxkFJyPWwAoh6Dal13vL2/u7nMrU77U/VNQ0kteMD9ty15HjnD9J2
YnIxcNkyCWt+hJ5gqKP9sqEddgoSh2GzUSlEpI6R8zRqXh/Ek8TT2qkmCgpwhNtO2l4y0jSusJKD
0QRRkfke2/8n1uTGfCJZSny7MEOlielbodvFOmHuXE6OaMXdXmxTbI+KmjK8QhGXeWYO+pA5s6PX
1dIa/dUsXgPRWmyZ0g03aUd97mday38sXao2EnOh7M+r+xlok5nz2keHSfYg13eIp6sx9/QcOru9
gz5bY3fqiUMSSFQBYxwIWoUk6iWXTyZuM4/Ylw2KRZMvivJUppquZ6zQGhDLlGERcOq34NEQIFx0
r6w34ZisrLjShTY+EMQaHdQkTdcrx+DEL/XKIOMrf92Kj47JU+u2JVhKHYhzS4BsKHXeaE7b+PA2
jEfyzRqVZOwEWnLO1aAEbmZk+LTtSBgdakkv4qA/t3M0dufdasvU64lg259X+QpbFE3dHreXW4iV
xlzJEJ8Rwc2dW6j7ZzaIYbaYSYm+miDV89fieakkvoYp0SKKyAOelpW9WF/jkdCrhFrNy7lhJc1C
NGouiHzxB3JTzHwQaQbaJpljP8JNmFOcYdiEWxR7MBrOmHQ0PZmTlvAEJbiST3D9KL0A7u2bdLHe
uznHpj83bBMKbDF7MxspVfeFnRCSmClWkHCRterywnYeBnBWQwgqhNVK1tTyYpsNurPibA46MRp7
oJBOJgo3yDqcFVLQlRAJXuQibfqJiGUKf/U40h4C2ZrvxE7f4YRmYA1Deg1qpYXpqHgyrExpd1Yo
FPYdjKZJcJKYaP8/PB8tyA1m98LOUnlXGommxWiuEC5HExiEvBpPByDaVSKETyWss5d8dAsAqAkg
we4yU2aQFkCBGIJ81Y3oy3Eejplp7cNXbl45Wo8YOqhqvmaDxI6/s7CxgEAsPrhQ2gYC/oLW5XHe
ZhWixKyzW2RZLHyRIMdyJp/Il3aCXs/PR1h18GoY5kkn41s6U7wL8aOYJ8yeO/K1tSD9zSvAlOtt
oAlFWx3vMi96+csIOd+QygOx7Vv83z2sUgeDnBugbcoc/v1LNnGvvFPMKfSt+oqiUkT/bppcc/55
eQB/hY4M3vS/0/Vi4X+Qvqt4ba0BYO755N2RMIZrm37D6mkXvgFj33gAyFMw+UdVdLEX54q3n4LA
Xt35f6HSA3DMuz8+9ThW5o4u3eO189kC0E0WJ1zoLQWC/xplnpbLx3Rr3y/EX/4+FB9IyGew9Pd9
90MUhfVG5u8L3SDKy7oNJ893qSPBg25h1BOzDP3arypNYyH/5o0CoZLqge+xSjhyH6Teor0GkI1F
ROPIZr9fP8Q3hUy79BHiQB84AQL43mJC+lpSR3abNNrjLDBhYjIwK7E7XhoWcN8dlLGz4tA3d7Pl
/0A+88x9pv0shgIh/OPldd4qgyNUmzY9OhMpMQMYGZWC6adVpvUra6g0ftp9f4Ybsj2qVO5or726
9V/bHzy3udeyovNAgIL2Y7y7sexEKaFhLaP7VbDixQ7zA9XyL0JmH/7j79VnlSMrLxIwupkytEmX
ntCMreZ3UfOHTE0nScDIsX+Ghl7HfH2+833iUu4Yg7pcKpsF4Ao3a5Qx6L5NmQvi9+CCuO5PaIXE
nTuU5YJxpOCslMojj1myEbFqDsY2mSCCUte1cFmS5v8Fp9KypSmQmw7jZS4z9rO0PVPfZkRlDjUN
m8iBLgwQ/rNVNaTohxFSaCqrqnIbtpHX2wAuR2jrW6ShsS46dqY7jtjqb/lGnAYfPbVI+Yytxk/8
tSCZkauyoTLNypdaSqNGFmwNc8K7/kZ+KuKtj841w1pXMfnU1LonHuNHufU8Qv60UdlQX84vxVDr
DzuJ9PrjOitFn9ujwtHZYuNQT8w4HL50QsnHBD3ceFZRXsE/kwoBOEjLuLNs7WoGJyaMVhF/AiBs
dHPrzgXhmrTiJ5BAO5TAoLoLXSZwoihsStuUTPdym57Lu1JUqsYSgLjBItFfaa4wpnxJLZhYEOBw
Q83L8BYqHnybxMNTz7fIqepPmUTF/mOmU57JtMF/ePvhRNkmfgvrN9coJooaFIwxRsKpymU2VPM/
B0ZU2TvTAC//FJLIX7igRcdZHzNw0P9O4EL3ZqD9uUBF+7w0VLUOaEAGhD2+9nZG6mCS4gLGQYkV
QuvjbjtgMrwkOqYMzFhD+LfPHxXELXR8V4VDLYxqgZkGD1i1RMq93MrbJz+RzJeHAaLnbEiI7V1f
sJGWHCCChYtDMGZTS13p7WFU4u05UA7UoisX8PH0opmjFP/p+M28DhnUo3kN9FY6RJh3nszLLMMK
NztQc5LFCe64m65YVlp+uUJn6aN4vmZ2ApUHJT4qWE8kj6a10+eLhC9XJs9wFozmLKG20GVbzZUs
4+pTeFVwUoP/IbibIuoknelYjRJAn0a0fiFsiYeoPKfdLJADHSRwM2PsZGdKd0zupIoBi8Vk1Rrm
4DP/lTuiUWcifgvJ4BtqR68HSe/8O0UTHDhlQICDNhZFHlFAwSHtGnOacZLtOOzLjJaYqMke4Y+q
5FEuzkXOqI50qVRorhnjMsvGT9uXKgInDUGcxdoMJVL3LkiCVHUDccq2htQZqXO5pqniQmyrvj7l
6YmyqmHscziUfSnFVFmKfpTBVsvJNsmTh/031RoW/v3MIFYtJ2jYLAzeqXDi6uASh8TQkqAmcIpt
H9F2imgd7x9DJWYyvCm3R9e1aGvHL2DoEZd3wgwUwEeNKs2koI8Ba/xbevOdoB2qj8OEdRMElwmw
Fa0aoGya44nIL16H4rRCf9FU+jfUEkTElCgm5u72Fn212jELvk9pbWNDPMxqs4cf2RTEzAwPICes
0hQzndikXv7nJPAENh9tQUh8bGhhKgl34Yj2uA62mxuhKGQZWXBOex7dC4Vl6w3lHGvZs3C/VvCM
zYh0JS8txLFU6M8YHPQjAHNV9nTOWRiT96lKJrRnjkppfdK9gaVtxAEciJtqCn9p+OLn96ilrHon
60+Paby+VImNmmpv1kNZlmU3Tnx6sO2Xgo8sashbkrL8yiQo1tW4uXdjrWqK4dsIuJ+qidObW7n4
3yk2N7LGpbo9fTPJwTmQFq/MK4+FH8DJQsQLCAEw6anEgS/nymbjuc9kL/QbqTuoDUFPbU7ARbVg
SKJ099Ja2z9iyx/ABMbZRfVn9gC7d//4UtKdgGAM0nFv19JEjFq8NCeuL+xYKV2ij7zBLIChMFuE
RZiOfnyVjo7Usr3rUmyKiPASX4a2WUYRJhHeBr7pXy+g4M02yTJeLqu/QHJbzf0OovVfNDpHMcEH
lebwJJSZPal9Gkcn7fOnQYOramn4K3gZ8RgnNfPdDqXHtpNE+bLvOwrxcU/ET+3ADRl06/ntZaWJ
RBGX0fAwV8f2eUgZXJw8K1PFKHRsOjzwylSZnHK8X0tq49ZbmxvuNZlCC/MB1sf114CwsQ9vY0Ps
JQ1TB0+Hcsuk4RpgEHtcmVABDsicusC1eBOAYzKI/B0z5Qzjxiaqt7TE25kf46mFET/N0/b1GYdy
AQTiEOnolJ2JNqy+lmXkvEL269SCuZ5+vv+KFxwh7Fj7D2riZJIC75DGhZDVb+I9vWxpETWQVt4N
Fyi3TB/b10FNQiXNFTe2xdV2w2q1NhNZbgIqpr1NaEb0FrxxylDDK5tXpBDdEdn6O8ggqfzM3fEK
6RHmx29jj0aFf7NQ7qYHFka8KWh/3etd8HPzHXNj+WqN5vh6Qs0DjQxLfi1B5S5QfioAtfpxADoO
L77PenNg4J/UbHA1OPqUZU7yUlEFn87MKNgApSUdCjlhAPN7WdigA5YYMEPfnUtrap9BI/LGnrs6
TmmtN9aIpvOmI6csLwfrHFH+kecugnQO5eOMSZ4cB+dH9Xc/dXMmVE0HjcFK+4hvDfOkNEq7tecN
+ED4J2sF8wLt5k6au4rhGGvnhBth176tPCC2U0NmMFFEmqRhJRUl7LlmXaJRMUmnunEjjxugD6a8
AMc3fJw8RTWlF/Bt3plWJdT31u47ko052Ie8lNx8F7gTWZ7K7/h0Kx9WWPdpokycpBBQrLja56gE
ZLzeZvXH0897MejSmvdWIErdfbytOWStSZ/k+/bAskwrVa/vKv6dBwkUak3Os6r7nZTTiuz1CUfX
5Eggk31R66VSD4Z0p/NuTT9dpPmVTBzW6OqYURI7eZ8ZUCfmFLaShOiiAsgu8mc4EWVX3F12Qoen
oDdGa9SrAIJ1gUeq2S+Wg+aW/624fTsxPIPX8a8sH+SxA2/yy5oYiapTHwKWWo+ez/Jb7y5+pInh
mhjpcA8d7zeFPfOaal+hXW7mK7sVJAuZVvDfIQ3tzVQ7tC8IbKpGroztr8fQdXHQMADDmLyq4Q6J
jraLDacLNCCozgQ0UKyYxeHbObPbpqRtrA/9wG2KziPnJmpbgFYu5eE7ZU7YDfKT45Ku5KlOl6Fv
ina3No3BG2j4KAn9wVwCBua8EpDN72TnLSVWrZJffehRqKhPG8F6enT1EJ8spU68ehMVvwShsAF6
rLoMG0oo1enK6qoML8QtG/3DCJpogTEBCuKQvaZgmBl6KWUPEUw9JaUfB7r3mlLmPUXqmG/Q9PlS
8AHE8Fv+vbSll+mUnhh7/OApiCTeEPztQ1sWTJDc+Ca6KUo+c/42NpblUoOa5940Far6Rpm9rdfX
QFEhrciQasFEdpYaqvUEqp/DRcqgE7u0k0Bhi2m2Mn1QEyZoqn6s0jdKS4NcH+++BmB7V5NwXcbr
1Q3pRNqBoETEvleVYaEpQMcHlKoRG3Otf39BkEcJeljKsDpGZjnZyFXqc5hJYjCDV+klc8wqIKD/
3Jzf//OYiNDn3klx9ouTGt8vct9kSseNNuAmy9xDE+Du8zGQUFvYOwXFysNEHlwz+C7zDWDGU6Xb
Jln5hvZip6tvoeElF4Zm8+/0XJbxUTvuv/ejgw9OHHRiW3vggymvbcpjTr3ikA/kKiUZXnSP9Eyt
oJVHQnSk41zQ5cGwIsCVtMgRu/1Ci2+yQkw5QQI10bnTDxoTm8bbWylIzaFz2Kyh1DAb/TbRLY1M
rMyq+dQZJeI8QkkH90xUu4ijuhdYHO+LInWZS3j/hlaN0UBm3T2l/ad5V/dGDH7XzPG6XXR1BCku
OTMi9jO41MwsCXjIZTFtRq8WrjCElkpMhmyGt/H5WNb1ikd6yOM/NkD4us3Au+hgu1vQ/6albzYP
zBRLLktRcqNMmEcyT/mHT8N3rR92rST7VIeEK7p78rDZggjneTPfuohTtL4eBC5BdyhRkND3bRaY
usjp2r/OJz8FA67KYEDDuGKb8I01JFBqZPMOnfP8PBSyOgKn+hJ4EB/lIVnQMbsDiVqGUWTGmUq3
J/23V36a/TAxy9IwH4jUfl79sG1RxhHNXMEF9ev3e6ScMrbfVVFGaWkghOZ3byjDIUe9HLjUyVMK
0zA1ewFBG9h2KGPDMnece9n5y33qKE+vRvYl2MYUrVQWPu3270/5aTzr+VAjk710C8a5VJ7w42Y+
cS1EGbmEZh1qJ2pGxDXm0jJhFOOyKmC83GUh2bSL5v8MwFHjMeTZi1PFov3VE8IRBmqqiGJ+zhJI
MJIRdlKkueD6jD2SGK+BfStRPuTo1ChTkrcbwC0b9vzik2nbzOFgeA5Se3i5HWtbXbLJ0RXsLKYa
PhPPkS49Mr22fhvt2AnCo/nrDMMvMjCo+aF/w96fRGYNvbEs7GkxQstJ2cos6aSpKokI8KB9wHFB
DDQcdcMXVkHNmRHSscJNgZozT8ygdvirsuZlrxMfqv9Q1x5wdw8Ka9Vuv0Pt5woAN+Bj3X2ptRB8
mXQ/zVhHrpwzA+2hWRgeg0Mpn0NQcXrSF2RflASTXmjJ0txaSvmhJLmftnrjO/ch/VDBsrVsjYrP
kMjLsAHrUN84reEw78UMZOF88nsUjgE6oHTlVbnH4P9qn8pF0TeTA7mO3TiAiu5cpLy4eZ8ppuHC
DusHRwUvbLe5p/NjlE7ajY9b/FH0IVUTkrflr2LWRTHdWKPdV6hIA+tMB14siTEqb4ZlARzVcG1w
lt99B896y2582CiLvhlz7VdUEcKQTRe3hl8RZWo9wQgaee5bJ03nqaSQaw0yMiyO5etu9ZeF6Clx
PDq8KC9E3dxWWWnABGewwxULG6sFu6PJ3V+s2W2lPDVFmGo+qDMGcVhEcvZ0MASUrbZr2qhbCHZW
dOBx+8G8RP2Om71wITPT4T3bsiZ+l5MvsKTZ3yHbeYju3kjG+qoqwSn585oNgJB2gMOX5tEOKHZZ
USfknOYbDNR1Dr7Y0Nw/Jv8PuGGDzKJs2TMULYe6YSvRG46gVILSKjPqokqBTS4HSfD2u2bms+/R
Vjxs+DoNeoN0Dimu1X08ojzSqwqmzBteYSffwvP3+nvWEmjYUce4+2hvqZ0EAvuTRWxLB2ApdrNw
YqO4yYZ0Kctn5fjOHqoUo832Q3nN28l0HQ946kcsYZF9EreIU0Lkjv/mKC9FFD6gDfEEW8g89NV7
zaS2ueMslGW0ccigyFyNVjDg72rEOISx8vKSZf2DqHor8avhuItSD+L+5sfPu0n2GfU3tYteCtkP
PUYjsMGEKzjnQ6CQQGhKOmzxLUr+4PsRxGz/WqteAMcKktAWf1MRCbsuve/yo8yRD9cVOTEGi02o
6yYFgDHWSI+sQ59eN2Vut/7BpRQ1B29pKcUDSRGv5MYNcJlvp8xLcCZVNb7UmQHFj/jspdUv7eB6
UPhaP83SVEVWuppLu4kqsoUPBdtRJE19OSiULq2EyPhxC9X7119YBEyK7qBily19k1FUyb8kKSao
Esfr3VrfrPVPAGFdT2DDJBJQJrJCdmH81xQnJWjX3EX91IYk6mEKhIGjd5s7zZwfust1J8CqoXjh
QtKi0tponugXwvF1vC2VzUzDZQn9IYwo85A3hyhtvJYGp/EExKhdZ/NBy5grHplqlElA4Wj2lXgP
9eYtYHLK7RcpmA6O0bS+cIgCEoNFOheHPNl0yjpATuFHyW76B1d1Eb6xdbRBwl3bSTTD3Eb4CXy+
n+s+uG791hLSCZGJUwTyqKYBGq5YY0Ch2bg4pa9mIsYHf7v/SNjKYXFWzmeiLEPO+RuQ1NvGVty2
Y/KFItpkEUL+9GVyLBURhFhCc4ocFTTtSuJ39JBE5zOP8Gn0/J7RigMLQhS/QLimOiCsQEqdaO5V
YrlR0dAl9dGXN4Xr5EjzRXLHnnjBRSIy6ECgvxWhmmxQSihLo5Vc6gyhEzAZpV/CaCFrCNz8Pngs
czDYH36Ogn1CqfonW+UYEu5gKJZ96X7Gg2kZuZqHEcB+lYfcnn4y6deIr9SxL8kOhzf+KRP1RhnC
C984sMERomnrGO5pOhnjekQoMvCQSsXnQbJVjaX4cOtMx2RGT5onWbVSIMkeo7eCjuNepEZBrkYr
NPIpQUrk8JaYV923A83dLiT5DcQwb09UYqBe04AHvf6ku/12J9+SHxWb1/QU+4yPNnDT3EGDu3Aq
M8A/XJ/H6hbJ7ey3RGgmI415+O4N0MEy8sHSzy4lA6eoM/eBye4PfgSTnNrMu9H0xA4BzHIjGePY
czEqaP4skKSkoT5wbJCLsjT/am4A1NmzWlEsRs9wjNXJ3i9tLqNmmkFwxSgemLIQ8bO1eUVB/G1d
ngHmWvpLPm5ZtfS4oT4a6/lBuNsu3ig6BseT01aX8VrXiDcM045OZqT7sSQ0Tz2Gn712ZArnTnGj
CATifI+Isfl8c+lT1Ottpfa7nCF7JTkxjZPmNVLofl6E0I6YRXx9fDxhDx8mM76niEc4D3sw35Gj
Txnr//kaje8A4SuGzG9uZtfDlLdpJSSICC/Zd4SmPfyUZgiIqbFxldxB+MDthIFuwFGUiHSCqZep
rBBjPhUYD1EeClsVRO6ZIa1FECPSbQjpQ9w47xUOC5M/GXd5xqBZCgQZp/sGjgNNTksavY5kXjpo
xHhlj5EAaFCt/SFssDTn2OWrnoaa3Zuo3URIQ66GIavODxJEVdNK8NNnROm0xVIef/hMAbbsk/Ba
Jw6MPrpnfQseBtCXt1aIfrjkQZibsMhVSfYKuhWgzQ6BH+/1Mb2eJa7VIRPQfYQevW06Tf/uFz5d
n8qTjC/e3vp9z+sJo95DmK+uOUr2LZoFvgMv04cplfEje+v9wqP5Xqq8MyL46ZjYTHhphdssYEIB
tF2cFJnOzsvlsmMKJL96nk2nlZMF4hDgKzoTA43RNaPOvY1oBdwIa0lU7/EJ93p3N16FhBaJAw82
yZ+CuzdytMF6FSO1yD2+7BFcWELS/QPo/68U6XNAzorjJ6mW9PJDKrjoUgjUDD/zNqpjm6a90RUp
OOwvZAtQX0RMX1cIoUnnZGLs+uNI3A3AkLQ+3d+fDHvVfgSR47G6EOH6uVpqrAfaSk+W0rrLjSWK
4xENbnOqdLRJRZ+5XjOFvX1E1JBnXAdhZOmjgSiLLTDD894JLcJspng2SLl8DPLaIMD7D6L4e7Zx
WNeu5UN2mOwMt8t6a7JzhTW1FUBOJ7HLyH31KdqD7Xr6q5+MoLJwesQHHa0Q/ZwYlQGYkNdYBBW+
R2nR9Dj1nRtPYQWyLCnpgYSzLYibqfyNY00E4GXv5Grl2HHVFQYd4nf/BiPPuTAwTNzbTg5SHsZW
82gxd803QAg4IxZvUzF2Vqk7Zq40kKLwUHyL51t8YnFzeKSKYuK0RZ3XWVRdOIsxQvDlMmLF5x/g
wGYdPxpBJsTdQvsBuaJsLK8G78IUpykKJvHSGJAW4qKPHHiR7iG8nRqYvLEra4yNaGaL3EQfUaG6
G6s5wDL1LhwRXGIH48QjzboEVxygXaaPlfnvtJ4ShTqlMAcIsbGf4j+f12XAY5n7T5BeQfqGSHLs
emlLQGANR6WQoy4QpjQAWxqMi7g4pDTdJaVq7AE9qx7D6PoVb6ZVgvWRcWZzEJaJMPpxcvGSIwr2
lsgw3Lle2ibFJScuih3mbMyvw+/pNxw2F0nBJLh/rXJrwG8LAotuSGFHUyNLtpe4vVtDTGRgc0Hz
s+fvFtaWQDbGSxgGCCFxJpxppukaEe8k+ikJAdttqarABg+aE/grgvwtpmWIVIE3cBzxTjcmj1v2
SimF/DTMQnBHiZ0pxaclnICK/k8hUf9+ciGkGdt97JzI93YuIjFt7UZyAkzcFNIt14OdDtKG/Pcm
DwgagnuLC6CN2EqW23nb7wja7CjVS7Lt6VfwSIHaZW/zpphYbTs3ZB/WO0ELVRBwAVThyoNJ7wcN
dDWq0lt1EVh42YuRhL/FnlTRK/9rggowhFcm2/QAasliJ5XjRqTw/IV0eRWVQpDDqakpkjIbJQES
kn33eOqXtiu4f0LU1ieMUP7QqJyT16xvuKsuO4zUq1OqYRBDhSsJZlXH1oK+NyQHMTrChVicgrzI
KOeO2uLXkRZNusQBKCdxbgTfcKnhFhbK5gVX14qOtKTdIjp+VpVAy0c3/ErLwVGXJ7963LRpkTof
wK5Foy0+QP9XtFuXjVUNkGN5kX3e53vtSW+fX87uJeELIoJQ0HIk6yxe0I6d6REgIJqHDNjgqeHp
mdMEKzdBwXisgxFk1idHhbswDe0v6um53WKQeMewA+Il2gbBrIAq0/yv7EBzYWG7M2XROhEWdnfm
lc9UGqJ389CVQsBQX0Y0W6KRPOl6Ix2n/toGllE2C6dcTZxSQ1Ajx1TMoOV3tgQKzaApWSzUnKy7
xYUBAJqo10TvmovzNQl28bTYhK2cBAKWVjBLp58e09fmW2KNrm+W+gP+oh9O8Q2V60H0udVDwKJv
5r2dH0KRyPH7CvqgaD5e1Z9G4SlpykPVsfWWtC1tERv1/mwKp26ohNzHoq0UPINM83OW305RIcm+
jBzPfRSsQ3rq4T5dq2xfgJpuEcx231yWTp9ay9hTedPWDd92+2/FvbHIhQp9H0eoGabLTvpTjarS
l5P9x1T93hxiY1m2uhAHaPqPkKsZCcpqcVQLk1vM6ttlzQ5nAvy1eoGPD1VgG0/6+SnjM/zESKYD
twfBPd8I16K7OwEW7+neznzPFLY1jxKhn9Re2NnqW+9FRewZ4+IGoNgQG+Z+aG6bdQwMEyWbAQoJ
1OpEfKQrhce8WwHXzR3nV3O1BgbB75cR6PeI9pNoafsdyh37Lhvy8cNjIT/7pRANyPNXGWuL6QY5
w7+3O76QaQxNwea0DYXTYszIVWCw5T35LYoKb98Jsefmc65BdRrH13po6JPwJVieKZvs3e8NyO2u
gOvA6X8EszF2QDI7XGN97kYx7PDMh9wkuWOoJVt1TwAo4jnlZiFtCyHXTd8nFS51zxAdMmp+rsEd
orJk9jVC/cB4d24tM3K1e4PQUGdyrsif+GUN5OTOt3Z37Se9/Dr7IPj3AX/WlcyiMaBdTm1xH8LA
TqOEKqvzU1f5iJ8PrX2mwHOGnDDv7RIZw80RuxOdZbzLfFh4UosrI8hNizzKVrI+XT4AZQCj9XW9
VkiUBlxDbv5WUikF5H2aqKrpLBnppAbIq/EU+hRBx1iXZ8Dd35HvdP7ki3Q54hoaW924qoec9HiO
3j5kxnMVzcSOMjeIjc35sOXNqYLL37dEriN9lA/6ZgALKNcZWWM+YbPFqOJDdl6qLMgWJj15KrPM
y9/vWQ5rnAahKEvbRIsS9ZwrzUAFIxU0gdghndTFO18gjVHoKS9vKVIr9Qh1mxWRVdWZp9ZPsVTm
+LRVFv5PNROtZ3ywPAuFJc/ugbhGufCSlTPKv6tW9Cbwo3uhTwy2mnddgplKdluNovEjV/OqyvPZ
Y7lBN5c+A3Pl4jc/XnXIhDs4+ShCiBU/OqbBuh4yNAzpbA8DVG2dEh1Qu44ylEXFWgSwCM98MhIP
BHB6U/ub3ToB9n5GcDi7K+nMOfTNy3DHq5/1vWe635goHa8kGOtpX2hVlazt5ftkb0zGYCXm2Bem
/zXqwOVA6FP8V9Dgr7fBLJgtOqhEifck7e4SY07DsTVtATNISQAxerwxK7siXkC2EXR13feLUlLJ
G4LXdTq96e+brC4NGleq5m8hIeGfYAnSHW5VqNr/v5pZugF9rgsTRV41ftdkDYOxBDNzowH5TDmp
Qcq1EWmqe3hzGc/aqXrOOKi7zwm+m82PapAVBQa585k81FOUGHFpJCBckZMf6FW96SmWB39+hwJM
m8gB9/Xc/ontuSnd2IuU7pUtLrY4Gh5HlxMnU+CLKkqOtw19jKADZrXVV8um2WklDnKO1K3SuAle
Hrnp4d0YPeL1oGwdmNsqMFRf0J3uE893d+jEIFZj4xpsvQGXHvRZQDiITrbaYPD3lbOKuviStjmP
2C8hcILyncdZjMM62MlTakyIW7J3jDPjidY2YqygpiPlUowEnxJeky2ZYq7Wtc2UncAzcPHAFm/Z
Cx4WZdrWbsH4Rop+o+NX9pC+3FFIcTLruGEaVY194BgK8Gm0ZR/BTR5jx2l13BybfUIIlzUpl0ia
Wh/HN3W6Idjfl13aK9MGTXmQl8ZhSujOl3th8c3ux428H/ZCMednmt8yd/xA/8p8Fi16SR41QvGZ
IiRpEelThXOSe5TyGdkOVVhOeWlxU7VIIB3vHF/LequTPktmn2bzhGthz+STwRMfNnC1+S/lqGkF
M6f4NWzoEtm4oIzVvlMurV270V1vlJJUjo+6F1xA3ZHggV2Sm+Z0wyEU57s6Cr5ZurBm3Kzdzaym
G+kn6e7M9MsdHUuy6yri9/xJLL7/uL+SLDkeLyLaDWgHAvvF460osG6Zjl75xOgP7nektOU1MYuk
koJ95dGHdqrBTrzz3aI4CmU0jyzLRn6eGeIyUu0UcCOcP3NqASiMRH8+C4wCOUjWwnq/4ScVeo5Q
X1AqC+8B9cJTnJ55ajLwSfr+ay6hDPPC3eEG+pd5OhW0tQwm914IDH+mh76icoRL/MM5VvuBh30A
WMPoHvH2KIgh5AOggOkmrOTqN5W+VvGvVFBl2v2eMxFBh4dYvZYXON9XgHf0fHYrijpaO6J1r7cy
7xbTcna4sbsikp5k+iOPBxGBtLFxLy/IknUoyTJHJ9F0Wp2Xqc4neeLkw6K12iQd45hskfO8fDMR
RXDUTsmTePU9lmauUbjnG6YyJwVrAenK5wxwcbJDGMg/uBdVasqnN35DCqjvsjeNHor6DIKqvRxE
Rp4rwGd/7gysh/Ydrc6VrrAFRgSkX7ubKiGJMO7SXyVpy7alcaMdTiNfZwcBx2GHlmUtiY7zmnZN
nE7tiM0/RZFyqgop4lnuYgdXG7varkZM2qZ8vmIC1hUBhL6boqK+RDo77TsuHZIDANA3YrNt9n4F
BEnr6eDTrWB9Iy8I2/7y0dJggnQQtGv8ftKV1LKH7uE1xPsIcB0fj181PSBN7rkTRfv6JoECv0VT
OZ3mHO88EK31Hg3QKLcTmiqlMlNBolTE8solhVQYNCO0DRE3HSLN5jS5I7QSP0+80OmPF1MUph7d
cxa/UTDH+C6eB5VJk6ksZ2neoF/NLArHnmiMyIDNKG6LkUM2nfInkfnDrsJxKbvf0+sX1AZgsPGr
jOjY8PymTsWVQRSLMTxYEg+5Kfr8Rgrqu3Fnl2AD3IL/aLPY4QXaDnJ7OpwzmLGz35J0XN4Xv0Id
/iduVDvc7xDxqE4NXvxoWJpAzEQKpKKM3EDCMuH4qCQlGFU9koXUYLmXONSEBAwyZKXmyxglqv1b
CLSMERuL/FlMdSc24FnJwwFvDquuUV3H4OB4zR1uXa7jqUhr/mYnfkFZLh87Y7iRYPX4nTeNO3Zs
3xoh/qcsBsFikffnt/QhPSbWEitHXl/nqukgmRTIXqGQTmnuUyhJ8pLbsuB+ojz1Nxd3ccS3d3jq
ov2GQSgq3WqBmuKl/xufVO+CSVQldFa2fMgXQzcNnIRSdRn3oSngTNOeKShZOdd0kMWtvVVU7B5Q
vSX3NxLtSmQhdZyLxXNaIjIVS6yQpSl2cAe2/oeU1oCUn56bcoKmYoQu0BlrmrarjItZV+U3AqZT
Ggf5QnDBPxwGYGNYsU0qUt5L7wDACxBeiApYRwn0RKVjeJ5+KAryhDB48vWip765ecIarcJOmZre
LMfN7eD1YmxmcOuoyTeBNF30AiiCfflCcJ/Qk5oIr2pJL5KL+AjP5zPI2xESZ+BrCp+sgd8tu3dj
0Ba7JdnorOYN8zKQuzmZty3Rm3MaVhzkEtiwy2hha7WWEz7eXSESaqO644UkEj7Z+9Eqbmr2eppI
y6IqmcEvNdaQ2OmWdtKR6O7aAGy2IZoaaQeVXfrCTpo7MdrgcZnIxtaG/+UCejBIAAhzOsiItcXT
RVb8JA6eqwcP0H5TGZVPwaZZ9CM8MDwyxUE5ubQwmwBO9zmwR5MFj8NB818c8rY3gEkgjxCzflzP
p5T5zojpfpOfG/m0WULYeIzq2AOj0o/++YIhwQvQKsCfZ88jo+28AB9m8Afce/ioKLnHCLOLHiAg
1BsFpJG4ehq5gk7/6mqAngNUBsNCrF6M/see7dG+2K0+87E43mziFM9ddzbYOczNrTdnxGcWlHO1
xK+NVl1kRuvhsutKvuBcGzFeuChLu/eDZrY4ZP5Oa1zGuRZDNK9JYGhJv+Qm1WKCMBFGcvi/LlQs
bazEEW28f4bwbCxQ94j/XzZQVIzRi9X/UOxhuTO9Dw9wYNB0miRpbfJLUe0sLIPW/TAunx1iFUpN
lTzt8ZUy+9R2sZNTc+o2LtJ5qoDEhJjN3Hb2CGsdqMuXaT+M7SBdkZSvBCKrWkZbUF5SKJMVOXwQ
DQ641XM/uB0lgF0e0kiFwvo3oni+FMsEdBHpPuXPlNBPsHASOOuxsMfn+W77e32NWeuLNovBj8JT
I6thCmg3uX0/y+eXPF/5oTuZ6uVRehawyjM4RUK07njzR92guWZ85vywXgQcraDOlHZN8u0Ylk5i
4SESrJEFiX4FoAhq8FErXJ9hj/YZI5ZKeV7jRQ6oLmnF1R9wu67S3kgsVW5lSBg0KzjJ+W72mryX
aA5azmvcTb+l0sLkuE5LqMBrWKFJQ8rkUVncQVWEqwSN8lbkN1LBHu92LWkynrtWDlO3H65pk3Bd
VpzpI7CwuJAJ2e6uMWqDJdHNgGVfvSU6+JF6ZWxT9VDHZnFOUDnhZ5Cais0gZdrkPBFl4JqZK84i
g6BZ3YwWQgKXhbugqZ0y8KJAYPARuHIuWaUKWMP+u5IwUQDmDGLO7GO0sfBmwT/fL1Npm6M4KQ1/
y0KgbWSoMfQEp16wyTst+nlmvJyQIwxKpmqA2f54m6ICFfbfe4yOCINqQbrFMiBgcjF55fc4NZEM
wjYqWqMpXfpZFfkyeUUzMaEX+yR3d+aEAgOexWlF2NiQK34oxL2e41QAdc1y0KkgEVLb/Lg9gH25
FmnqlYj5XgFkpbIDwptPzXtUJM6kphxDUNOQYgsVCEl0i6lWZAErNaBr3fMokrmsoIM8n/wbdSJH
xSnHDHd0EqWpJOCLP610DQLgP6GnrccaBcKtSUl89SlzpYxT8otWEnn3RIJlExxEXXC/mJeoOsUj
v4lGcC5DJq/wDPc6Ou0vGZpXClzlc+/u2MX4UeFCqNKpTkTXGhgRST9zX2Bo8UfdR5TkP7WZiBsw
X77VPRV/dWsLvFuRZZJO+tGbIrcMovk9obqzdQHM1gAYUBEw6T/BAkdB0Jk+yU8zibfrbQG1RjW7
787LuXfY3yuSJ1Up+6SeMtfwsRNLr18Lhf3LtFYf1X8l5GlaotQYXdLmsXf0l1d5OctpTYZijUT4
RGMTp6U7GgkkITCVrxewgjZXjB69lT8Kf5QP6Ro/1LitOxZjqfyiiypYoFEklmIFDSX15/E8e7EZ
ZRIl6hCUxEpgWU5saH4vGN1nDFc6CDtn3eBUWEum4tnaok07Rasgn96IHS26UF+sL6TMIJE1DV4X
bcosQKph1jvHrxMTTg3qKu38E6pWuZocaQCbe8JarCBptAuXXK62IcOv58JYcsxa7Q1S5Vt08hF9
XCz0181jExGAGhvP0OatyOaLl92vnjJ32EMSiGF0qn1mfI0hUWYKk6JOh/1eE7B4Uw1kXKc6YZ9x
B622Y698Z5NZs2v2QFU7/f3hIW4ooKdFEjggWip4o/qwwLzeblARgZxAf1RfIHCNE+kf406tEXsI
kEwx+eUAPPU8By3z8gcuGse9cDD6qoI5c78K07eU/xhxaLQ9qTuFlPq4kW6zdV7gRtCis5InaFx9
Jxq9PiMrgC1HQLOsitNaEx1iHB7dBc6T9Ubd1Trg2TqCueLadnKgvETuxesjkGcpO7oxPWcfOj2Z
Lcv4XDZJiPlO2U182txQVIw8UTIq6i02bkrrNYa+dJ7xFmGA+OSNWZhmbYu6rad4/k2oAz8YTZ72
tsKoe9Hkk9KFNPyg1dpNK+VEQDsNfOr68CoqrPtUpyA7MN3GHF6bfl+6TpQ7M4saM430KAe9qGDN
Q9VUrzKbGtvYvTkmwUd9q1Kl1UqXbxAjBGJ+qQdZEwA5SC2P1fCOayPqc+n/4m33za0CQKAc0uUp
6Ds7jzOsknmQWOvxaK237C7JCJMIy0YQ9oDBjTR6EceMKfzqvgEQ0z7BJGJJGeq5RHtoT/qh8SGY
mwKnAfmse5N2FIdu6XFZPJqXGMuqXLgOuwkmWoITfumy9Ptx93EAad5UN6I29n4PX2m8oyttc2Ik
uUDzo7icQ67AcXP5LWb2sFd15LUUjy8hUoEez/LxFpDrjHiY8LOkMYgyINPImhHs4G27YmS57irT
TdAeWOnZPEnogUr+xjxk4BIij4kKW1SOkpXx/Y5fv1QA/JTe2x8+wSBTbDBd//ljTKiqqXEMVNNa
1pAtVSVtqMWDblZ2T20RCogTk6kPNg2N2s07r2DEAFGih4K9N3Bso0iim9ZVIqijq8O+FSG4GXCY
YeUVeC5HXM0reePQXz3zOi/9Iwu1vPkoevvlfDNaRAJKIt9i36bc+i9vCCwjzMUnu4byKP/bvLS8
ky/+jAdE5ByUTsy8pxKaZ7oFhhFfHKpEzQQjOG5cdzdtjxCE0+6puzZ41pBR2Ah1Vbwv7vrPfMWQ
vwQIx8/UnFnLI69cdI5Gwry/UJuyFmEi0RV/LKre6MioBqz2nPj56Y8Y0oTAcKiMrCy96GW2heGZ
6O25PPDfq0HiAwr0aJuJnz3agjwci6tnqggh8lmXDAPyHnlM266ho47ANBjYGYbi5etjv6b+5Ldl
K2vu02yiE/N+ZeV6buKNoPBT+xbuAStm9FwyAexdazhOHXf7dVRmflPtPPUbeYY5EPJ4+IY+/xKB
i6oFlrePm+nrYqSiIm8Gh89zaxb6L7u7hye7NWP9/lZsgG+ud66PTDcJ1oiSSHkbU3psqXO3UjcA
UZiVfN5MbtG8JoidqWVZF+OAgTOKdl50CIM451E+hmTiu92lNJSbu+/VYKTEoA4gJOKPtM97FRoC
li0tyo18fq93bkALRr6U5u8YlHSw8SE1V740X4MWL4jJbDk6fzqsRUYcw+WhsFvI5gHm8vpw+uJB
ioJmJevNfizT8BIVpMrkOqg9iBZ6UP+t3iJTZixPixScZ/qQDT0wDMpeRcfs+2XlDgoAnY59dk/E
rFaGsAi3GebeplbuHru2GbgsPc9fpidnMSsxuxaQ5OnhLYDPw/IptD5GxHKeFXWwbMra85ww9lXj
ibglK9rMYb7c6fLvhvBFsIcAFjMYl/ywRPRw56pptlUNRqXGvd+5fXCt1W7Dij8Wi1iE28qLUmp6
CXGJGd5GO7ccDZ90B9DQiL5dKn0Q4lws9gL9pIx8VttA4lbfAsZ/8ZtECRLG/tEjgO31FgMk7otz
B9Cnwh65GYSvCVHl7j4kBtLWcIFZy+iJuoWWWOFKd2AM+O53H94R797LLfKZ0kYQfyMp5s44ojw1
FHORT+fHrYnWg3zZSeksaXlxb6AQQF1n2iRhakp2btSAHZInylImiYi+eaIPdh903i5TrT54XoL8
gHzG9+h4+wXeTNbWMrmGiutvgKLXnmwQizTCY1hu1UBFbS5Hzw3dvdNOiUupXwMzIWwQOKYaDK1X
RGh6IwRkMf/s7pBJell1JdgAumI5n8HumfXZi5FY1S6ClUFPhs/LUQUX12bpVt6/smrjciFIq4MJ
sr072xMWZtOfLpUkejU4defGzcxrxi8b1ts3Fs1oTtD6zr/WFHfiSxNBHm1X4myHjT+1la/miEmk
SgV59pPGiIQQZaqxoMT8tMucGq2TTVNUtayZ8gDH5EBfzbS9UUNKhNzRA7wGaU6YR+quRR/MIiDi
CFOxdDrUWaMpj/txWsTJoA4c09Gn+Fzfe8MM0XW80nxKgsbWG8Cl/Hg2A53qC80vKbdlAX7qa+lc
gWnxHecvXZ8nwQAWaq3VoK/xeYAR5qCcq1RtbWT8eH4taNKV8ugb7GHsWPAqqGrKYR6uGEcvEfCt
zZI77bc29NxkvFR0aO7CMpizWJ+Lbqi/pVnC2zeRf9fhVWWJ3+nDPagtTM6Xbk70jsW2HfWN6Y9l
gZfxv0JtugiH6lkPUitTGb1TD63CP1NVxT0nDjCo3L5SrVCizk2jBK/j2Txbow4hq1hhHK9zUG+p
pqlsXLXUDG+7917aeCHAWHu+EvMP2P1x7a1O2/nGKEHMfB8E+wCTC6jGDMLYKih9EKorM/a/w5aA
xdZfjYX8Lkbawu+8wwKWZ0ERAPws1Vn2CNt3DVdxgG8k64V1vRwPar+nsNbOSeBM/Z5B+FPeubZe
l0rHDx7CPIbYIL/n5y5hrAlQhlfHW1Cl9HLjfYUgpqSIcjBlGv91b+lAGtF/f/zFDH8na9oqcUsp
uSmkhXnAFiIf9dpiJuogMTviotuTua/xVvUsL/Zfl9rkTpo/NL6WUZi2mx41DjEQ6pVL+MmQhmJR
G8GKaSvKEz2aJhOYe81KhKfGzsUcBqQMTbv5wCBgmM5AFDFBWhiPFG73iO1aMyszMnCp0zGoOPtG
Hh3F3D+0HyEMkRvVnqhWmv1NfjS9LGMd9U37O+/fatRfLax8cUyzJpjm/i4HAqXjisAZL5vYXW5t
KsaEa4CjQWV9R+lBx62qZ3QD+ov4XlnF8jAE3IJ5EAVJnr/RuQj6xgJzt9wpRkAEfDYHoBgmuYqB
oiJd7I1dgTb82GPRASYMewygFdEup1JEuyqP5KW1vddVjQK1JGCCxOEi/aZv9GDHusALBB/2Z1DR
CKGR+TTFXIHLOCOwGVFf4qaiW0Z24vCjGJ0M9fw27LI1Da/G+TFMkhJ0tBTPwlts5ujTWkj2VWb7
fHRiUuRumyqHzifx0eSfWqpMlPiJcJknwvqVZ17FlZKRg8t7KKSpwF4/6qyE5szSRUrExmgi+/3F
lag7KbRI8vvcCfs60FgD/q3L2UZ0DUUx6ZZjW5WFzfrDV5YnC09BcyLHCdxihYcFheQAQVY27hgW
pZxqPC6QOQZf/X3zaHzRm8Kmi162b8HxRKSs2TrDJFbu8dXjZHCCeiMbafzN5QVXGEPQ5NHwuha3
89BoF3WwWHwBQMDPMhVIK5sY4TME5VltEqygYUlgd3KZcL39QwF4QoP3jdJIHm0V5UBiNSgBn6y2
wpOLwdiZHP3ymEg7KwazA/pgnltSeh4G5goGqjNilBhE2axJIorfR7f041opDk7Qn1IzbSMQz9Hx
fnOaVBGBDdWM+wlc/FCFBXOz+KwdBjijKaNVrupzZiNWpqhacxR51ydSd4DLkuGduusyiy8MBY5s
AL4PS9MFmtY26Nw7q7b7fK+alZFVfjSuWqS2aE1hmcVN/H67iRTpFiz+1mv9JpH+SA9Zi1q1OVEl
Fu7QeL8JQv4wWcSRWvpR6zPguxTnaIDzQe37Ji7yQLiTumNGg6Hp7ZLWuhhY7t3C0leO13PWy2+Q
kgMpdZf9oQy7H3TWUpKYlMTwDSuuBRYeOotwYWlp43OFwNIVs+uZ0upVRYW/pJLjhRx/2FHSu5u4
bm/BtICD2Dzqt19rclMQs+T0XwblCH0eFQAV4mLsRV8v/7byP2jSeuLKPkzoc7PVokRCLpvI6psa
tj9zGssI5UYZsTSoRCPbvyx2pu4x2EdSRwMri/2MGfY/0HrsSN8bfs4O3DVAaduF+uQ2qas5LYth
k92M3KKFRuRIFivkC+viIt5R/TPhiAyyu34ETRJPOWZ1n8usLu9YZ+LrloA6aA1XfphHsT2xRbl+
/uW5X0WGt6f0JXYTsTA7hhapFxXWr1VHMeWUIPhsJhEDNhJYd/ZacEpL6syGuFpJMaSJNZKImbga
ufvmctLNKsxo4qYOJsySCkBmnvLwiVX6mJaj1pAPmapS1hbc/lCF8JEmrvPJx8ata4nsHiyhkCyc
NqisKx3gcicB/i44p9REKqxBA9m6Uo68N/Q4tTJuNr8dyzmWCe+VgiITCIU0zhHBlojGbfUDH/ET
hVKJpm1jZ2wRWu21U6NhBFYXzezUfypz8zAhUqRjnFU67TB2fps1OJohM5sOq7QjVl/XyCCxUtbn
/DuBXZQGIDv4rnwwBzT8ixYtoe64FZlORu+BHa/81GqEPWEc+7BC8JSuRaSa9gAvaCIxaCzKZ4Km
L8UyjryewSYcC3AcqDlaqIHi2csV4LK2cUHxXc/Rze2/T7pNuJRS8YYAiXGCsEHKsAAWwEuU5Cjg
FyvYFIEGmS7szQ5ewj5l8REhwvDKiPitnnIUmMQ9BulqoNwsvXlWIVdynFQByesW5zZP8tceX2gU
jZXkL+NIttzL/bRFtmgiwG1PJU2qwSkubLDAKhnSvH61004xCiLN6hIH0zHu9cGrE2ahW/raIeqX
6d5EOP0a7t4L8IcYXjBZWeECgOz1pl++Q/vS+YZ2kSFalEJ8D0cRwbsguY1NFlo+5KKfFB+5K1wq
wj/vSvGfYiLjKGeGwHkOqRrpYAtW+SZwTcc73CwzmpvQjF4BcWlafayOUagkaxCe5CISVVXml6eO
85W/C8wAr6Sa9sLlSGS/mbMcaLJww0qfp33IyLRFhAeCIsh3je/mPgyI3gfEGBIoNG6R5FpB2Rhc
W41cTJAd8wBEa1YV+rjkqo5zDbdW9cNdTHgwODzdiKeRXb//TNcNrUco693YmSaJVuS4rGnX9YuU
+fGKPRR9vO8BB9h1zuKnPgKjDVmfM0AtzAcZ55eXYknjzFBVX4+bpBZL04KKaqndR9SnN9n429CG
DyrKOVDEeg6REMYyf0WpHpHYYDxvAysMB3n7+/4QaucexTz8v8MsZ6SoQMLxbzJNfdijv10rOG4D
hfX4iWBBqE0kvk29hGlcDMuSvAlHwrWiEevVmqlk6MFah49NKVAQ8gKv90NZW+OUIoh1bf8xHyxX
FpZBclTiNEiB7u8CSy+YEsPjWQ8WyeceqUJOVSJ67SvUOEiRkv93H4Nm+U2gqIrmmlaq8G2pjGWM
fPjZHnCV33e1zGnKNnElmd3MY8BX3F+iPJ+VIknb9eRRYRDsHQGbzDjijotdOPezM3Gxi1JtVUhf
SZ0GfNfFcW47z2FVrbF/aTzJtAm+kL9bfz5iVdoLMD+7ifZJkT0X/eTxgbaSz7H7Uqr5E20Fnc0f
gh83M+SvW/JSbfhAF5nX9n1xa31Y4xut6XU/mrixXSkobCffo8r5ClJLo5f6bETnxAYh4vCd7Mlx
s6fQOEad6ueTyACZ36bzscBQJ12gYBOaJSukKGNhfoe7zP5ZLOfIiOA0tdxDJERF1UEA40ao9w4Y
ExMkpQvi8njbJDGuzFKznUibNSW1tWLlqJXUWInpUPNc7uOYH2CD2y2DfI55bRKn716jC00oUHpS
Oz+0q84v86gzjpvlDNkzf4p8CgEreSXmqlBPV7Cb4OcRp5AimVKjQ8t/92OMJ8r1M6Z7oa4pHriX
O5afDDYzCLu2zikShuV+yulyJy8cTvfKFd2uNeiFGDmSsDWewbtbTxqOSGHQU/0O2nNvzU+vaPWJ
inulPJi3eP20GIhDMmknmZWZZ26nbQUz+oixZVuskbXURx/O2XomMQSqNkC4GxtAONTrE4uOWJrf
Ji98ueTSgng1q8O+14FP7GtMb6PmMfzXQiyIIspC5g0RFOeiG1jpm+9tJlg3k8Fqdnr+iuVWs3gO
ymY54wibDmTn18H4sDtSqNXDs+nuvoHDMzebWLOwhWPDKa92q4X9NAlVosHPxokiLsgaJec3mRG9
YYXVcX2wY2zDXwcHgdK1ScTm4biAKlV/z+J5hvzegM4871rncKnROLfUrJ9yLYchsYgPvaU+zJB0
bnqOsHNJQN+shQgHLf8ei9CIPrezT31qKQCKC+pMxiOeFtDSnjmvd6ysW8qtTPbtVuw3TSqJ7tvF
ejmvXeAfecyha7d9sIad8LcwuD3lqT4/GLC1dHnlHDb1bMvAphD/Z83TChFWMCvVhcB3wNAKyn7q
ByV20fdIP6p8Tbcjid8O3ORKHEBFBVmDPfyKhfukEQHPxKKikCdyYVaw/T8rAfjA7FnWiL0YWcX6
UbIvU9Dkncoxi2rbRmZ/Qurzzw63Qxps249LnHHuJ480cudH3asbrH1Y9Fki6DzejMhr7x+FzDWN
zalZjSi0HLHsWqZlIaNhgdBh7beroPueStRk0XA3w6lvw7l5cDYbb4XqwGhiuWRx3LWhuq7cjs5A
Hw44l2kjMSxgg+TqTBKO1FIBFyPlRAK1slBxOPPoYa6nTKCh7FqS/b5bwyAWln2VWBBV0uLy97jL
8/RosQp6Dfc2EOXwxySVyfjCoi4XPzVkWt8EGF5pf8ySQ/S9WFwp3ask3A8il3tHj+3OCdFmPiBL
eOd3c2s5/v2Xdl4fc8ddet++RUTBcZ/IPw6BXd1Sl7GGrMzum6s8j7cwiWeGOJ56Eb52awqybxjt
6Juz342n/jtXJNhO126jXwn0/Mc21rztlWGrguLqwexF/bq4YFze1ZsWm3e+TKEYKa+5ZnI0zVCv
0xKzG8tpOF9u/67wIIWaROdPghYucHCVwQkrtxGKzWHmQXRoREsg98Bt70+ybaYiKWsICfDlrxcp
F/+82PGFmQQ7kbdqanICLwEiAH6N2AixWL1dqEUb70YMoKp/W1vn8cvNytGl03+eHDBEbb6KYef6
61sC0hu9yqQFXMcyfCleQ7mGxT+Gsl8hNXfmyug9g1Aokp8y+5AOqFGjD+gegPqoNcXqD+U1JVm1
PNCUwi/UXi5E/pXR/2OVaoqiMqzNjlGUDGR3LmEig4ArtkIHBbwV9G9GJGNbbDE/EAGRjuQz3h4k
APOjDymT8V3tZYoJChS/xEQLtamkO8+fSws6I7TIN8qhPwmkbACYtmhSl3r+cYKz05gu2H+pBpHq
MNlvE/l7772XKh9EcrooVKxIBGcKY44yZesUU8Jw8aLUHuKuniRUW/uCAhr2bfER8ZKprXGf/Hm+
ov2qCvw8xD5whpmIImdX+rzRH6pJ2d1Myr3kCNQIicL5/tz/Ody1qERZBqxsAx6cfnUWjx7ufH16
lauado/aYPZP5SZjd/9khnxbxyHiJvqfivFGYSUMXfETm5P5s9foKXGKakQVZ4Pqhq+mQlQBYped
q+GEBx3UbSE4eNcZv6uHfv2W84AYGVQ5rhOWvcIxHWOcxB2ulOUwKGjOOhhtFbCQKCAWTtnOUQ8Q
nybpjHyX7Ww8d+50Znw/jAw2YnnBOENJ3Mg9z1usO/3hhZelxkq01jxXzLdnB9Yu0R2pXQgBpU7d
UZ+wYXPjiVKTWxR5dfyj3dnb9AhgUEDbaWoKyOxwdhYo6HuhPhqjOCn5w7kGIufDWy4EmxfaQw1V
wIoEymSF9Lcf2oSus61LjbkDFvAv3hzllW26ztY1qv9kZXt8dQzlAByY/9SAybhN2WZtNEv3vuUB
oHr5/UMMp95234w2tcjn/AceV57b7NF2GocuY+pDrUK0zMbDgwl+zSStPcJC/2FKA+Ulf2IWRsc0
XcBEWVgXHTvNAJyB6yy/deBsHv9hX82HMaFVSTA1cwgUut7GszVBLJSD1xFs++krH3ozz0WLnwbi
r1LPzu4Nw9JSGoNvp5c9UNiUBBknEJyWjE/ekNlQu/Rr7IqNaKXcsrMqZmSfNk9QUqorTT90K5gU
aFU+tU32xwPSN/Lqb+0QOJJAMa1yFoCZ+/Sh5w9bjEdujO5i+c80ETAkT/EJhfwbXnYRjSQuGx54
Sr2PagWKUFcceLggZgbaors3rnBn+iiR7DR3/c/vSWKu9CF7A5qqF457GreiuOS1MvpDuXKBDscH
Kyf0K/n/7SrL8t4qTRSMEn1/ieUtZ8L1hY/ClYJ1JlYirMTQSEcl1AF1JGM3tO7PMYeCDEN8iVkk
iJAkoSGRmX/cDC/ND+sABePc+o4Cg/xzgAbqIOVYC9rC2vZJHHxDYnF1YLIMz26c4wTfnooX+Xox
RqW+nI7lvRD350JHFvSm1WacwZeGUpb5HjzJftn/FPRbVf/ysgSpGhT/CbMHQk9VxIfstDB9Jhf9
3NKca9u0sQmP1SC1cQGm1Ghruivm7W+aSwX9N9v6c8EKDNNE/YifqMSCmqUxDWd4cO/vZVrjwESf
OzR2oNuIzh1oIkUw3Suf3rUAGNbcDGoAPih+x2CgmlQOUfLjEoqCWdF/YBWz+6+CUAPoWGEdbSqj
8TAcypCRU2pOaAYnQlbUFHnytuFGEvwDhTOS+dtJYe2B3uV8kU9Wf7ljOnlalLsVHWf5s9KqlBJS
19tieK/mWbZu4jMdsbAnWb8ZPsRkZJRL4GZrtKVqvj9SBzxVexvnqut60Go3HcdS7KSQ98mhvbqS
mMB0us37BLpJqsgAtS8sc459wz3qK6UzrvQVO/XR6V8W+dGN/ka7mlODuzujdPA/iV8SgVnCjzhE
YNiJygFav1wN5qRTkRzh/D7TdYXgIhYxufA5itn+tJt1/xbi+76tnc5YcFuZi9MHM8MymO1l+O7N
o4E5Z2bT6d2sSquvP7CW1194fqFuwufxgvfPOWPYjelbhZgG35RQ7d1HANIbQTAC80mp6S9Q4xCw
isK8/XZvcdchvEqTVkMz1BWhIB3Tr+Edp71Yga8Egzn/n5EfIoe1HQZE586LmsoK9DxslIbT/G4m
hqMowxtoEEgYVtAS6iJuRkFbttUrjn8FrMo9DP8IUXeFjNQt44jmeL4TRoW1vlBOZ215c89YHuLX
OxzKYWiAYaj8e8O6oNHoxav0L6Cm1c5l5PHJOcEJkeHiOTeHgI8drUD9ElUodHAtp679hapPKW/o
1tzIagM1zwwa3z+nRuJ/gCDNfIdMdi5guhBKVDEleGWNNVxG1jhIfoYVR/mYI1Ipr5NWSpEIFp1d
mvXmfwmf7kBySAyMkiFFLW75Q8UyBlUnVzNmInDFVg/1UNJde00qzKiF4vivco7Q5S99g5hE1DHu
FklCh2Rr2Y+jXSOKnzDIMGKz9SloCuSY0aAQ9KWFGSkUUGK6aUt3IixBrDn+vayIrNhIql09QLPR
8hNO/eecdKN9j7AS28CIJ8j3t6D25dY8cvyikMmugcg7VxORX6QAfgJyEasO+PNCQYfHkItdx51v
xi6a1hEdkUx2u8L/KqWNKNgIBepHp6vMhkyUZhl8DoGddpEWATKId1AO7F/b22Qwn6MeN0xdmr5W
8qMkJL8K6z9+TtK22aybKeI36QxtPmxiBDdcKOjwOCKobdjJA2bIrncAtU41sdHxSCCIsQ/9Jswg
y7TrJzQQsFUPRwJjPjIR5EkOxq1gu33ANpH4XwgBFQtytWqcakfkGsjgVnzeDKBXsP5H3bOOU0Ao
sS8i8sieZmwwc5y+LGmCAdg4e/zYxz7fQY3isXMFjtHMVGbgphJ0ICmWlXTRQBdz+pWxEPriOYgN
SFeZNDC+GpXm9r4UTmq8U6z70hsD7l34p3yO9NWG1xO6P0zop44kgqXL5s4E/cKXPo7xro1eN6Vb
5PH4VjCjYJ6ACmmww6rM5KIjYZlog/BLKalGPRHEU5fit6FHN9YrN1xE1FizrYoahH1teolyQx7P
InP8mg+FneRkCclyN+LN2x8E8Llyam9etQqrCfg60lN6Ufwa68Zst/xO9SUHLPC2Mh5FwPkbnFrN
gMWqODrZvtHG+AJPgjfCqQNfvKxF8pOPzgfwmZ4wlT/f8MtITaIqXKy29fWi86v9cZzPRWAMR9V6
RbiC2WCe0Bj3H9jiJZ4EOglKS69kt8Jg5EV1T2Tc79OAchlF78u8l4ysI/Xo3Z4b6tFr5WmzOPxJ
ISv9Z4aKGZkuwf+1DbwV/4rB4Keqg7ky3Xzz9nCuftvJroaWZleoJmOVxSmxlsUkfP7dAP7rMkMQ
kU+aK/NZo+xlORZifDWS8fjBBmv4BCULGXPeSMfgVS3ME+x8HugIYewBa/gLcTDilmR5PP75cJdV
EmigcKcsVmf4cWDXPwV668OYjZxcAdgvi75w2rWqaSJL9puMVfsTYlXwA4n4UhfqYbRt0njh2BL0
capmqWzlm/h3EOPfnCeoY8C5MseY4T84obE88nhavF+x6v14Hu4lprSpGrxS8MAhtEOxiglIMdR1
6x2w0PaaIg3AVbdK+adgpw5QS2Y8OQoOwPdFMzrkRhV2mYlwewrUi8TNafBC5APdFrn3cgNcle+E
HggAk/PyIHUPyBCf/gvZwGkoizNJobLXFcis56h3y4bo1qvFDoD6NbdegENOD3xB7V1oblJpdAbR
1vTXVGxezW3h3sr0tkDGOtB8lMb8QVMG3TilikjHBte+7b3oOrum25mlFUvli8I6eYLDZaSC/NgT
N9E4lbnRBQ8mvR9ahWpeeESLfEFQk7o7ywohgWjKBboFNAwfZD9tDTuKSSUJIg7NDFuF4fTG503s
364hTQZx/BRF4jKC96KO68L0BZOVdULdxiMywxbB+3XYIuxjn+hJMmgw0H5/28IDBU/rvOnzCE4w
MFIPKgtAMv1AU6FImplgT/5JzdPByh6QIO4q92piA2RPi3G8PqRdpScY8yynfWvQx2TRRLMDoFAu
oIzAMEf0Z0UDcJrXyR7uEfILhieHYajQNITpfseScuoFlj6S5TQLU+1SuEbdcANc6Qw6gxjh6Pm5
xxmSX5eEL8tQZSaSpXiH6921hJMv8DDn5NeY6lC1BYwGlVUIOm0ahK5LJEu5srovGl3/esjdCrbZ
9agMT+WuxzDAYAz58xJR/24o/zWaPWZVWwOjGUzbp1IvxUG6dkNlL9B2lBtwKRbAyTEGsFd86eF+
aVC04frdfIzCGNmNSbFqzFb7CSD9qJWroGuLU7GJOz67HIeAOpJFp977THQlMBXSJF2hLCwf1dEd
dDD0hXWO7nBW8XC0HIQvETPUeOwIjuY1OVUpG8oYhrrp5DgmigRi+CK4FYKJvRuoMIlrLgoef2Zf
8JJbxRUd60GK04duvfCrp2fmeaDa+7X7S7avka5Cj+bhxOCAqCUD+9NMthmECiOpWLeOemkz7BGO
G/Oal+P0qXmNwSmJSyes15RAjpTv69ZqMXUQ4TX67aSwo+2u9UOk+4HT+rKhPfIPXoUZ8czNnIIZ
u8lYj0A+WZCJx1PEM1HC3QHAPp1qLxVPYeKNMNz1sTc9SZLNm3khpcupVjeO9xI/4v9THYdilqhL
cYx/4CBhOv3+kC9/q/A9NC6JOTw2XM50Ek6YgQ8AageVRx0fSKDu5RkE7WAFO4HsvVAQ8qvTt692
IuMAbsOXuTb0VlUEGTWXo9blmSFPhDBv7ohfPZJSHmRlrMxpTY8x5hwQAutZJXZDqLb/5sG8rqFP
rV3h+eINZzDP5+A8xeltC1uk9AhhtNCq2qLcO/TNy92ji9LCs77lHStttbHKuymxM7EZsph3NRn0
6y/vwMkRpYZ+nvXXd2DOnUQ++gxUW3YoUGqVctSOXR0YUF34nEfXNvPbtHDCMOfeorMLPmeyhk97
2iSueCpWbmukrHjHq1I6vdPVCjPjlFMqvyOE1RXuH9i3yVlqWFigQb3ppAuga1vDCLwvohJRRYs9
hDc+tWc0lPsWYTCTtHmNObXtdlJrsyTWNYEJ0PNJ1watIWeRuoFICf9ntE/emznGuVcwH7bI6161
ON3mJSiHhWiividjJjnPchJP1KFyKl+ftwnsAhRG+ZbvfNwLTaZIDPWI1OHIHgYvVXjJ0ZeXjywN
F41jM3gFwRRJxzVtJJ4l5voOt0vF5h4EvCJKNf8RIvaCoEY9Flau6HaPVP7aTbFSglDKa1Xw0yvI
ymzla2A4Ms/93OkU/oTPA1I/iKfz3akPXgxzzTC9IgpsKIUoDQ8iTloMySiNbyqkqcMtE+juY/5E
8ZjQuJzqW0Q/Gwqpa+lPpKaF/XW4TZBA5qHqTBbJF74K52D9A1cU0hHeeFfPcbPVTozDulwS7DzZ
rcJIVgUVzixzbuVnq/6cIEBuJlJMbrRHH6EmNK5HWesaE0hS0hl/O+0JRSlBM8BkI6HMv5Z9HvDq
teJGJXtWmqwWCP0roX5ARQ97jrZm8UH0pHiwbux6IVluv3tUaBod+3f94x+aG3v9U1BN5f6jMQzt
489kdPGQPazFteT547X5hh/dJkbSrS4rv5iLUCtbTL11Gzr7FenNpUg7e2E5tRp3uwPITYvhjeeE
hYJsYkAmLp2GFpaH2JY/gcpivwAQcTbHBpX9uv85n4gY8nyNdBMmg+Np5QJABSITsIuwlNtodV3+
5QddoPEtBU33wkO0HxOezvzojOxu3G1l8192kCsDOAXSL1l0nZOGgdP3eECaFP+U/St1GPrvaHES
6YYOnEHqnsueyUhtnAiwt6FcmZLrQM5vgEdmQ1vS+IWWgXpFoZtS9Wlu6OSc3OVLyrawAxdVfrB3
BC7wPUAG8e5gsso6pZxKys+iKkBKvDiMaiDhWNYlnePq4S8Zd7HiXpfxcY8GGUZ9yZDQxjEBZ9Vt
I8o/fjy8a0X0ci16SOPBVMLfPW3RHl4/Koh9vGH60I/NiDv5Nxi3Ox91ZDaOG7K1ERrTchp27NH9
CVUZAA5fCIW0i+pV7o61gYpn4/UooZJVVRH/KDRdPfluVYIIMbqE6ioNVTyXqaJ9iSHdNjP5sZfg
M4Y9svNC6ZN1zTo4L1s2Cmw8pcnNqo5eYpvDErjKdc7lvbc42cJ9aB6alwYWMI5WrMuYKIg4FtZl
/qLjMJZUzqpSu4XoVlToiCmJzN3SmDkgo0oVO/ob56jLPwQFvsjKENLVeB8Du5sUIkBmrLs0Ohru
YjPtPOKeZszpGDYIMYvDCjp8uzYL2a0/XoFNr4921D0DrXKpCjs1Dq1/5Wzi9VEH3Gp4o63vT+Ny
pLZbTaZMMJQ1PQxSOn6oJIXaedpbZenU3vSSdN34Gg8UBtVX/cEVbrgXMD/07+H2wHqSqgsqeF+2
udY9RwrQiVuZvYxuMSo/hzQCG3jLgoUo3c2tHYowCPoBO6vonOTrLTZ9QTaTY6hufkERjq9b32sW
4CGiiO8JISzmHSQkK/Af8XbLrCUBUnKzeW9s7FcPhT3mZEdG42exehlDCDHbMmD209r4E2tq/51m
d8Nezlmo3fS/ti7Xo5ooTO0of7EzBxvJslNaXSP2GRFle1TnPt0078LxEFpQid0yZvIQyD9OxAjX
J1RSbZcmZOXt3Uhxi7MvEQigx6KES572IagvUN69KpJGLecFGqL3s+Cc6KhhPD2YRZlkg46btrHD
0lR5zTnM3eSU/inQFgu6gCi9LB4x5ibrgac4xKd6XUl25PHY7jU8gXXbmuBsgcmVyZ8y3tpNE4+a
z/4GzEVVs0OCIG6Dyutcl2tCqaXJc40uiNVZrUmFd/ceKyIB5jpOBhvS1bKiXKOo7oRUv4LN5hve
UE65iyL6xl3jaYiJxAY+W+jneQAtv1fXQnzr5skGbv01xHEvM2asTMVoJ7v5W+H+YhTpEYmp+BfZ
B06ALOWfmGgeqA+opNLT6YnE45iwYEeJQ3Kmjh8PIHqii1krq6xj0tLOydcPuxqwSWF75u3O9wUT
fdPLrP71pjAE/YM1XdWW+7Zqw4L52dhPlKIcWe4vsAOgRwyehIST2w8HO4H7N2sdUlCZn5f8RxrC
woAcvpCGsSWry9V70rddDYcFgmanQEGBdUatxFrdO7TPGe8OFm+/J5zOZdV6SMMgJd2PN79+M6VI
jWx3oMfUAEVRpTCCpG5nJv/j7DCgBCCt0VFzIfYLwhTttvfQNDq/xLslktPo1jGYlvWF7Xzr1+WE
taLWJhLxG4x4woVdsEGho8kGmX/oX9MsyfPFHB3Hm0MEXc89r7KxOL0QOpl4ijxjkRw64tEEA3uj
bfX7wtZpGmQCH+vVk0FWWjj14vuMCP+UyLgW/Qmf4xLaCOZJPUwWTKIFtmDeVbKvuLnAQ9jPSusA
AMfrIcmimdI3IiDzXyVM5w2B5NN5aA0cUJhhe1CbU6+jjUF1ChsOZYAOKwh7wplz6lGUEN7gDTlm
tAz2/Np1VOGsD+HliDYrPJ0VQz2PWNKPn+eyOdZN0T6Rxk4jGNE/ROukYtTGIMkyUHwo4zy3HOwK
PV6iYzUk/s57BH2uxyOYjZYa9UzZjbZT3GrCHfatezB/E+qolOYAkf6VcupLULTfjDpq+UWRyi1S
8aiUlyVMU27nIkC/xLdIG9sZLsJCaLV0sPc9SpUu1KVQjugJgkHgncR0RxKFS+/fAh3O3S5kxqMd
eU3GO0w/J1kFOSN+8oK+Znkm0IZSl6hzNY/WJSGsrZ8xFr0h8wEoWCdgDKQ4fYLvcO+DUmGyAv/W
8PNoEr4VZXo+ObfbAO7yUCSB93e6lERi/g8u81QZFDmQR5OJrg6nR0KYYcq0HqAKIDH8aHvvfkhc
iR52ShVj1ZRvZRUfdb6Po7tgo4be67dS/1aIsURoGT4vITRdTbYME3hbgC1GlXYBxqO4hIq35ndd
NE0LeB3tY4smSxkwRRJFWcY9KE5NK+e3RvNB+54LAMcO+VQ0LyNSKouJhmwSfYrRZwJFHefJB9T5
oSD0sn20294AJ9zG+SfjsrtD14CLAEW3kik/q0UvfWGl3PHIy/lvtNzoeJo9RbPfjGY9WBlLOx6d
ycE1yVeQ6C2udS9bsZSyu1T76t9AOAGeKjqqAJDcMG+W+6pKj1OEiRNXIYkypjOejJSLis52zXoT
tBMF/WP4fpIzQQWOklO6EkMFBcm7JrzcZM3SPaFtaM0F96ZsCICYT1jlGvSW8qqhorFGZidiy/7g
FaSX7rH2VYGnLHeFlX3ek8fuo8tC7OI3z3eA5upURmBYxMSIvlJtCwpZXrdvBJAE+T6NzGW61yIR
BWj79AhwHHXnokX1uqj8m//kWGyG1jbm7VWbGnfCuGV2RCIfcyZxM/Ih96v9WQoWnz+qdBgiJq9v
ylqJwZ02R6vmEWkrKiT+XBINk7UpqRi4aM5NJ6QtKoObyDOhkWbQjO/x/+veayuCCEMmj3amN/Jx
60xNm7CgR+tQ4FQGtVQdmm11bldOSmGGba3GzIaZB2gzrYUYeebB9zxtpWVwUjbxLOhSxe2c8SXO
U9PufQyuFcshe627qv3z3SKQviNA3zVV8n7pVivkDpVYSpD2UKwyuJ4Qug0vv1ZkjBMl6NAyEcTp
FPV5CbmMLWicyFmtitnppLPyI6Lx5wTTKobbjlhovjECEOFf5oF2F/1M2Q5urW7F+y+45pNNocfY
BC5I+fXB6AgZ39yUWLBK/0UypiYwMFjtMx1rBTldjGh67RGsTOlY06YnwN0TdN732dLPkKhpI0iI
kZET8hYxZLXaaHu/0Vk5c8d4xrkICUtp2zRAnJtIpDWMoDt2m7T/V5Rz8D3yoi2mYZ772v+guyfo
ebKE5To3Qo0JhacPw6Ys0P2g8QZMXzvKq50qSFTBcJaYt73qoCaKs3B7lUUiveb60wEDOQQOersH
BxGiwJ03aFd8MJoZDgbDVRSj3k8mEqmEnQR2mczx7mhze+aR08IfGJWxvZZvW2pWtanZgAhqVIvi
peHkYTr3A8uOsm2zBot5jAFkDmWsPu7xCui5krMVQcLUym5u5q0UC0CCBcRGcIZlbUqcN+KU1RdN
1j9JjYB52IF4VssEOfBY8foW5vbZvL3R7JCuDk13qHDncxtX9gc1Gb/32pjgZ9PwodXCMi0H68kP
px3oQ7PwpjDlabdUexOGMuhAnS4FtFy0qQyYbhsST43X4UCqddnAW1H3iHVLYPreyjnxVtF5OoIb
JYWk2AGEeJJrKEIio4mUdwt9ai6qokhRZ7dbA0qRQY+NZA3qz1/eZrVFD/J71C1nkC9MYNi7q9/+
D2bmJZr8aEW/bsbtPIZCeG64A1GKPrTzstBOuTUyxbX6sT9+RxHuki8yyqxzC5JKmOHaqlOCKOze
IJkqFfbxhmKg4zUzv/rniOVQTwksOJFZoXHvI88ut34s3aJ75uysZNiC6oqXurXqGfsohpewDmB0
41+OH3m/KBxIMwqwiOG+aNRGMivIIbQ8vmOBIG1yTS6ViGDXQ+7p6eFZtM/zEEMhkx7JWmmB8uhG
dp6G5dUJDTKglnvL9G9fqV79TXUOQPYLhzdkPVgIaEuPFdvEYRnqPzYt8a9DJaWP72Zxww7YiHMt
eKyiUcN7xycksLNDPyLtCDRUJTWKKaL3w3sV7lU3BZRf1/w+Z5qoKxNj68GP1yDrU7Ckv40TxM3s
Yk10QaKd8FKM0MQX2GdNlPzNfM1M1kYklLQIDmIjczjUYiD8S2OuEvlMdFUxFwdEHr17122NUVsE
7OQ/GLIHrFMKAKiBFPCRImvKawT3DCU0AG4JDFONv6UM6/Re9qT/9UTi6zGQEzw7tLv69/cSNwQM
Gasebg8jmLxUrY8drB98GD4koyIR0iKIuYn4ZGaFuugM75pQXZkkLOWf4ZxHdp2icoHecvdcTIEJ
RACMtAEHB0Fzknw++Kxdr2V2hsSl36xQJjP4SRk8i0BtP2qteDObYzjhreS3/pXzY3RsfTMSJTwY
SsYaIUSg5+u+7DJubKYEIqJFVuJRFUaYaLPfNqkm7eJfYPy60Tocip6bRTsiOxIhY/8EzUO+c+TF
yFBkHZtcwD6tMSN8ZbUd04dmDLYaByEB7x8yoo5NUpdZ64bN29CYBOplzxPycTKaqbkHgwiq6bgf
YoGZa51SQ1/ehHbpJrok8KhEnpKQF/2bZ1XTDZ16GG1+AR9WE45Mz9BMEtF3EjHpgn4xkCA02RRh
lbadpcFXUSifsaGvWISA7h4TXXkRGnTvrwK6Xgw1/8lWzGZahznNvTtVjKiB+a/ufwihCMbDdCi4
pb1yY4IRwJas5GrvIWYCOcjKd3+mM9jJytNixqsWs8k1ta1ayucOM8clzfg9tvIwFW68Qf369wG2
763Gmqno5Pn/hSU4LyZf2cJsaqGgTVx777IG4+UiaBMV7FLe3XrIUSSumBwR0ytgFFVlMwlbD2AV
3SUjz1nee/6YcwjHwa5yQRGRw3YBRK5m+xW6OaIIJU3OXRXe3FKzbU7/C7JHwSpVd8ji6LU8t+i4
5yW0l6ZTgtK42hBX8azT/01tO8zqX8ln3UummyswgVAa7aqykSI61xbcS/3uVB1TkdPmVzeoQNEn
poCHQVRX6UCJm7tbtz3SKGgWBxafrQmcNUB2Yc/o+LkZTh1EvTp7wMMemQhRk2NfoKIG9MKrFSKw
qHLNNYIhg5LIaLVwJNwNhGYYMESchI4gCMLd4CBM71VlKv/g2sWB/vjBxaF43r8jUmEgD41W09Dv
+z3VaRqoCJSVgwBUko1EycyA3OXi/+NHNvVrQuENJiU0uH5jfOBmy95OYYcK2au1tVZhi9f2NUB6
GFJhQh//16eMrv5SnCEPmfxKPsOhcfI7ms+C+Bgg6ypfZ2PF58CYzLlJxk+bKzhdqzDI2bh6oXsa
XR4Lkrk3PqNQjbA3AkO3jcTyLMxVGBvkUKVko6p/0ycb7Kj/UDeuKu07uHv+KKu6xNsbQwqPNhx2
GLQ6uwE74a7OuJqsC+hwvw7JbRPO0x8tTvZhTJWtE2gj6LBtvV9WnXoZfN0jiJWDol5OCe84anBk
UzeNGeEl0hg+9lnAp53CvcG/bKa7PvBbY/wrgJ1NxKaRuKgUa64mN1kYGphw8QlqoIrGb+1/eG2w
HB96KIQDRC7IeesFqFLnW1PGE6fop2WbdWBE7ZnhV3jDXR8EqeINSTX0OLv8QsIg9S5Y5ToBvr21
vEra2r2OFJxQNsbB+RhwZ4cXay9yvPhO2JnyBY9IgAm0LOy1hdwdrcNqClNVjFQJxrs+JW0ljXs8
OZYyJQPKEdQqjIdulqDC0Lkzsyae20FX0XaTFIHkaMD2nSsatVpIOcCSkHmQ1uCRQWTkCpp4h34l
jONG0mxz8gRaAvekuYSI/Zfbw72tB2kxdCJeLFUAYC7fHyIO/fuIy8RdvnRX/fef19K6oh7LvRhr
RUiZsl8X0+aLNFupbEVE36+nU940zNcQmJuvoeO6K2Ud9OiVC5FHnUyf4uDvL0D/YarpopN2Q+Q7
/41QL43k5+rUXR1FohmKGW641npbCuQ8VunwuV7uiUEkvV3AfETO5h1a+IQkp7zcB4Ajh05nY3up
008vAWBN3xiyfFHzGwjE6T4//HLwF0MJBZ6T8HwA/HgtGQzDesMxZzNpa1zycjMYSAww+yC6M/KR
/Z6hBcBcuQi0Ic2Lyv1MwWaOPiBWzmSdDgriaI9DOtSoNBPy1Rn6NTVxNZLZU0M2sYJmpUdxCGVc
V2NcoFeKpwtrGpSipTeuqM3+HuQIGaj57gtz34ddi2lNGpn/JOyaEkP8UEyfhP4aM07S5FOZoYkG
Yrot6pFuslrfbOL4IbzYWCeYvV9HlqxJRYn8sGHSLzkTK1tOQMWpbi0MF8epKRtcU3F2sjz6DhlD
E94JXJQToaNtwZQtjJGdwq9kXyFeRMfrpWZCHTnk3G21jbMhaiEu57ho9gByjIZaMGojfm8HknPL
VNm1MPJFMp++gMaBVhXO3zeRo2SpehEvlqbRvYILJ3zCxpZJX9MKfoZFu1pMzm3L244m/LZto4ek
JlxJu9px/9bOCYz38APwwHaVMmhw8OjDuCXRNo259w1ejD+gfbFPvT7LdsF/M0z/wevxiy9MTJoV
3j4L/88Cd4c4U/pBwK5GR6gtNPoVPyR7R30EZESscAl+q05iwta8rKKL75/MKpB3zqw/tgp4khQE
g65EEtxELuiBPoAHfF8u6LQnDfEi9jzHPXzYXgokRKOTT4iEbaXwLJ15cmJacpU/b1JdDQxLZ6YX
00AKL4D/MwKj95lqpTpFYS6B+1b0hLGYS2luIYtGNoyyK6yMuocrzB4Laax9q7ehUTLnsJR5OqC4
SbRr7kqdmO1eyfeoEReW5R3EMmetGCkdWKkTPnjzGvcZcayOUS9atSGf7JRC1l/ScE4oz5bPTcTa
14cLYx0HDbK9eu8gr7eT0m3XwvrcqX+aHzI227MAa0xNBzsyeO3g2/m8BhKMcB5tygpfXm4CFLHO
ZzsWsR/SYLV0FqLJe47pO1mePZUpfvlsE8pAsQNzenyQxWGmfmmZwDlJaKhAKlSLgnnJLWIOPc0b
Iqa7v0n59/DZwhA3vwoIfcbfeWTeIpbrf1rnCXhSICWH+3IpC4Sk31MHQr9VdIjohxCK3zZtOK0D
ZENRgBsgBbZ2bkUEJ73gR8niWMtf8auxCDRDSE92ILtNIles7xuyfkQ7VpKWf4vgmaOkcdAvbOeu
peeMug3icx9J+l88Rd6JcEJpxcP/cVAYlGMmqC0l4DeGI4YcKxjh4qDwtscVVUlnlTkzw0xJzoZS
9ItQYokowXW0JphrunzjYhHw36+jTnzqRwGeTsfiviIMV0j5EHheet9vAWWe6yFy0ymlrJTm0f6B
seIsQy22tCkSgMVVK90n5Wz+/PQqqtJ/6KNGdWcTLDDED8ZayHTTt8TjLYSXJVUT6WCZAKWqRoT7
B1no/Nb3saVsztXvHqb+4esSAPFdMoW/yjHeom2SNn6zDpzq+QsgDU93w4TJtS7/SQ+ULXj2lXmU
ofbvXhpXE9vxM/+viKrshogNxYjHSPJD5Uwm6y7iCfoI7XHF6QsYhrI76qGFcLRVJUvjwGNKFh8m
39yM3Y27suN14y5oIdBdDINOn0sUvVZh4vWFDcK0FWf5QIbfkvPp85VhlKKiYdfdzOCTHLXtTo4Z
BuZXUFsknzSoklxUIyrZiwSWUPZfPswaOoWCZ/iy/Cm8GtKwZKT/jlZIZjn02YAm4+OEPqqZ+ese
35VEdn/OScGfuWQKZExgqm+ysGPMEuVehehPNdPwqZml0rV+zVsNkaz+xgjo8+JPUchAlNj0zLm4
2B9I0RaQW63OoAx62k21zRPL375x5w15QS8JalYSTqG7vbuV084zh8FI2YJtu3RHyzBVDpRd+f49
KLtW6tYxBm3raItiiWt3vDXCl1lpu66sJAT9QhqSzbQ/FKm1kKjtu4zSGqOgSHUxyyEONEFz9Nnq
2achQUzQiGuPgj9eMf6NPl4PJu/xP1Vs8+DyySZ9q9jNO5CWrXs99wjF8fOrsi1doeGxJTXt9j3r
sD1ryu661ECC3H4Q07epHKSDeXeboBv3ffgZwB0Fm1g9Lqxc5MzrCbm9yFhnruoqrIUvViPTnh8p
YbIoPBLfnRHPFzSS0rY438/L8xd/3qjKUE/7CNvs1BPcOreJ9T7dqsdJQztJmA/1t9zeBfzqnURC
I7WZUcJD2+Os5LOhhrz8hOhxCekkq0oH6JVSVVk18f2A1n8/qxU+iJndqVxTxJcCLekkCKeQUVq6
mUPa5zns6rC86bqmR32YD7jdcbnrKXhZMw0UBv/+6/GkkhUckIwMHPWfUYcYdt3J0efix0xqV/bH
MMfqvPhQVlJGZX18/PoXJKOyn3MWGlPnaQWI87hLTv9NfNpRN8w13hcw41HUbJzQQWyWDcfxwX4W
jZA1oJ/lvy73cKYYbZvgFqO1NsNM/rvkBkifKNS+8EXkleluksn9J2B/T6I7dChG3bP6sjqbszo7
qtFUJ2m4qE35ZGWCqstOXwud2a176w1Ac+Gerj2+P87kSTtbtoiZCteNOEcF73cj1swoSLGjE8qZ
0Le7+2n4BlDims4hI3yg9m8IHWED5GBBrDlYlccZJk7e1lGFTi6bqg6lbMQYH1MzfE+9j6a9Lh+0
i03RbywUiPLMZifYmR8AOJa9qNOPByv98DDmUJ/Hr0s7Xrxd8PSmyLPJD8QiEjq+Wd6793OcHjHI
0QuwAF3Kr1pV3+4t7IhTAhJwxeiZ62NSGktNV+0WzCROa92UetEIZATC8wJzA+LmTdRdqUvw7CKT
k+EJcn9JCGJCA2PE5fLCGAPMqmRxD8S+K+/7E4ztxS7Gtjs/XsCaTmB26BP7EHrInRqQ8sPcnhso
WNrWxn4Z12aRjduzU6FIB+v0ZiKe21cyibIHTDLhC/8afaEbUT1NRGbKJKMxKnaZno5isjhj1NAv
bTgRPP06mLpNWgkHrp3AkYH5vSi7AmNGdWU1T534GhlizpcDWfe224n5o+LMaicYYvo42hwWpYqw
L6PKpvuWSvtFjtuYNQiPfy3InWuEtRi46CYEns9D+LEtzCYw4cMHPkSZEIm+A/serLgptOxKcHts
1Y0stlg6QRdN7B1K/fjrbz/93uvc6ITNIEKIeBR8274M7dWjlqkqSLI7CsiZY/VB5/WPkD/1c6AL
T8NvX0kR4hFFSEYylG9qN/Y4psee5rkVl5GYd2zkQp1pJJanKnlqEzh6OwJ2CmRZnrm6isYHfQbd
316Lq/xQe1Wn80WbBzE/7xhSyDG1oROp1f8gIUragzKJaZiQjRvoXG48Aiyk9vpUYTzYRNn85kjW
UoBnIa4dPdV06VdTzfDb1lnWPsL0ByTyJv7X3fD0Aqlu5wdXuLNB4wTqbpiU3Yw2tR1qVjg50tqI
xQMDBWkLR4dAkIfC202kDGqcJhQkfwIpt/dF3ykQXaSh2BN2T2SQAifUPwy3zJc/ArfUKaR8jCjA
uBBxsCxxiWgWn0sP7A15zrsL+HGtjsYHucIdJIZph8K58P5/v5Kj+xdfEp15a0CGQcZQdr4Qe4K+
AuYvlKrxNun7hyRV2oghi2D4REx4iNN4eXNtOLt2/vv95TykRZl4KP+C+k5tWJH0sjcGkHvvlJvW
bFnmEyuK0C4F83+MUNdfFOFdBk6BJcJUXcozRhaOucDi+qDt1qJWeHp7ncz3x0wJl9d+hlkz/ZBl
Q1EgidwJYW/KFPIwXU7BPtS+KbnpRSp0DyBGGKfsi/ZWLNSpHdbXlyC61eni3uPf+Otj2ouNlZGW
2pSDZRrIgH38W1mRoGzMvmaHwYYQ2Mh0+jqmtuglpj3QHKsDUrghzHPIT2AiCmJUEyed05iLqaiK
ybA1oTpM29dLU8hTXe8E/xlR52vilb+U/fFbHUfKIKEa3Ydr0MDtIkRjwVWtpxwZs73+DmDJGrFd
tavb8MnH8XbXI3oCEIocjLXvSMZGVXtxpoj/WF3RRUW88jduaoyuHSyP2uJn1oXLKTj8jm8neaAt
KJ3HPNUwRd24JCdm7i0cqtb0CpMudm1pMLUm2cqCjx8+RHtE+OssVCrcBKdg7uT8LY8ojXczpjXE
/UToFBdHco13HsUKuGW7eNxg6PKtXdIrvcB4KLhIZch97MlsnowSeA9JHwu9IQ1nlbtmn+46H/+e
cTCMnoJzObDGg675GNdZ34MAZTsU41SpvdXN65+C32U5iDvC3g7VlH3NtX/IEiSsD70oyX3F+EXR
symYtvcoCf5uURUsADSb0e4bXZCY+MS5uUPxvcYd6IruXJ9okGFeOAYNvKbz1TjHHGu037aHxI5a
WpWn0Jid5hDG2Nuc+OUSUcby/8svtOQ08aPGGoolH0YVvSMZtXO5xhZHsGwuTyZdDAIFlF7Py7EV
xvchM1+N40EyHi8I+gJNRPTBELdVRn9V+75E4Lt4ijtjWKI5Gs/wfUjXjdGjbWKGKk6OyMDqNF7E
FQXOR55cgrqhOmZ0dUaS7tn/jOSVaYCrxhOCpHiAAZAzzBRBtbqij1/5DQZzS8gIDFN853kSnZiY
WGMX2g/R6wIig3t6ETWMXGeNRmoise5fhtIEB6Ob83KCTc5VWHnDGR/OF9SsF6BUzBNAoJb9y/1+
dPe6JSQYW50Gt8bUxWY/Vd5WjPwD9WG/9lQzVzv2iAocjj3L3TkXkpZoFxvtt15O1vKkhzC6eh0M
7KZ2ElQi505JWqr/n26oh6q05y4qZRSEp4XlEU6w3BVnz72riHuP6Ua9dsC7f1RmypjAHZ7XkpPB
hO2U5K5cY3Z3NkXTWEkOBN3kM2OX4f9vGQ4DZ1HG4vMrn6xnybe4OtiUDTUfsP1xXnYVTRL3U638
qj7YUs7FX3Aod4sT0xe7G192kPJh5ESxXWHpWGeGBeApCIIMeNrsJ5ECDEnifU4K4JtMg/AHF6+S
vk7lcCFUUDP3OFBTV1obgWTrxR4fLN8rQzzSNd8FPlpOgOA/RWnjEwxPwefk2/gJgNHc0Zczklyp
Px8E2pKQ5XhwpSrljZyOi3lineDMbnAVUGB29oWifCdJmKGzEXb6GYKOetsOBP5sxa+eP2Bc/asC
C94rJa2RJQKDl8pDFe24V9ngNoB2TGuJg4ALJnF9lu+dEEDOoaSbRCJREBFcWgM4Ptcshry0LkC0
tGgF45QjmkEqV3js5GaY2v+caO5UUkom+Q5ksboBSL+kG3Mp8VX6e0BZ9m+nIGXOIJioMICo1wAk
oCvUnD7peiSRYTBlrQ8R4mkmbSEflOjdFlhIKEX8Q08sh5TAs/+CwP1OHPjTZYafMsX4oE9iV1Pz
+pd7duZMsmySPFMYdpZLcXkjtotqihB7QP7Yy/2cUETz3EYblWZHsiXuJ+nAmqaq7zyN3ZEdZ9lz
otgI5oKawmA+5j810oqr80LwYOBGB8cTM9htEZqmZCANjcoUml2szLcO2n3t93TGiZpMJnuiXcvJ
3H+3PkJ2aij2KY05Pd9To2i9JyPHqZhlC64/sZznDHhvXT/fRwDEbbz4fB5/lbT6jJfcJq4BH45d
R+7CGAbWRB84oXNEzoUO1VPm6GDoQDwcfNMpuX+GDOiv8zjvETHitzVX9YSs+CUJVy8vhOqisVYW
7dmKRByon56gaOfiIXXA+E+4Z2VsYpgkE3I2lWjEeZhpLT+4MOavgm2LH7GOCbo8uyBaQXii24fc
owHWwzyO2ZF+q/jri5YHSQZCLZl6q/sX84nIZaQ45NXBRtvojoTJI5dv+iiY0M/rd523NZQ6eJVI
kqYxycReZtnkruc+2cAlWvzI70FVoBW8e+1GRArbMEUIE0rO4PyvlDhL/djdAVyOv/vMDBikj3f7
Lddq6itVIVn51C3PUVgC5jGUZkPTfkoAxd7T9loTMVoGio2crtg2HbOjwJHLObIamflQ2ptw9ywa
g1pofKbMJtSssm5oNWRmS3WKaEMBZRafFM3nW1XGClAhreqwYpSpLSjJtF1Emz8LmDaLD1LHrwM0
fwLWrpWsC+JeFbDZse+AuDKIg/5Gp1wBHy7zUSQdnPmlqd2B5qX67qilIR1fLwgeZbQbScfJ25ZL
2hDPVdZ37aogO+FphCpXXGFPB+YdXHi9dgDsPOeXldxnMIOGnPicX5RK54wmbh4o4Lm4uH4DB0eD
MNLqhY/oWXcpOvRPD96a4PJpeHoGM3XUmbAtIWybVh/oWHP6EjqLAd+81CVo+B2M92XtsBLNhliO
ExY0j0tCtN9UBtRyl7ONscY6Ct0Ki8SNnnbWDY4Os+Oyi4zEUjN/b8E4IWwmaZahXM+VIHZRiYF4
FUfE8lX/0xFFg9cC7i9GkA0KCrRPVPPDOwy5ZSlWUF7QFj4RPsGGLYWkIq/gOR08P6NW3tmyycKP
1mK/pBzcsKux5Sc3uz0U5TAd0jmuXEzoW/lYd1wRY3Yc1SCIIlhkXgJCg0D6hIb2lTE4sOq3yVRV
whosyOp2NwLJWv9YEVLsAxKtZtym/MjIHfblQCNGDm2vm3w9hdbiwTAPQPtFkgTs/Di0pF3ysyT4
7F02z7FFzMm7bsqKy/c5McwZ+wlgAoA2w+O774H+fRTPyALRgPh8fHr894Ti+ljq2f4eFilJaASB
QABuEgKbR0GFKtdkvVVTu25cwi/NFrGaEsPcI9ckfkjocBGG5XRqUpA5NbyYMMnCL3gD/XIzUQH+
20h9JhVX9N6p4mRvXYGKbISsV5DKCOORr6tRW8jXqE9b49OJdsOsHXKlAy+Ss+FQ0wnDP7W7ItfS
xqiYzo+aBQNlAYCOEI0YgIuk3iAJDsxfYGA89zHByE8QyTcqb3ShDTy64nN2fNLJ2YzaYJ/1AXLL
6rOdkAJbII848XwaTkefwyid7LGB9SlmRLUhwncGd9dKgkh5rPtQqsZNqchmtyhg8LSQXnTnUZDu
qTncnfXS3FYLSk2XwZM14QJaBuI+NimCOEq70Da6J4SAxjTbOVHShLNo39UiXzjR6+nwbirrXTXc
GXNHSfzjPMATp9GI+QogB1ehGQCiNkRhejEJT+oBEDkvS+KnbsrFXFClU+0WVHbcMBUzvTvau4Uo
uGJudCtKkMcBv7YrIPCtd8cfxVtVf6597zO7eR2QjZFnj2jyPdRDDJwjv1uoAm2yGNzMjHpWmjdw
Q+nL5ovlFcWQlpF5AytgC98FpmuViuT3sMP/aDhjUY4CRUX5w0Y4CzMc+UaUAaGUUOL489tRM9im
VE7cdXN1vn9easTPRh8hF0dJHcDSivZeo46gsnET/Usyf7RBnxtELg+Mr1fsmUyJTbYacGMMzyyn
CZLpE7xRvoAOvI50Gk7ANBO9FRNcacJ2n1D8Nn51a38qt3BD3kOKKc71Y9tfm0PgLLZQwMs/lPN1
CyUvkjKFuIShQ6DltFqzha7Wskm6+LnnEZHuCxo4Z6VkPMo8B6Y0KZqMdOJJz2dFNCR2Pn8sQ0Cu
s7Kx8v6tVxrUCry2RPnmerTOb+qQ4PjSO2cA5LK3N4kXXo0nyR0OhzZ2KCjfzBN/t6kNA9/8+X8X
cJXGXvPtRjE3h0ZOS8kHHFvmT6gY7uuZ1vHfvj3gQXAn/4SnXuDegVH+Vid9duUlJWm4omSu/F08
ZOG6F1BaSz+L8drISrAiEmPHGsvF98paRNBs5J6IlWAaayL5cyRmKeQuJN0DVGIymmRXp/uzjQKh
2FfzvcrK3D5dsI6xZjdzCXVNcHVgLz/RD3sKpYsvodpR95DslGiCr9YzLt0j7bPFOtj7w1V6Ubcd
KmBnXsqcMApnjmD80x1/otlAgJNO+HoaOFc7+CO/Quq38vDjUOD3X7Iv9dlZFigSGrtvEErzNqL6
LPgVtOHHbU3oM+IbdJXEcx5CTxnYz1o3s6zeZJExrhLAfYzqNpqzpsaa3Rs3f2byVMjop8QrGDT8
B/l0hF3YiEIxCOQm8MJA4AY+Pf7/GIOx6ls4S0t7uCMy8Ipr9njOjBJrqsRrT0QA8mpByqL2/jcY
2kDLK8442MptSa+JcOlXhltGWSJjf0hHw+rx5U3OryfFxlFMR7gU7LYURI47c4bmz1mnvnyUIV/l
Lpkc4Uu6ipyxSvrgj4N9BT3Njd/BPak0AhQfAnuVZnlr0w0g/10w3lsJIuAwLHGlLkdBW0o0mhjb
Favwgke/Vk9GYLrI39OZx1f1bi8Vt8sWrbESkFfgSiKSgbO/UIwF37oUTFhamDg3hdJUz1azNqx3
CkrcTGCOpeN2EPp3o6FAcq0VEFtt8OoLrHCGl3w3jEGWKXL0oO7fMRtaYflnXvCbB2mWDdt9lV7k
46I9rDffo6rVtrSY0HQFn2jgoRUyn1FuSJ994ZsVMAkOTthnWqn9HPdfN07rhzuupK/5/e02LdhA
49fg8tSGxYCudINxVyASTEnk/tp0Xfem5NUaVthN1XDxB60xfTaHna8zr8BDddVqqj7M4G0CmWuK
G+lXfkWB/rvdzK42qpeLFBkdav3k8V+Ek5JYOv0v2lE0sOEH6vnDpD7nCoA0We4B4ROUKX6GLT5O
UEJc6FLyDcmQG44WbyJzrx/xYZ/pOYIz/2SKvAEFYoyk5CixiLS8qru9KF3xE32GScCkVw9wyZM1
/8Y9zuEP3ybgAcXQd39qx6ba7fVKxWUaapJNuX36/BP3my6fMPGGXZkRwHXVOjkwrenI2HNEg5K0
KVf/BUr14Uif0pG3xi3mnRI7wh82EnaPmlIicCdcsRolJPXu2gGMjCwiL7/pGn1SKhFrUeYKDOC1
kqgbA6JIgN7C6JFxvFfnqGjk972DmTm6gxj3NQHOpqD6Zm0iw482O2Hh3EXZci4vUD3tpszwVSl1
aa/rUG/5qcbhBCTpT0dv8/XcXgaeD6kRkbgJm0GWr/vOnTNd1Wr+Rzx5Q+4nceLEzK4JP8wFSpsT
0/GzsnCci/0kMzkfnBe/C4un6Orsi2ubecrlkreonnSr87vCluyDOtLE8w0ZKlFjOHmXvT78m5kf
HSUBaqm4e6VD9zcfbycB7jbyQ7P2PFKzKgbbvtFmEHLxz0l99xS+MGxySZy9PsGub3e2Dj5MbA0j
j2jOXby4phAMkCPsIEdu1D9wv9xzPo6GaaPjIKHWvrx5re3sALPejAPxmP/5kRXiKSeIWv8NDewx
Is9c5yVAu6ted8DoYisDOV58hlfN4bfZxRrv0Vrvnbx/HlW58p8xTEgabYSO9WEaxCrW123he3dV
X2Zve54J8zUiTpR7TrHzv/YzGNhosqUzMEonkb2Qxf4l96hje984GV9PEoRRZl30GBUEW2jZ+RNL
fmPC3zox+c/im3vo2xDnIBMaW+tuTt6hIyme0u0mj9PnHqzQCdAzeQuqBVnl9/Dn43ypdbRW0fZe
DvU1G3JBeB6I0e4wZV3uDKH6rH07wZptdZezQmUtz2e63GecsEkemgJNA+0uzotwcjzpzluUcCFu
V4nZATWs+3tiM/6K2pdOVSOz1OAtkcCBau0yeqneYfLhOJQ1H9hmFUl99wTmug3usmJOX4FmdhRt
JyT3u8jwTGfSXDL+aZvGNpaPHCQ+/MNkBZfCtMVBGbjrFzcu9yuUZRhs/LWjyj4z3L9i6hPxWxCY
hemf8pBAvljuDlRdxFFRW75hLbob3fTavcsAfGURNiMw2358dSZp5rEhTm7plKgsiWRdH8QHfGKr
r30Rp0r+8b4WOYHZ3rrKJmRbb8SVrpgpRe7liwipB3ggtAndshT9fBIT8f3lx12f48nOWE27dq2H
YQpGv04X9Tr3srG5Ntnr8Crn3cDvWrOKNYR2CIpfSw2rvFwf0q9L0RN/GJiNOvo9BbFb3HmjFn5e
G1+tioP6JFlK9EFt56MujD4WnUw1qNga276NU0Na+7BwypmDIDGzwxxUuojC76luaLx+FIVWdCGA
6iAjXEfgc2vQB/Jpxd/OVRO8fvuVpsgSCTkaSKraMHQELq8ftJgVAN3Uf+mPdHtIk2oDgnaUnBYH
iQdHt21PSL0FNmiYEk9N33MqcLZytj+evuLkCAr1+WIjP3skteEcwMiujArtbXK5J/FDB9YuEAnl
y79cVpuy5o8O/KI3X2nAx2kTY298h/qtfhBeZlri7BpggzxlWgSsOnDyP2yuLuuQYQ+Aje+mbyHt
4JawShhgfyXZVGxaHTLO0YDu4iwL4c4jPcuZpuqsa2OGtKSU2rN0pamBW1Jb8xOrOfM+k62mfNdc
POcoMrMqibbTcE0rR1TxgOU64agCD3p3mfYIUeDwT+a/5tfU9rYeDWBX/0645IBpJHFiiNUQjvjP
zMb2BG0zo6VDuwIoZjNO9w0d4mClwd8M50H7v6JgXqGQfhjP90FLznDCnlBACsv5aS56ixbLO4Ef
E6lcADvVTE2/H4UX+iRtSJbp9PkCBGgmC482QImcOskqvtkVgk19cJuEgajncFu/W2bDvbdSnggv
6AK+UJjRK1eAsSAWZ13ycmUV/rV8JQpcKJnPm3kNag1sd2BqMNh/QqZRKVZ7IC2W8ykqxV7b8qug
mKGny24WFGShSEE/aOQ7NW9EMGxfPluZcbdZRbONThPcuSlztkJUke85CXDN6vD9sAHY2mywVUCC
OKMIXRijiAw7w00VrZMuQlzGSIhuIc9xsDNRIbKhmt2uuGJLjxXtmlpzXGxgOS3YltpylT3d78wg
qa6CdizTWTkgQR5mlOY1aX1wtrAAEeuoosCifSLpA39s1igwvINE10QRn0eqiD8VyoTb4Iz2e0zu
vO8++VHbLtCrkSwxbIDftq6EVYG4TiDA7SvmJm2rzRHlfX0uK+lmqKap8oIxwJMG6JvKV0f+jWf+
rW64FV/1s/fyDlUExWYh9+G/9gsqT0lxjMUPg5Wcqn28Im6b221C60idAWvzDiIFStsiacAq+Mej
8F1xkttN7Hw3iqmOu4Y4EowAF18t+q1UPj+lnYGZVoi83Mqr4Yrv3KkSYfLkbhEdizI4AK8ElMHh
gSI1Hi2eObQ1BNO6SgMibC/elaj37kvuRRpsOF+xu0Cwt5ww2ReMIntzyydddS1FFgN17uXFOyJ0
+fiFE43Lc0j+8kfr9nEuOnsNVqEWF6ZSJRX+OvO0dr1Ry/OtWZy//yKrp3Pj1GSYcj1rjteR8nzV
wNimpBhgrkIqXiPQd2EUqLverUBRPBcgs1t01/NuBY4UYggMJCQH2rWBRpY9dqpwmfhRXxYPO/iO
3EdAis9s3Qa5711+pK3Jr07mHPG1qEpJsdRKZEhPgYJTUJ9YRS/K4bac/ktmlu3TXEZVhnXmFX6J
I2VodSUKlge1lk+zUNju48xIbEod3Y9p+YuXRLDkFURxv5ExsNNhXFGpMmUrw6bPem/04avBsD6/
DJM2ICsJKmxHAN+TsG63nuXT8rla9EKKV8QoC83JE7DhcX3ftUL6vkKowYFafu9jP/zZBgtTEPb3
C1ByXuaAk+Kz2g9JVNK9SNDLFCF7KXVBRrae+p3vLF4LjiMa5KLpcMIazdl/D9uSLV2mVH1kEtv3
1N6aaU8rbu3IbOjD24g3wtzQ6Tu6Nlp5KsX2QoxDVVayQG91chEpSqcLB71lGi4tVDMlv294xzpw
2q/J7PdDSCL742AsWvqqiPjcWxtAywoFzJNRR9sZAMYauxo5AJF4pR4aNo6TJ/PyZjs4h0PLKXSe
1pT3r2unl011jvp9cw0wtfEs0e//Pv5Y8QvWq6UUfPhj2K8pMGLsqpHJ5qqVfWGjmksdQED+kTou
3vvfGg7ZsXKVM0jmGt/gVPGaKwbp1KTRmbS/hpk48zYsJhao+UGs9GNaneBLPtLrAlq9FemSfCzl
gAREAF9QaOEFDI1K6wz4+LBHjlYDeQhjRRccY0O4j6U9z4Dqj5y9YzMycWzILaVDNNrVbBuWBVEM
mS8nOjwRg1k7Gt9gMkdr+Cm5iQtRD9l7wf5FJKkGIzZra5Ng7lW1rLtx8irW3YktULLOw1fE5K1l
aawazDUkTuXUSQNIX7MCi5kZ1QS1bfsC0p8wh8ZoSUKhd9EhDODiz2YTQ2+pX8D2N0MIJ8WY1EGF
tSRjilFJPYu7Q5s89nwaTiDSnSbLcNPnRZUUcgPTXFEl5jyHEkW8BJGy7+XCKSrjFKA1G/2SUMR/
1MT8/9hfOySGIeQoCHo7p+ItFUvpI2mqgj2iIbP3hjqTj6Ral5n2x7JFe92kDrscW0Z+Wj8wCb52
KXxJC8PhNOPcWAnGLz/Mo0EHQaDioTS4Pojabrnub8LLzMyv5VXsXW+2YjPOjeA7tMYZQd6NlXWf
sbIXNyJG/XJYjqch3glN736iH28mSmhcSINEzmS9A35ZI7PMyf3fPC5JzLzEeFN/vxkMhPCXM8KJ
VqTc3vP2cNUpvxKCuG+F70fCzdWuebtXtP4fItrxC92g5RhyvhOmWGilA8tv5jAaurdVeaNkt3r8
6iNtapudlXvRpGuMw3nNI5ihTvPt0ILCMd+YQkChFd0GopUy6pOUPE6JKp5Cr57Yx5PdAW5vzjON
7uRCGSleaBXMbEZth0HnJUsBFx/W66c4XmssqtbqSj8vYWMypdkNfrIByEiA7SU9BiXzYpxwL9XK
JCTWyIi6+8WOp8ezskBNnkiBuFFaAOHNwZ+jjkSxPt1tBPRjzuB7ZSgEia6hPDtu426DwEclNDWy
IKWYUp4QZb01e1P3pi+XJs9cefpD9eoJyjC0eCojK5M5VtdQGOjtNcmp6WhSj3CXtoIBwhhcHZSD
YwYaAjFtvWiKB1VCO3vJw6eRGaUX5WmK6bvtyDbhOatR7+V8HrBihpofi76Qdt2vnAaQd3DYwwec
8DXGL+7m+WwXvySMFwP6Xmc1gs0oL3V7gQPjcqYkI+31diODYYzKCbStMOdYjou0dhcyMmEQCXie
SNCGYtzY4HXCdt6NZM1PcjZMJzvL64SFHiyPN6fFgtn0g9CWdG+NVJCTc3qceVdw158y3MGC31TU
hhOsg1YJIZis1OjBhoAmrS+XL0FNayw7DA1g18v3tqIQcZGerDKQhwKL7eCBrxhc/Fcac4Qm/R5C
ewsVzomuD3Oe6yDvnFyrPcCnRqO2bIG/HEO+wlwQlSdx6HjoiOlPANVOpA52ebo1B6k2wo6cqMS4
PuQsfDJdjGdaKdVC1GTNNIWoBdZNirxiRn9EOixlxg/DMUjNFuaM7JxJLKGkWtCMLpbtMWvYZ8Lj
E7xfMzTugBOO8xQmXzN/Ib/GlNIu+iGGQOdFJX9jvySPKninmOYMQPXWsaapUbwnvv7HU1Tkx9cX
SDj1Pj20fasCuZr7v7dSoEqT5d3vPSCxK0OzgMYJ7RLS4oJSKuZzuQ/y7NET1H3wRyQNLjNyFfu1
7MEplkq97SEsmYpiieU/OMK3FfDEf1FF/PNWU7rPiZg9HeJee1nt19zNfX8N/napYSoYB5QbTHab
GK/VPfebtelIwhXyWfMrG91bJ+gHDLF8t63GDJRFP6XAygGYKklUs490Si+HSNr/WZjH1ARuAmfz
4Kn1H2OTQpXxBFXDUHn7wSeHAd8ky6z6hWf1bkfttJ5gdmoEZGFrDXxVAQ40zLesLzi/ScVmi4Ny
QaKpQmsyVcaL06acY3j7XPAK6PhI5muQQKhA9igrJU/0lPSafEUr+IZPCwk72fqTuj2sdyV2FFIb
keIrdOzOuZ7H/W00VC8rYea+1c4HdkzhUyKihCYkCpkU6KbAacqnyqMPUk5pKLevIQjslZJ+pl1Q
EivoRol3ZooqgjmAyfYqJzzT+teCgG6EBPpc62+XDbiJe+P8FuFeUhcIAfYGhLs4RGyA0jIjUosm
fanfe+KkzT/lwFYLvS/wFU5qcC1s18Npc/VSS2zGFtB2NYNWHL++YaMpi9SF7fINOXA5Zz6uLOin
eJIp/ZxhD8P0qDc6Uqwzk225jqBYi7AdAcrHcNWeoxJ0vYLhKzvGxoyC2TjbkiUds87wh7iZmgXk
7BuLLNwPcBkvGItgMy6PPzjpa6oego5gjIQl9WDnX0OmCc9pJPnRlPPGmu1VY56BpdAL7aQZmVTl
uzdgeat984oz9bVYwXYbDjL/NjSMzUZkyicA7SX9YAyWVwdXlKgEBuq1GLFqApwzZkBgZk1BSZE+
DmUHHjDvu848IceK41J5YXVm/2r1mzcCXkk+1OS0G4eBGW48wucR08MeGXXH1QOlgScqMbKU3TVF
uPaXzkoxa8U9pGHRk9dmmMQ8Ptqz4X6kKEYRmDA/Mshf52NNURdaEBSMOgjulJsmX7fWnNOPv80/
idwVHceCffmE76ol0E+sACea4qpKZg9NSLnv4JVwg1q2vpM6la1Edmug5vTkIZ3pettX1ny9O8P+
/N5J9qQs/RtEMzw34e3chMdvk4zT0Wge0Cyx8gmsiTq2uQzlGmZVuVXwBlss45VzVOjlCPYdbrVe
949TmNphChWBLsSN0+M+y02R/reC0K7d7TpQ1YI58x6lGptpYVsKEndl/Ppf+cYBrdadXf/JhpbU
0cr6dVsxQSmsKVW0PlJZkztkQMaf2ftTPmFepCBCx540TMyNLZfi6gTL7OjD0gcQ8HE985wCHd72
0OP4Tkbth2ZQcpxnwkgBfQV/wXrjFClmBp7mkInQMQ75xHVe1I8pC4EPsYCejedY3q5zX8gkpL9x
rHfkgkoDJ8H0bn8mXJIyFK76/qfgSqMr9Hovmge4K3f3V+kgC83dMd/wc/jebugp5VtnkAmPpCXC
YUWIKes2OYip+pEdyIDTEsa/tcioYEbM4LhJsZ7SR+HGIq15YxVSV0mPsPeLx9+0NAiN9sfZHdZj
vvV+BQS0CVTR+Eb7jIG3BR7HEs40EqWY8EPK9iCo7sftNS8p81+83hrAmCeAE4X65+++Bid2yjEE
fv3I+Tx/d543ESczh8GfGcLn9zGOm9BJIZlOmvsZO4usr8kEOS0iEhQow7Jp8g24TCWbEnzKXFf7
IVOnWGT/X6AASWJGzaKiVdbO9rzmwwdNMClRD/DPrVn2S3F0Ih3JefLPz5UKf8s74fCjwKh1+XV1
xYm8I+gGsL9cfzrmNwYVZ2f/Vqf/KXgnM3ZjraFWRqRTyxKyOx237H3VkZjCCt479L87ya96I7aT
2nttXR9AHh1xE2jyxPrHbrL3HwIvpJ1xyBCYyBa17iBSCgSTqE/8/pLDEhNYeVJTHIzFBlv9/V4d
3ojLaQXq1CMFR4YPgLO/+24ofea66Sz/wAZHB3MsVyHKFJFtt15OjWDsHNlovmeaXuo1nAysaN6b
FaQoOGXPfBAyfeFzZtgfOZHMWxGEyIe+yaKUdbMxWSB+PvRrwg43sbGovKgDBs2gvo8KTvQs7Mdy
rO0Wwu05ZTLPQ8toKqC7aDJtteTFkFqwbYV+9tcXmfePPME3OnWyeZaEV0iJrgqk5fCboyed8KDW
gIxUumw7goJ92voFGc7LWwKTI2PPURr+9KUkuus4UaNp11B+VmMGp7uuNpSrM0LQOepOBs2L70tn
1tkeX+MENT+wKdpoMbWBhAtGFQspxa+CjB/VqYlAnGHuJ5x38WNZFnsYY3Ihbtvgi/vaGobaYa18
T+FIFICuMmawl15AKtdhtT/I49NZgxE2Ug3LO9e/Yh9VLlI0+pKOZCqRLSicSgh2RqnIw6HOwQtt
OhSdqbi89h/qgh2JIK+mGAdeTxxq+UKppRPYtN/0DGK4BbPjGf+KkmOwodEDv/+5q2lJQNQEJ+If
tHVs3DInaVm87OZGT8khukYJfMjp6Vz53ysq75vo7zS1axPe7MbvlflYkXR2keA0o3Cz4FFHAYyW
4iJdfsDyZGX4wLAHQuEzV0pcSE5YROZrzTBKZBtyxoZtepRAyF2AJ142clIKOO9SGhRCrHRgKmLx
KP2BZh3NNbV9nxnJGEXPr2+33a486GKhB24v05XM6ganzK/3ReH6Ynt0XY9mOyFd4eJxxnIRl+d9
odjv43yzqp4tKrE9mpZTlgTjnJVlMYl/2++BiAH0Z47UKrWRsxZ2t9O4cdzqAN3oEWl9nDYX0ylb
h0R6Gr/Bw2U4VYLnpZzAEWrVMmy1Qsn6fg+COMdt8Rd8pAA3awLDgUyAO85trM6V7V21Yw+vp+6v
oz9xmgkBHG4GhJ+CQEeRHaulNOgCll2yEXQC9tLcdCX0DVcay71WeEZ49+axQYYY/wjgYuSvAz+5
nk6FKfiawUqM2vKuYo1gOp0ooNcbMymy+QBWnbzXtSPrOw1i465UH+/DWrD7goMYeHq2b+0S65P2
OVezeBOZ76MAGOhRwcolfpBxumo4kYEFvkxpZ+AusERTLbsruZr6EZ6LejJhdmtbXZmlQ6/8gnVr
y4BMvOIRNjRNS2Wr9YSFMjSIcq103cdOgaKyVUsyI0Pdk7WhYxZcI+jHkHE1PIhwGiepVvfZUeK0
fW5Blzq+DomUsUdv6PkIPydbDx7vxuRmpNPXqwJH1rAB4janesHnidoYcKk+z0yHAAMqsTurSo39
NJHD63ozfVON+faYff0I0rsm4yaTxrxGgsuFdxM5hkU9AI9KKPrlQjvfzHygFmWMom05grYi7IfV
cHXtdcN3fQ0pEg9sQQDSd4JB/V+X9JjQ4FqmbhP4u/vTvCZsSxXgEXtCNAeGZkOLZLVwOaFlm7dU
++n4tJoe+ntB7yPkL8N4rtsR/aZoQqg6i/4aT+Lo2CUpQChKkfDLVJo2qEnXAW28ajk/V8E7pSKO
xDS6e7MlySJrRmjcDMt/j9AIUkkY0PWyNds/Dt/pZDe7LhyaNFHcAxLK0yCLcuJpTsftKo38lcxl
QNM0CXW3FXOa8vgAmPTlJeW599LtOU116q4nRWq3buwwy3M5CV0c0cWD4Mjxp1w7ilylpc4CBpq/
1p5Rmb5mCKUH09blTb3eUo3YHvULMzmalv61dNk+hhz5uvDDC+IY11y+leAAuVmMWhiieHEDjHeX
9BYNsQBj3ibsL54mkNlxSbjxhRs8/ApuEc77f6PQTzlTEouhm/0IMoDV5TeHffihWyj/7VGwD3Fg
yzmgA/+MwiE9bDAfLXoVI+ZF+o0JDohrv7qXAi4C24JlwqniAINpNm7p0nxxlSlZvn+zD9AG7oAe
NB2m3pRvkqmNxda6/vslcXVT1b1J31Mt8N/meOGJGz3KP/RJl7H8Z6ronNVVxcy15KqfASLBb0Ps
NXrvxA2WN0D4dI/O7WGg5woq+pVrPVeITkEIYUNeJ7m3lzf18utAs0A8cbpK8tOsUPySTcqsnVlC
MWvdE26L5FgnzQ0shE2F21C71YsETEXy9+6eMFefXIiztc7i/iX3caoPn8Yq1D1PvkuslOkAYPra
3QhBw924OWG9R5GvCmAXql8lnzQ3V26QjOFrN6O+hTm7iI7WpIAfXL2TvD3N9SAEzj57glU3wEqI
iDQDnVCEbN+25jpfX3RAW0k/JhmTqlvIfSEeisdjQu1LJ29C19MNUqPKNqwX/gFxlye6Tl1u+V31
gk1O72PO4A5wqo2aOaWUpgMEPtOw8XUdvmDVhv7sWtxmkjnCjZcxbgfN/thN7bt892/8qqIRz6A4
X+7BxHqgvJx10JCszVLc19vq9qqYaOJkYU+UQAPKf+/+U6cKs6iI+97aYJGA7bbLBXRSKDgsrAJz
Q3dckGDHd6DH1EnwDQeL02cMqH4qthp2g6D31OcFek4jP/znIdccEt5pVrYVx1r1z+IqXEY449FJ
aFKQ4AiUk+kS4fGxEzGesA14RR/3gr7+1cX2K+m+RyQ9oI7EsX94We68+Rxhr93WkTrsZpUCZFYp
3W5Xz5j4+JLj94xgNqEjSam3sxk6ON9bTlxAepLcrCmdhDPyPSouuQAIYg50+9iRNkgClEWbDn32
BSD88jaEVtDLSduAcg0qv7E/hj8zpj837rpAnNYfK9JvYqcMT4RfffdEYr2vi3/QGD6eDK6R6/Up
yBuQReDyo0oJhwujlJ9LE89QSmarlrWaFxdQrOxZFKQlNSL/3ZrJkgop1qlYtGPnq+y7W+c6R5yV
JQlTdABgUUGGs+9V7SHn4Y+tSBIQSjqwlcEHjYPIjrhVUjAwXls6k60xuGjUjMtAiVgYd48Iewo4
7lsDxPV9SJupUfkCtt4FkcR5ehwg+8q1qeLB5IGIrLzXvIO29ZyjTYVm8K62RBeo0m0ANzJwplS+
56vBrmUwUdUosUbXgV0ZTSNbawIYbZE2S8TF/piB/SxJPXDttYbxi0rfaq8iJNSSywP+Vjdn4Ppj
uKWhumcdzfF+gHdBXOtUub0teQiOX+htm2mX3diE+V1RM2vIvKcJKPeAfLvy83Fepr8zw2sUsYO4
0eWpqChScvjrNznc7Rnakq0h/rd8LYCvMNHY3uR4W5M2ON1gk2g+FpoAhzJoC28V66XydvDPSqFs
5XG8xfs9pBvmrtsqsWflEGGtEC9G6Yp/UKgyph/5dzPUMx2gMsHK2FAmA0Lzs7Qsm6NupeU5jcGV
BOoltM67Z/VKVEC6icO+S6ZbhWFDxnID/CS9m0XPsvLyzw82zB4H+kzM6aCW7e6cuZH0iPUTohEV
pV0NT8Ew2RMDLOrfwwwpBEmlzoQYuN3PGWBGtrJYvEfKlAy7v0JawceJuE3747IpgrXMok9MkbjD
fPR+4e2/KwxBmTo86XvmKth6b9eBMjEZEhWzzbJeuohrDeAmSfP0oscNXssH8k+0fq6I6NyVf9pW
zcnNI1RTwxxXWMg8yfZzu95OMNySME2vDT3vPnJCTm/vh9PelkFNTDUMLWS2IyDVAvBYioVDTA/g
/uza3AM6ZGlRJDc4UXri0vJGnsdRtFs//kjWogXyqumCvg3eNvnoZnrEqIXBSEIVjD+/zaUjlov4
Q2J8kCtboTSC5VvfVz4iMdtTVSXXED48gSJwEocnfglAZo6SKbsp1KnFRehWRuPniXq1Xr9Hl8Pd
3ZL7dcEDgezSBsnW2iz/BbIqB+IpqqoXzcKx9blT1uu75NY+ijz6poua3b0B5YHOKLg6IdlDoMZx
53RglSIPyVJqNeeTv7AizojhrhtmD0/GwrVu8bXh7/UA6u7Y5R/WUC2JkcD5JFxXO9POGeYH/P4b
58BXMMgxu7ErsO49DMiFmx6mNQfQZd+esnk3lU6RIQ783AouiYKQKkd9c249SRdb+HJcgkoGvzom
PEY6ScRMiKjXPK9DaZDv1VQJGJVeTUNrDDkY5g9oY9+/3ORM4sbHLGjjWTAgKNVIlqiu7YK10USm
FvPvtbMSogQblHGMYe6jbXMdKxxAES5K/N0ZSB8WXeHqJU+v3UgvpMgV03VTjM/wYAk/Zhrhdv1G
d2dJ3A/E2vxiGDGPX5/88QMI7k2Uk92AG2r2wMaqnSk+zIqIdbziuJs/bQWN95qAvPj82kqDvwMe
Z6IXIqZJ5cCnVA6HomSXx+F7K64weCr67vWQOUv12oK7di5KS0RoyCJhGBCQanGQBB7M/siz0i1o
7gHK36ZXjITkSxU1bUaYh7BDAjLobv5vQLQCRTMkkoYW7Ojpe5yEtt8DuR5Dxvu56E2fxi8PNXQ/
vGzj3Oq6pxzjjrtS43P8BglJXNfcOoVw8AiXTmRozSqAVQ6K7Bim5jzdIO3BiX9o8Ab4UrrLcwd8
HFx5UzxjFMYdl9AQw6qiSQX4TjjIW9r9N7OQZDta2nP8ObcOi2+H+6HX+oHZogHbrNIGkBXDFQlQ
XuDLP6AId8Gjs5wPYuNoizQhKL0yhoeywbBRAGwf0GaCHYEjXqz6dAfqNsq79iC6uee47bDlM1+e
gwBwXQThQW5TqbNoli5RsiUsxwJUS95JnyeMno4KmhJ5aKm6gp2dPd67Tb8Klk9JLx8iMlR5xetK
gvmHOvNHFt0pZQHJtq4hIelWqMAfxokIs8oRPnJ83+hW0G0tXQAa+zlJlBNPoJPjQkljXiht3oA9
D3JoSJgrNvI9VH0uf+M3wKRYI8Obvi7XW6upWVpO3mAdM4a3wFqRc3KPz0Yke3PQi2XZ9PuHKbiu
DU6miNqMI9rB7CEc+NL9t4qDc4WCvjx+zQcWJLdyIwtbtEaV3yFA3myNc18hV24YApglX6ZBGbNS
gZiAEa+iC0C8kERidZzHAk7p8+usW1RiWZYPlyN9SfDdGD3WEhqohFo16IH3tM4++lUOc+CC6B9A
kLHFTEvaUQZ8GxBj2tp7JJpxj/tDFCtUjB7/gIXgtZnBFnldAOAoueiuBYB0kRszrGm/Z0bLCq8C
7NrFmjVQTcT99qyOtCgoqYqxu4UafJJNMQUpvoj9p36Wm9dkLaI6AE1wpn73hwcpUCpz0GaNjKvP
Q7KPtpvlP79u0V4WXRzNl0YY9ScfnAzgcxHyd4UdkFx9LPf3T5tdSYIDvE3H+gtrN60QZCIFsZzj
jhetBNnFIkkqx07/AAqXp8EVvWGejN8Eu+mMHs0NJ32wjlqf2lkqUAU4yFZyPStSHuy1Y88bfE7T
HLQ2Hpuzn4UkdNnwQFncoFsvGO9PkJVXIUjmv/ccAYY5nVn+bKMESjRN0tO8Ir1dnXrj15BgmIkf
WRN/zBHRjuNrNcprrknppUJ4vPdjGy8EWC4njJ7PAQBxEm7oMWzgYTl+ZN/tUWq6TgtWEZBAbiTs
Bhmh1MzjeRqyZHIn+6lTiQ9QIw1OueAhhMoMezNa8tySxs27q6CLf7u6fUORdG4Opkcszj1DneFI
8IikjdLfqkYesfovZdCn0jjAP41LmODXGOF2a+TbaP3KYb+tzZBxSlr5VUq8r/EHzY7bqAJnNTiY
8y3e+iy67EMOA80osfPtvuNh8vbkbxn7VEr4Yaspmur6nJJAIZ9w3492l2uyDZFmevH8KMc9pjcP
ozC4CojxEFghdOA5N8TnZ5dqMQr0Ows1v5mN6a+Uw8Uv0AQb05aMbxoIGleb95ilCEOLgZzuSLBP
5SCnAGqghw2dSgmfcm6gRdSxM2EHVp04cwkv56DzTcVDD4PI+4HNyAubZpBhS4bCzCHGWXxIZJJd
S9d17AQEuvKFNO0uMb709Ii7+5h9Ba7+WL0/FIZk96yzKSR/ijwJ8H5WEhWkHClMMZ/D5oUvyZr6
YePX4tmwarWj8VoSdvugjGTaA7yB39cvvUovNtEPiGUdbvDMMvlN2dX70EB8pGKhZ5Wna16qi8Wp
J/C8GHqt+HpID+zMPnKNFo5XcFws+rqNqD4eL3DPvXBnD9NLtep+K9fH38SurA1ZTl13Q3n2hOzK
BmxNnI/GeSKipU8xJqeSxFV9o0TbReClc0/LoLUU71vhGy+gdeu30tuf8J9S9eSfWJIRHp/iGJd4
MvN2VKr9BD407patMfTuEGQlFxy8vJHqSADCANie2L5A//vL2G+kHxXMFHIgz3r4X3fMB3Lncv88
Vswj+X/f57Yjhy91i9/X0OqhizlCf3YrzYUgvQiVzollycLB1Eq/bN+I9gXvKA+rZyFAQVXrNVUy
HD3uF8xOwZNZXgnCwS+TTRDBHT9oBCigzuPoCR80tLUlXxTp8D+CEYX6CTmxI27mnd4VKQ4vUrdI
jYHSkuPZaVRnsnp0XC4OaFXVYiq8D27AJ9D7EYQ49sEXcOE//IQ5a5haFl53UWi8HYlOLTwvaUcr
v59HcPCkyK74lRrnzAvzcChAEw2ygWbugJzdvAp7QCQAGPHZElcoqdZhL96jWZ1zOI9lThXMfAUG
+4tcHZ4IjZJTPTqxP2i6Yp2gqC7Oipw7JnGmQ77Fv1stJg9IVX+maYmH2gnDcPna5dihZiyY6zSr
OeLa+HOHXj51JYhJ2U4u+aPn5fa535Gr4+2sSMVWDFhoOkwFDdHFkWpUeWCY0Y/7zlbbpUGM8ZRZ
OCpeUnCUOKIoAbMiPhHFd3qRkOYGfKMzH/kPbkNpMGaUMzcbxTeZqO0syTb9ji+80UL3rndRvoUM
KAjHPCiy1LjGI6314LJVWB8AGsVWlW37rBHZ2qUbHgt4Z8M1c6KRysOj7uLSPFhrHlUAdnNMiMR4
42YZF4QKzgGLo5Piz00dKhGy4IiB301WEn4vFpMTNcB51s8Qq8S19Hq2PzcMAqUSMHMbOnDALZoe
O9f1aZ18Zntc3qzfKlYseZ02BBZhhWCB+hZqJ3YasBrwES1pXw5jl0DITfyjT8x0EGSV5BjHCwWK
cOpIB296h5fipiXe6ZWyD2nhlnJ4EJp8/Rk0GRf6Z758Ls+NfDOSG1DOV2XqSQu6PGhUOhkbMX0S
1NVmTCCYDsxlsdryZh2ExKwJCzl9WP4IcuI5mtZBiJfXhMBhvG/vIf3M8T9xFrenq50oWMnpmnr7
Lu0yEsN6VQXKzcWTSFxyrfWDap4eBAFhOeySUqGQ+KurRpAskJB5g9qIgVr4gnN8oTM8WYBakM4K
X7YMR2tslgaraK6gSJNQ3kYiAANBGE85MmO8v4kmK/CMjY4/U5LUKwuoULx59LMfcOB0Djln4RMV
TnGZ31ABtCnjmiTMTrtBAMgpxD8uruKUkRnswWuchPsurngQUJOC8g1P3yjy8XNi5JuRUmk3brEd
C1SU+1AEAtII8D2bg+EciqgRdBq1TL5DNc4c1ErkjJ28pokeOzWuuuu1Mhv3SN6sJztZGBj0JW49
J3WPUiMbvNAHeTm19+/2mWKKa6Sjl3o7nMh8//a0qYyKB/HBsBhxn/k5VLBUNbrWEjwgXKDcGRst
whWbW/win1UZcyzO7uy9FzvaDLaMWY3ILID5a6dBVwY78QfcaOWHaZyeBgSsRQfdsVSYCy2U7vSW
Mj9XR77adN5x76ZAErtR/tVAzTXmNCrSjmo8wg0GEI7JiicMKR1M4R+EFTw2kat2938Au6u2EHJz
6YoLyApc6ceVwJT0NlB8N3V5jUeiVWEwsm82hhzPyUsx6laOx8e8ZXHr20nK3ngXYKAJcGfCOrLe
JSezMyIG2LbfEhIW1IzzbO/cmEbUX9VF2P90F098IB0gfwnQ4/FghSx/EBJHLDg8Hj7u4iH7D8PD
HP/N8RlITkMT5KFnwcMx3OLgJxaBDpW75JdWo97MyLa4f/AchFh8NAPRo6lzYH+r42BXFcgdd1FS
TWlo8GZAScYVX7p84QmCBs7ocNS5kKQFM5wRdNRzMPmOcGwcVp5+oHbt1fukWsrI0iWVCZ7xH673
LqpLexbQtbuabRnNRPTQzT5AAI+Ox3czmIqDHoi0rTFCAdBNlEVIPFRy62+gDJaVoqBFnO81oBfH
SEfTcXkUj0dj+IxOvmfHj49vgOcyl+bkOjY9KF4Pd1o0jK87lPD5uTiOaH2Fmd056IRz/mVx3Roj
JI3xp/YJ89EwB068b2ms15moGVYjh14vS94ZQfBJtcBQrgXblvOEKVFno2Ba0w27x2hCHocWpjZ6
6xzXRuALtcS/e6TQN6yI6nSftWJhyz7JvZd8zYJdQmbts+Vpl6GXDd5LMTCCd1tBxFvzJm85DRA0
eDSSVHA/sD7adbOZuTz/AF/XzoWdlvqj/lJk2IBkS3AjIcyrehfz/RQ071iP1kJXqXjFE6Go5R85
amgSrY6HXJNdZJ2CzHmJvD/MbqWqkaFvPk5LJO6FWbcpjOd1P5vsUCUqvdsT4g2RiRBVYdfQJEkG
f6OE0UsyF8Db9mfzO62BYKswbZaCl+wAecIYYuyOZAVsLlTNNqUxwqx6bfEEasqliMdEpdNFH3hs
KlxT2T5wwVQ+omz7SeS8jnTpce04hqEyOLNAJ0ANa93vVXs5X4y9u7MoFU24mUTPOzjdFdbQRHnk
Uijm1+KFaP5h+Bp+TczDbmvxkPNPEbGo14geXNG3Gtsa1x2pQh8AX9N77uWw+EEShN6/MUv/Vapy
0CCczXEX9T6jzrOxHxA6t78nXwY2HsLSq0e0aaXQf1tR29C2yM5aQCV4spOOaPXCvoDCurRKyfhJ
N+tCUo8XJFZylPWFlWAAlFXdhI6rpbNzQkXb7OsVj/UIVeNyWG37cAjzDHUr2C2ROQ6qptlE6MJ2
FC1Om0YVxW7zWLgpUw3NA4wj50SoUD+6hIWIUx2G88V3jLZ4t7I9Fah64dxLkbfW/X2QZtLFzOeg
ACJOOxLif8I6aFlLWc0BBO5tbvE3Z3jw7a67lE4sEhBANnri78+8EE0z1thdGWgsKRHAKzKGcPf6
YPMQnErpYhhdmh6MdYDV9RECiUVzOiBQ7YRWTHrxIrluppIP7a3YZ6GiLtVoz8RHj4dXHscxLukM
aEBeQyFRLL4LfeDNHdt1g3l6iM7bPKh9qobZu3Qi44oN/q/rDfCbi4JMhAk1WCojm7MJQ9k043bi
nBL4vFzFMOA8L5VwdqQqH24aST61jHBQ8Oo9PNNVnF7XoHAFTwAHZU9WXQ0SLALFKZVjAPx3b7IK
H+Cp6W3VfnPoNUYcxcVMuJu3t7WKvCGCI7mblJ7LBYK5shcMUIqfyaNzbNDaJ3dS2H43ldR2AyGA
dQHPI58BwnsHifI+Ry4HDEHncy4xhAtDXrUMsAW9vW29cbS684SE+mu09hNGEuZf7UEMjm5MCeaW
f1zs0SRAOaDanJIMQSuVCSA60WT7bOqgW5zJo5hq8avwFpM4+Af30EWN7zjNMUCd9Op8UlTtu+ZL
tObV0pY+hF2fXwjr9qeYe9Itlrsi3CLY/yah4K2VR395cykABg7o39yvXYNL601vBCVTXXjIuK8G
1p1S6wlTVeAJx5uIajdi1cuRRsFVTWMnQ0gBaLNExfeoBB5ArbBTHja7JK1CQiuDJJYQcKFYWCOZ
3HYKSJWUu0D41ejZ6qVK5kGo1E7YPOomBghm+wcbDkLCyVl2RSnzMt05W97ovuigvhMd1szxi4KP
mOHqJHWgvHvivDqLgC/ncm4nDQpHU/OsrVg5/h22cBql8ZJBfOvEXFE06xqMW9JWInvZKMP34Xk4
ZG2pKylnPn/0d05uhSTULRHqSw8mRA/7KwndJCeL0iypZLjdhkup6B5Aa1SgxHwiZclhh7sY9zoz
/cz0vp4Elncl4gHJdUnQMX5uvCpMvXrtiFMobWXdrGaZp0CJMVkvYB3w9uvI5mF0WPXLRdzZf3qI
9deI1iXmoIah8FF+ynlMiJkTjOmuellhHI7heQ+Adpx48fPCy4CJ2E+PAr0l4rQG4pCGf4Or2QOx
LHIeLo+djcdaRC54I5M4TvGVzeI18CX8+R6h7/Jul7T0SqHSCvf6sfZJKUqX1HN2nXOkRlr9L2n+
8ZhkD/eRVx3F2vMgYwbiIdAhTZCbjDa++Y2oV3SDqSn9fLrGoFO/Xu1VB06MVdSW4B8bOlly4n+P
/3plK5oJPZNB6VJOhtYjg9f2+LPdTTS4EU+8XJmhGby8VTZwwy9ygH7YvAfAj6jlQE9hkmC0qnto
/3p+yKLH9rvnp4NqszJW5Fgt7jJ4IgvzMb0EK2ziqrKSdJx4fqS7RjXIzaoKFq8ifgWouTgQK8R7
HtCoDWOmLk5I1RpcAriMN04AnvygS//43r3IOpc+vX6yJhZGfzkdM0Sytv6p5GaerOl3sU/dzlCW
ypzlfoNfBa9TYoA26YDIUqxeRaEoVY2SV9CaLDMApEaPexTGLZbhtlMzbGg64Ymb3/4HD6hgFvhh
lP5H3BsiRYSUpBQR0RFVbRjMY4m/PKCQXxcx5/2AVomkRHqGce0TadLXJOvhyrpP6T9hPtCKH6Yz
hCmvHiUJF7X2e3PDpgXSad3EQNCu3WW80BbgCDZ81rTk43U6vSItxf5k2Wba+Nlg8seUX9nEFZc/
m8adCpYmsVq7zO9VuafgQHtHry6jp7g9/NTUHZpebg4KuzPhZ39Yu54YYV0uBHYk1Q4D4hYskx+A
EaYVzBv0WWJrDHnj/IOspdO9bVH3ORO/jIJ0CCqpWmRmt37XDYGGGKXGI6cgP3ulojrU42dmDzti
e9n2Q8/ElcoiOL2evWPDHLJegDHI9IWj8jv0azd1fuMZLGTwGitMiPrheEi0IGscFHQw+47MXPVp
rBvdd4z34LRvrZNwpNY017+HkDvcvUHqPzlKZRbMUXLnx8z8GZ9kEVwoPBru8j4glLLrHPlUuEaO
7+kgYqGSELXxVEJL0h0KL1kV99zkiQRWLMr1CF6eamU0fm2fOnvS/fhkLsYN0vPpcNHP3DgYlFDV
m5ZAObPeNIKHUYkbEXk9BJ15s6QszHiilgI399BaLuTSwx5UHn89HCXBrORpuIV+rTKrotWOzlun
cvqSSEoXuAGPwJqMu7vj9sba6Oa+qSBPaXWGNhnAffg6HA5NtAc6gb8FKmjIBxQiiCBBj5x4xAgD
Eh3FJ13G/i3ysp5+gplhk+qWzgtkvKxqyrWhMfeXukWFAFoSVD4Gn5oYBLe8ps+HuLi/rF/7cRLj
dmPUPLL8zMp+CkdtTYaC4NI6OBPOO7AbQMdM5Ty1D8mUU70Ue5bNRk8tsMFqWt26lBXTA+kG5kn5
cY1c/1CQYR0ybDJaG1vv3hy34jJ7GYpDqte0VxT8zGxpqVbOOndg+dGtXKUpabSHSYNkQWCEpN1g
KPQXmTXs2X2F5RjidhWfo5g5vj7uvfr9uTqnw4M9BoNiqkI5Rhn0w+P3eVYiJ5/Bl7G0bNLE9k8B
jDuFcNmVyEt3aOckgdBl3IU9PFKq9bXYVtesD68/V3O1lNcb77CzCe9tmGPZWf5X55CONoy1hJOY
grSk/srGLKCX9PMB3oaAbvrcVvbe7RZSbju+xoWSUyydTlpcBHR/KiV/p11qq3tUZJpeRrFV5af2
IYljL0/YQrYFvzclAmYOI+XF8r7Z93R3NUgRWqBq601dkQuDnzgkQxiodaA+XzBlXSW/7q/w/qev
vSbrL8fj0IWSw++IpQjEtMlctek0Wnnk15gGQNk8UXAKv9yAJTOfsGMtFTn3xmXApdhCTJxq4I7U
oXIjXv78X0lp33Mj5C9RGTQR1IFZoknQIwzNeAxqhO19qRffDOTZHvYrHb2ZS2VD6ZadL9oQsAgQ
VSSZuC1aB0g2+zH68JA2HhNg+XPFQuzHczP/rf+44lpMC5xmiIFKPjlnBuXIIi7Rm5zLI7SEie1x
qOc6b0wJ1rUPVXVPAvEhDFVvU/eZdk+luZRmG3tndNFnM47DL6vySsoVJPtC1jxyt5gMBmB3Uj86
PgFPEcDukIJmglD9sdgBkZbFz4k+TLAtYVoQv6f73H+HfrK+PprVRR4y8qJozb536WWFNX/tPADX
H+OPyhsS2Cwf8ab7tOXhhSniUh+qDVtHhXe3zXGDC90txHuLYNCfVQTVPLLvVsNcXVNCzU4F8uE7
LWRFREbfBTEFx03xIg+DgYVWJgOmb+rKBnQg5WkYdnlQOeHiBMtFWdNYUq+WzkeIa3YpKDrtHgIG
B0Q1XVY6nZ/szvqI6Wd1P+QfhcIQAAedFdwxlysYyiEnfL9uT9w9hlOgNOHqzQf9QA4VBKU6SLAa
rj6AK7vPuPqqCKNyokNC58KwIgSI91CIl/CPtUkbIh1kQ36jv0J8kC6RIM8SjnJKTSFZ0ocLe/JL
uIP8dzN1E1y16A4Whx4QxuNLvy5vzlgToraCr/MpGHu1BcvBf5HSFdtm9MRJ3ZvOKylt51sZdoYx
Tyi6KWZ9dFA+gKQUIqoPVOV4MWfW9o1ilIUxZsr9qTYn8DEP3N3qmEf/PjyOBU3IAmb0iYgAkcZ5
iPrRyVRD/P95XVcxi+WMRWn7O5QrFuPJ877Uj1cOY2WfPHa5+PEaVWyt8HU4Hi520uLNQoqvtPZw
J1VxZTLhVrY7s3TvXhOK5/l7+Ke3f6lTWDLre+h6rMgoQSaBe9u3qMixKu0glxMtdBguzpqGojh8
QUnn6TBRuiQSEPEKAd5lHt37O2LwZvk7qCMl9miNgmKei2x50auyE9WwGZHrK4g07vF6+LagtG4D
IpkSBN8Ul9QpoL7N0DCLAjsHkFSu17K4izVjxxIHjkFLglU8xeqpBJTQwDceXPakDAbXXWzE23qr
lvvFdj3H7ttqa6h6tOSif1j1K1fq1o3WL9b5svL4jUp6/hm4dfiwv0Sv/OEfUa6CPB8J5ulcFzSe
vhZ4yMo8jLECKImGz87mm4i4lsPaigzqqIzr9WdwT1lwUWf8G3kRIkWX/N2DqYmuif5xX1itGxSI
3U5iNONYEYcqriPKRPWeQsTPKYxpMlx3G2LffdSQBGnx/CG2pVQ6im3RgjqcT9EWFEDFswARDMaG
+Z62r28CHkfEqtfhzDT5NgNrv3Sw1DmPVp7Qcag3nRRkgQJ6PZyDdMC7FDmJOA9vH14ilxD/PDWY
D9y38qb2RoLd3DxNmVUNBrsYuzSa4PBvuZowZmJcQ6Js20J+pgkn/W8QDraX+uIhHCZCvoixngeI
hpjIEXbdbHyBQMWcmtxJ4B5IZHQA2DC4DwiAjR0975DEFWeJ542ULjUQGMj81tg/IEr9AYkZzRxj
rynbWdIEGxCD8IsfrBaQ41uUO2DPkm3jmMHeXl8DAx5mYprmp/M37cj8tEOy0axtWOVw/pYHCwFh
7fwuF+bgyhWev/7zqKoViDusl1ivcdGiR4pSxhd/v1O9iqeMISZ/Ae73dBOmKlbbkO5Ib98bqiUA
1fqAmjbqhW0OFiVoJV1exHjYsI0xFXZZf5I8VlTbHYLZXBTmQunPJAoRjyJQ9/e8L4Ser9K5pL/l
r4Y3a1GORTe7L5JoxlmPyXD66zJhQVmM4pVhM99xC60Z0yoGcRljSzWdQLl5OtagensSUiDw+JQJ
qZEYR42MNE7VSwH0fKtrhnT3qf+Trjf3ft5rnwAWj8it0CGqj4KUGkNK3J3gmNXbANMi9+2l2YT7
6B5KcNG8TecEvEG6O0RIRdrKb+zpEcDDPDRv7H0M5eaz8MiyGlUe6Rd+Uo+xPfJhLLpxe5NqQQ/w
jRkHLe3yMTrsq8bHcxibb4/Z4BSZAvu+55EDfcIppsb293jVRejimOFbkWZAijC9OaJzf3y2HhRa
En63JWT+guqaId6YsjHllTPzeD/2NDF/mrpJ9wr191L1wlchs9bIt/S5i4oh1sOrMIBmSroHhNh1
1U8le4jnHModzlx4u+/6YeZnuCOQNLGUPFlURVXAQGOkW4xU2dtx38mEWFYlWqb5RSeNjLeJ+OFd
TlEs7hXOT7AHiTXAGD3NU8m9zvZd9aGbdvs9FsSTmAypwne6kCR7tpMuDfNHFhEFqs4PXxMLvcKD
jI/PVwPAxLRTbS0DoUscgoyaS3ZS2wtyAic2HiepDdYHuJ9YVFhm+NDIEhCZE8JqnI6/2hnQlCg/
tp8jn9iqLbDaC/+yCQnXNqgNFd/nETl0I+PlhMV7tQ5nXCVKU506MgHj7TeQN2VpTntct1t9MzTT
AM00FdM2i2Br+R/BEnffFi7OWHTSu8RDTqste93VCzzQsGJmeqWYv7DLbd2Fv+UxtKTkWqIEyz/p
/d64e1ZXgN3RLYykojANLs209UybHcRTz9fTbu4qLgvv1Iyh2LbLfVaSiu4zWt/ZWBO6llA4mQMp
8HRWWJg9bI7H31hAE/SpZAn5QgSLO2+IKZ6pFB1HyTPADtJCNsiHK0saOGB1eOQpI7nehyzbD1Me
IonQPY7w37calsRByhzPHpMWPQYOZKoDPqOLFqkO6ewrtah8AgLWeCxWZTHy2P6kV5Lng5uEnvog
T1p9FYHpfm2lH2T6ElRqGv0GH8YUOFanaaAyrmRHTmI0CzrgsO2S45bA0U417ZWWCR179kaecded
IZCc7PST09i8jDU3ggh1vIVyifP0bdfQPolNersHAyXvBaS5zmjiIKezxOoto3WUSwhv53fHhWVB
ltDdpUNdC6kbDzDwo5uJTersUb+HIKZSeif5Z31pedScvzcV2rf877VS+zaLJpB63EYmK48Ngksp
3EBERwU0SxPrv66DIgmT6g7oJwBy1hsHg5DfXowUEhUnxrKxPHm+9Yuvi/hEA/8v0Zel0WVQ3CAk
JCzrbN5+lIuCeO0dDewk0F9kcEzXpMl6vUev+2jtYXqdyqY4YZyYNyRziygIMe756gCcfpaRR6r8
PEDHSvQu4kjzIizy7sfmVekXd9HfTUGWCu2r28Qn7MRlQj5eqgb4xfMlrlbnLi2VM/Ya0tsFZp1t
ZGcrgaDdb7yHwTKzHivkkgakFWMJZkQtdJk7szrD2t8VgZ6gJSQMOLyshJeVfUGsYmuons5qMx7B
k2x2aE/y69R5qV2YBO8OdNEbvGM1EKD+yhc1U9RdlxkDypYyANCXb0AX9pAhtfr/gMa446m0Reth
H9DZDFI+5dadRn8I6JmQj4ruFI/93tAo5RJS5j+Jp3wIFMKDZR/Il7gv9JVx3kqAJJ97OLl93Ux0
fJgudlUHl0oBxUQLicTrK0QdSZpnLw/o/SjKeOQ8pBn6w4h2aWFHco+GS0QjpKnDYd66WqkVgEtw
mSMavZolrNFS0YjKQ8HkZfgTG4wzB7Tuck2yA+BAs6PYiHM+eoxb+YyJ7vVyLMwLciq/s8X9wYx2
Kz7RjUKUFkmELyuEpli52EiyXo5pIv6xn80qF4zsyJCHh8dGfUPqtbMpSmzJdNNr/Go5bHzeKoHC
UiQvQsK7+eHrhSnR4BqPdYf04C1vDfkhCmb0HVJp2wDaSw/Un04gtFWKftE21fPl9YyEB42al4NS
Aqc0e1JyNEPIBdQVMko4ydqjpNbxmyHX/068fW/grmp7oiAHt+1oFkWWMcd9iGQgL0R5HPqo6xEJ
G/d2tzHE5fb+KFREXlhtip6gNGD9z6uQUNzK8IZujnqZkc8r6e7xmaCv1yth+lzkaocCDFy1AuvY
xM4oanHWO2sMAAWtMvtzoDULBKnGvc4nnS+VJTTukGLIa02Q+PtL6wJU9xjDCah6yo6PzBACNj8B
0ZMV7OO2a0erGxRD2Uy5jog9GEAyZIaQWZl0eqwaHt/hZcIU+GbrDky0Wf+SI9lSFRbOrGxdiUXK
xO4JBM1cIGm/QgOttZ9JcHtCNHwBUawp3wzpEsP1HkvynSOFhozJ1jl76wboKJ4Sc1fn+zfRyhUX
z0YOFIs2/bTrv8LLuLlHqI2Ekp7zsiDXZBBFI8v4qt9d3yPH2MeqSKAp7ivocPD3sxSDsrhRys+4
jEeqkVrEH6U5z2VoGlyQ4N+pDVJBkn32Xw98TmgBfjiT9/Ab+BlBxNTA4ZXPsTmNYPLbgXMAVK2z
ev1UquHIaMiHBa5FeUd1mmhp2jmDpcjCZvjyOAEr8HT1NIz5eAIYbfjJhHxmODtxf1rvg2l/HzXG
WciG4sBYjQin2e0iQ0oT5esbCfFqy3YRGnUR/WFCGGYA+h+pRCXeeb1TpYPCWCG/pn7dIy9rnhQ/
btXVheCPCeYWE6x3IKoQgpiefnCUvV7cZi+876ueOc39JsSonN2KVh4DDrtfq6v3k0Z3I6ly49f+
UzN4/Xdu5S5/b+lm0FgS7a84uLLLDoKrv7jP/Af2wYA+75Arn7iHiimqQ0MZmXcVTX6mzGq4Xj7U
QOMZb/QvfXZtU1JGPKQFt7i7P2XQkoGi4P7rGKifJYek5YwSSOjBnbpMl3YUmCABbZC+CZ3pAEIs
ENASds6FVwGL807aVMc1e3wBdo3G/0E8znb3+I+fJwciQJT+ZyMLeHTwC85jycdQFg/McfzEqYPh
jatru11TNRwqqfe2uSYGe3iZqZPmqr19pSz5QiCKsH+5d4cqVHdd9TbhDmFrSMkfnQbIMNuIunxc
RZ8bHvpSptQkF9ODpDQS9oeKUUk8itdU/6QgcUeP5cKfzX9NraMJdCh+RPtDiBRWAoqE1kcIa6Xn
H54X/lUqNxhc5gDsLLAl+wza3PnYiqx/t1buq7suXXwEUGlNf+oGbJyPF6V30QSlJpvAR2t5nyR3
gynSvK+kspeqnst9dUfdJ5uNr0qnNY5RUWydTGwzV7GY4ArOvZttAFfn+A6nUjQaPj4rIdpFfvGE
EAxM1jIxqdprGw6oVQ03Zd0Y1/IzMOEOp8NTlG1M8v+NeWUahrXF7AiTRUDAS6KmwJRgxpE9AAvI
NF5sB4woIKw/VJWDLT0OpMC1Nxw7x0WeOhVnvbpkV8sc1/8iKkz/VuKK+24WNxT3Ck9rdzMIJM1U
my8a0iRyK3KbPrNlEbvYWtV9k9SztETHD/S1rcX8qp7TKpWUTTwz1aG1TYpZV0yZdUUdfg+8+/of
xaDjZjEC6MY319nPRwgwpAksP6zKdsXa8102qFYXJ9yqIRoR5JzkJMLcx0yruu3cvtFD//xId0Bb
F/3Qhuya3z7472DIQ8EjB5630W16bADP+o8GtX4Jb2Ixp8NTnWpqtkULPLdgfsyuCmGaBuS8sdY5
1Qp7S0ciIgbHMb3Z7I44LoJu0+IUawb1erPecZYHi6l/CA9ojs9S0RSYH7luEMJvBoDnq25LMyWw
a9cUDqlOPe6p/q5KdZQHoaEqY1AjwlS7bLRTXULtukiVkPSU94QpCSiPQBSk3AYnt+xSQqfbpm7e
mBzVaG6UmDma0gS0sd2cSeDb2jS0QHSz65y2//cayy4acu8tQ6yBj/SovA9OP2OjHbpY8iktrdxh
plxgLyu2DNur7pR+MlPUwdBvyKwEEvxBB9ptjEYWucOVzCZU069JJythL6A1vy3dj3TsGwgKRq0i
w8U1ls4pSdr/70bRG/8gPHQ2m4BvmXLA6eEZH+gOfNUy3OmEJ7yZkC0N5oU3sym7hDmjgtN/GxSb
MjEvgKBcB1eRzTNA5wjUgRcEr3stysGEVdppTuai/NBMhwenyKE+Q9FCA3//PcErMQBOM2x/VKOt
s5cmUYhlhpdHyFUlLRHRWb4dxEvNj+2UO4PsyPu1FowbrYHtNg5fUuuhFPLv26gA5jDpTStxnsdp
LVYhaeSUNB9FINnCYZwpMQ+EC4IekQj2JwtbNG78jWLpAr7A3GUCdCuW5iahg6t+FWGh2XJVRUS4
3+FbFqCHnV93UpX9JiUZEdv7m+uGrDuuQQ1x7HkL0OIIIpJzbwU4TPLECMWT2vd35YNhvYfDigLn
JPfTV5C8EB9qW5Qn5J0U2pPtpaV2bSO7JMx2rVm1H9bXP7Tqf9RlsnJ1IspYKoP5O6lhxvmiuO4V
9m3DtqhlavGSATmXhpoCFnCJfPhFeuCIZbRSCRH91PJHcazBbz7mnyqbht/V+uj2ZqwR/SJ91JIl
JWeV6nE+PssORaVvNEMGB+nexxbLVuSO4yWEwPQ4T0KVlE/Csa6FC59sobLc//ocK0RQbmGqjbo7
0pq/75GvrQcb/OOVZBYkcLhgV95hsEwLkaFyYIH63soo8s1LiZuNq1kHLOvuTuRyZJXDO/hpYfPk
eoTaxNanUVop3v3b4MelIzWEBxZjEegs/S12P6hlbxNy/a72FmHcXB8OEPMSytwCzC4qLh0lS8vU
rVz1U27Jgzz4oReehZcOyinkCU6dAMYTrm4Sx6nrwWWtjf589UsEyAmQd07aYtQI+ZMTyUe2TRm/
MT/X6eNZ3x/KsPvbu/aZVV501DMBKBnNYr7dbSkZSVSCTBgjQtCWvHqKUjTFRSpS9V1yMOhhBDWU
gLLVZusawyxY7798DVwKQi4upN65KIoRnl8gI8sCKyKLjJNrpGXaBWPoVfdof/8B2t2RmR+Nas3u
+bh4t3L1KBquoSq0rE/oHzCbYsMyPFdZFyr9KWlyrflFPhinKz6f/aQ8yhrxd/TLqNPWEkQbRp+/
bW7BhsieOf/aHvYRrf2LopKyUwhd3Y6CCh0f/IQyfMHnvCaMRW/ar/ZK/WL6/CPvHGuAbHwiaero
oSa14ar7F1u4SH8QVoB7dq3mkTYGp8ff4k+gP891/nmO5H0Xm7BsGKi44HBrLwAA2Q/G6AADYs2K
wFtwhR7Xx9xD/M1iMUbiK1pN0lmlxtJiNzsZhpWY0CNOsJKCZ3m7GnohgCSKSxMoYYWY3K/HNqSO
uGNKjM00/vljEzZnYl1+mxD8aFyCw65v+957Cmm1inEaILrLlHVMvnLnDZkRweXZ0YnQShjjoZT/
jmwKs8+WLE/54cuLgefE3pED8I2/8XOCeABHqkFBRO8ONHvWNDR0Ma6KiQ8Yx/WyOqimWdHcb0wc
tU2TRJo5V/bVYYROnfnAY1TY+h2DUFdQAxl5PzYdZw01bKtQvRgzFoRiykHkye/J2vI5+yqiaHUd
ert2XDYVficdrM7zuhoOJ7qefP0qHJ+eZXUbSF/CW8XUqB3NczapzVfwYS95zAIgN5cA6NWkP3Ic
+ZyPrdx5ffrL934ChKu2e6opE25XhX+McGF1/BfTfcKTOppCrBw6Gr/fCZo6xf1IUeqIlUU8n2qp
s2ScvLFuvmK+fRu8CeH6BMT/bqdXwi4ayO0azItp4GCkff1QcEnYTaYymtdai0iXml9XOHmwr+qI
qC+4WtWfdXHuI9EmXXSFqWfEDijI62RPT6/RBH17DOM8lc23AFCm1yiTlxtsfnZbnoiUO07lNDX7
jj+yUj46Xn+7ERDmTK4HLcYvjACu74B9xNunWvtRgizkGSk/J3lmDlpaZyQEoKZuYJQY0GKAF2hE
IuM85rdSBBQmyRAQ/1ToQ4dFPOHEz3K8dVrT5KIga3b2yulnrOVMOf0cYzkhXshfp/f2uqtjSHBz
CcA2DT+rw3nMM5KpODpaOhSkrQHWdDwt/d8rOhMvy4fgVIG34X5ge3B70wmyrJ2yTKZ82FTr171w
fDIdzinWDiiCJKaZmGrYRNP59/1mwPE+QPTRueeSy85WcXamCbBXdf5BX6v3XflOzB6HJ24XtZ3Z
Y3ttJsDhwDmLuPI+2659CuwqALD00zh8bdRwGfHhJCzEWKaVYvQn0uriG+dUZvgbtGMQZnKPDPLP
DWbIrfmNXx6F+csspgVpSXgAPi+8UHZM/nPjQERpn9KVqRcq7X46zazGzflomFvzjLWWcWpg1q8i
g0YqSS27nV4/wdQGL0aslURaqZuDOyZbwqk3NtmmSD3lbK+uZeTqVJCpothaXkBc2b7CYYmQvGel
wGOiLTvgpXTZewzaFUEReWUKtTMYmANhPZgHGDf9fZ54QqYKrbXhgiFJ7GssMRhDs14MFU7X5GLe
wWkA5kwPFuLUUjJIZl/yTy6WaDCo4NWqJfgTWMDsaqJQG5sMuLVhj0MIhIAPGlumYIFtSS6RI+SX
V74zhVFNif8zwH5giCmCoqYlR9im932hr2KHkVTzow6dT9ngRSobeR71j3uHSZN8r5pQcegDqCPi
ku99jUPNLA9/7mVn8cbCEvvmWGOFYy8p3giBjJGl/++/LbFdS/7isBwYXU3Np5xCuduu1fvAnrZr
59QahGFpVPJhuV3HwndtrIWPNjmwPUGVJMBCWQRfgzoq2SrkyHv2zWgYNP7QEmBasklCSiCjDPB/
3VQdmehzzr25bvn8ZWW7e1cwAbe2MmWLzONB2gChKQugGnlbYhXMm3ydk4Okhx/yauo3qemTdBAO
tzwFMHCVZSJtZHYZSEATBHPdvsSrXoth4eweykPIbaVRZYslBpOneFfd/LDJdc7t1+5YeRkocWWr
fUSqGMOxiwMyytazn5niCZDrlAv3NsoexZ0pvlcxooz7T1MSw0TMxLn5XwwefqhY/PYppV1/fyW6
nXCRUAYicDej822md2ew02UmgdVn5g/D5PQmgPlO5b2vxU0Yhb8vFM/ilI/v/vYxuNPGUmLKT71J
HoexxlquWbeyVEsxOAKjOUtk0aCBqkQEMnFeaVNZoc8bXzaFtq0dSRv98/oroQ6gHkhKEDaXQ7Eo
JMnL8KxlAQPu2X9LMveo14MkXb3SRK/UKIrGWPbM9xln99pQHuRQstxotcoQIcYhXv3lcBsAXX4n
m+wehQtac1pbvHEIxh1K+A4BWUe1ehSkKDHhToLn23rVL8Un85bNCQ7S52Cut1Enlhr7AA5xBSq5
S4Trvqo78colOk91sOYxoGBp/DrC1vs7f7jxguW/0nAf+2WevpneytlNubK7KZpemx9Y3xaPejmg
lAHjvgxKukyaL8MZHm8rzphs69dvToi4ZR8RifQOcJPeKlcR42Hx2k/+TrqbpO9I6h61qSkRVfYN
69w6Qp0mKIDWmD8WSWpdzbcVRCgmj13z9juBxX+THw2isJo+cHuEv2A7MprHgEUDTbSSy0Gr3u3t
QoEbPrIS72r98Qq/oe0Rcq0H2TUxb48Si0jLQ/SoVvhBRTiJ73yrc2NA8YY0cZGwZps8OY7qAsq8
rSJlKvbRr/TxppPFkQ4U7GsTowB1Rdqr5ART0ftOfHdFXqjfOjRefPSE27yU8j9kVaSQq0dQxEPZ
oBp+BAIscPlytdsm0S8nonXi/VqOyrzI6lew6fSZdy5CdhI9wF72+cI/eSh7u+nisqRGlf/X8U7o
52wmhwPtTmPjF7USA0onUN88UQFOqJWdatPteE5B4uLM/hfoS6wnuIPJBhncsX6PzwEcNYo9zJHe
bXfuLo5+6OSTuhsM3PEpZfKcuk41yZYi8qRyzVopgPycjRt9DVfel5ZsyMvjx5JJD86Ax/wh1KKs
liZwtR3MZ/fc+rEVQZVBPcQp3b3Z6S+2794SWObibv1S+rZfEf4zzYURC2xLcmf1EfG1qUYfdCQ8
fqm8ctsNxoQPD86rjwy1hZ3SVsf1IViDACVVsxfESCdN2u4wIpUagcAy4Uo02vceAv1Ruts571F1
NYMrgkg731ofu36hYHbN9aXcYiQ9fDUiG/ogtRE3Luzu6gQ2NJjkMTxJNmbdmv/yMn9jTzSG2vtm
NnEaqtLrvD3qXl/9gonLHRTgcf149a+NamsRSmK2uzMwabIeyOA2X5hRgmLgSpEzqZPZCJxTtlPM
KofEYWgoicX2QyUUSxx8ORK85zffR648GHZr02OgPejrIOcvVfLIBTfyNGGVUz+ww4IzLjsskIEQ
zmF9B5iJ51E/5o4I85zSwWNhGsUtklAWnnatxMjgggbvurAcsKTYO9Q1kRzQ8DMWKwA1G1MFoerp
3/VbpktGJBJhL1R6qGoIbaWpzkKK0lPQTi2cXvQo1fcR10lDiJfRomKfjnXFefp4qfBAvdDHZ/bC
17oWoh1eCbImUadsE/hfCpiOZQFtzHDXnLNNv3ipX/U2S7rUrs3oPRsI8hO42IRHdoIbfXbf1Aw5
3x7EkzFpmU62pPssAYgEIAZhvvX9en9QVeVHyM0A2z7FqWlpsMMx1MLlT16DIkbGRhcOSMR1i8CW
0xtMqumRUgcj4rxRIU+8muNVr8Xp7adkb6RmiJ/ldbIFfKlqVEc7KdbieuEX7w9Hq31OMbrXxdWR
167A3dQ+SVxjjkGH6sc52+EKI3P38EUg+WT1r8tQfPcBHIYl+ZKkfMEvFDsWELjFUdMT6jqZXhYF
22bjeIFaTcfqFomaPWfZj/wT/mabg+2LIUyuySDLKI8MeIrzBoarIStwNEuSA+kAPxDb4VrPG3Wd
g/FIwRBL9qcGMk+9tOXo2avWFwaGGhNssAJI+8vXcatM8bRTeuL5+87pT9/dNZV30wMGyV6orDMM
dkHS+A12C/0kwaQt7nKqsHPXkAmbLAWM5+yywbYuKTgO6KzXqKDjTuVJJuK7CL4U6nZ46Ml094/S
mWRPqqNARtNZQpM4dHJ1z2QLaKa5NHPiMO0ZblGdgbsKeWOoEZW5bymLawhkP/148mqJ0wISqlkF
TBd5B8y0YwzR7VSPhEkZOEF+GXq940/8UHnDiUyOBx4Rlwv/EzgkhlWYiWOqKmSaAelN+j4n+RC0
WqI2S3UsHZ237F99N16U4F7WI+Zh/bP0Wyi1UABwBA+zPJGH61rDFD5wXlMB1LmwI+C8AvbbMEge
+zbjsiA111E72vxsIH1Sh3BnCq2Mgo6SDLS7kEA+l67Q6L3nYtWyOG7+KjPmiU+UQtRw2LCR7z9A
xxc0w90Mslf4xza9F6L8gFoRZzQP5I/78GU97HqSa1fUyL8LEULm1uLeNs+BbKWCHlRNoyUmYgv6
qOhX61bJuiA/4VsErCUkTObLzmF8ZSJxin4in9aWIr2l5Eb31dSELY8y+4gU6NYe5xk99zNoDwbI
u4mL0TQ0++xlzIoEoAVQxGMhJRmGycwaI0PvDsVBGENhPOp3Qyrs2IAZqmuBfoc4Y3WP9r3HU/JJ
Le7hekHH8xU59iLyv4qWK055wuGyvEgh3sA8L0FKg2vxMIVlAPYShKGL/RwwZZVc4kjc0sFLImXp
KJUlQkD0Pe7tl8CJrjba6OhPQPYUH07MqL3AWROA44iDRD1hprvU9dKGt7jBW9edfa8n6yrdOh8b
cWqx/W9M/yuJbCtP6saYxg/48Kqk1H9GbI+tk4jhYkVE91ydKW7b1s1eSmqT7v8BB5MiWerP7gnD
WuxWO+TiEJZPAiAW7QwHwfljP+0zbtnSeHPZJIWpsyOB0C+jRrq2vXrDo7ruL1JQ4urZRgYvMkH1
R/CmqXl47G/qUuDQU0rZ6N3lUiTtdFq0kTUiV+Bq/uqvPg3vO53IO9tXZcp0kIV+7xMqMkDT8Ng2
j6NH9J1S/fJ+ZGNN73Hl24KUsdcAM9jywD5+By0DBmbjDP1ChzB3yZROTCAHLD1vsj4AEsnMQQbL
axqscKzlshfRN72zXGoFVrp6prbtJarbGEtj5erfQ+IbLwZE6T0i64P8oCq6ym6wFXluwml7gB8F
Oqgclgazm2RDqL78KezLk1ObtFiOZRzGD9DDY9aNeybKItdovSPgRCuQdoo92SMLKD/qmqhlOu8f
8lhpFDhqtF0z78Ft5kJXd+4EUuCuts0CnxSDfGSP4iIFkN045TpVCckSHm+DwWcc1n6S8nh7f8gY
DBI6uLJ0e+sSQ7xKMo8hnJD1lCbmKTdCMMep1RpIc0UaPomQnasdNX+zO7WEZScmFVkOvp72zCQk
/Tt5oMCegRDKtAsIlqoLjDe24C/uEb6aVmimUA4wsswaeqcIK39Ui8pzRtCU8vC/KKiASvLNrZO+
B2s84eAHNrYIGcJPqdIScTxXDaT47iOr3dwHl8NFLks1BDY6kF58DpZygC9apbjwXvEViZz/7W8U
JcT3l1Zvzvny173NZlBHOpSQh0K4Hc+k6McOuq0iFUGxYyBHSWP90sSZ4CEXjcik0ECAMvi0guoA
SsC7um+ZJj+yK6A1j309CbEVVTWuoZY=
`protect end_protected

